

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589;

  NOR2_X2 U323 ( .A1(n473), .A2(n472), .ZN(n474) );
  NOR2_X1 U324 ( .A1(n533), .A2(n567), .ZN(n572) );
  XNOR2_X1 U325 ( .A(n364), .B(n363), .ZN(n369) );
  XNOR2_X1 U326 ( .A(n308), .B(n307), .ZN(n429) );
  XNOR2_X1 U327 ( .A(n306), .B(KEYINPUT84), .ZN(n307) );
  XOR2_X1 U328 ( .A(n485), .B(KEYINPUT36), .Z(n473) );
  XNOR2_X1 U329 ( .A(n443), .B(n442), .ZN(n533) );
  NAND2_X1 U330 ( .A1(n566), .A2(n565), .ZN(n291) );
  AND2_X1 U331 ( .A1(G232GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U332 ( .A(KEYINPUT47), .B(KEYINPUT109), .ZN(n377) );
  XNOR2_X1 U333 ( .A(n378), .B(n377), .ZN(n384) );
  XNOR2_X1 U334 ( .A(n362), .B(KEYINPUT31), .ZN(n364) );
  XNOR2_X1 U335 ( .A(n336), .B(n292), .ZN(n337) );
  XNOR2_X1 U336 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U337 ( .A(G99GAT), .B(G85GAT), .Z(n370) );
  XNOR2_X1 U338 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U339 ( .A(n439), .B(n438), .ZN(n441) );
  NOR2_X1 U340 ( .A1(n450), .A2(n457), .ZN(n445) );
  INV_X1 U341 ( .A(G218GAT), .ZN(n446) );
  XOR2_X1 U342 ( .A(n345), .B(n349), .Z(n485) );
  XNOR2_X1 U343 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U344 ( .A(n452), .B(G190GAT), .ZN(n453) );
  XNOR2_X1 U345 ( .A(n477), .B(G43GAT), .ZN(n478) );
  XNOR2_X1 U346 ( .A(n449), .B(n448), .ZN(G1355GAT) );
  XNOR2_X1 U347 ( .A(n454), .B(n453), .ZN(G1351GAT) );
  XNOR2_X1 U348 ( .A(n479), .B(n478), .ZN(G1330GAT) );
  XOR2_X1 U349 ( .A(G169GAT), .B(G8GAT), .Z(n352) );
  XOR2_X1 U350 ( .A(n352), .B(KEYINPUT93), .Z(n294) );
  NAND2_X1 U351 ( .A1(G226GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U352 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U353 ( .A(G92GAT), .B(G64GAT), .Z(n296) );
  XNOR2_X1 U354 ( .A(G204GAT), .B(KEYINPUT71), .ZN(n295) );
  XNOR2_X1 U355 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U356 ( .A(G176GAT), .B(n297), .Z(n363) );
  XOR2_X1 U357 ( .A(n298), .B(n363), .Z(n304) );
  XNOR2_X1 U358 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n299) );
  XNOR2_X1 U359 ( .A(n299), .B(KEYINPUT87), .ZN(n300) );
  XOR2_X1 U360 ( .A(n300), .B(KEYINPUT88), .Z(n302) );
  XNOR2_X1 U361 ( .A(G197GAT), .B(G218GAT), .ZN(n301) );
  XNOR2_X1 U362 ( .A(n302), .B(n301), .ZN(n418) );
  XNOR2_X1 U363 ( .A(G36GAT), .B(n418), .ZN(n303) );
  XNOR2_X1 U364 ( .A(n304), .B(n303), .ZN(n310) );
  XNOR2_X1 U365 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n305) );
  XNOR2_X1 U366 ( .A(n305), .B(KEYINPUT18), .ZN(n308) );
  XNOR2_X1 U367 ( .A(G183GAT), .B(G190GAT), .ZN(n306) );
  INV_X1 U368 ( .A(n429), .ZN(n309) );
  XOR2_X1 U369 ( .A(n310), .B(n309), .Z(n501) );
  XNOR2_X1 U370 ( .A(KEYINPUT111), .B(KEYINPUT48), .ZN(n386) );
  XOR2_X1 U371 ( .A(KEYINPUT15), .B(KEYINPUT74), .Z(n312) );
  XNOR2_X1 U372 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n311) );
  XNOR2_X1 U373 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U374 ( .A(KEYINPUT76), .B(KEYINPUT78), .Z(n314) );
  XNOR2_X1 U375 ( .A(KEYINPUT14), .B(KEYINPUT75), .ZN(n313) );
  XNOR2_X1 U376 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n316), .B(n315), .ZN(n329) );
  XOR2_X1 U378 ( .A(G78GAT), .B(G211GAT), .Z(n318) );
  XNOR2_X1 U379 ( .A(G127GAT), .B(G155GAT), .ZN(n317) );
  XNOR2_X1 U380 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U381 ( .A(G57GAT), .B(G183GAT), .Z(n320) );
  XNOR2_X1 U382 ( .A(G1GAT), .B(G8GAT), .ZN(n319) );
  XNOR2_X1 U383 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U384 ( .A(n322), .B(n321), .Z(n327) );
  XOR2_X1 U385 ( .A(G22GAT), .B(G15GAT), .Z(n355) );
  XOR2_X1 U386 ( .A(G71GAT), .B(KEYINPUT13), .Z(n361) );
  XOR2_X1 U387 ( .A(KEYINPUT77), .B(n361), .Z(n324) );
  NAND2_X1 U388 ( .A1(G231GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U389 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U390 ( .A(n355), .B(n325), .ZN(n326) );
  XNOR2_X1 U391 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U392 ( .A(n329), .B(n328), .Z(n586) );
  INV_X1 U393 ( .A(n586), .ZN(n558) );
  XOR2_X1 U394 ( .A(KEYINPUT72), .B(KEYINPUT9), .Z(n331) );
  XNOR2_X1 U395 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(n330) );
  XNOR2_X1 U396 ( .A(n331), .B(n330), .ZN(n340) );
  XOR2_X1 U397 ( .A(n370), .B(G92GAT), .Z(n333) );
  XOR2_X1 U398 ( .A(G134GAT), .B(KEYINPUT73), .Z(n391) );
  XNOR2_X1 U399 ( .A(G218GAT), .B(n391), .ZN(n332) );
  XNOR2_X1 U400 ( .A(n333), .B(n332), .ZN(n338) );
  XOR2_X1 U401 ( .A(G106GAT), .B(G162GAT), .Z(n335) );
  XNOR2_X1 U402 ( .A(G29GAT), .B(G190GAT), .ZN(n334) );
  XNOR2_X1 U403 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U404 ( .A(n340), .B(n339), .ZN(n345) );
  XOR2_X1 U405 ( .A(G36GAT), .B(KEYINPUT69), .Z(n342) );
  XNOR2_X1 U406 ( .A(G50GAT), .B(G43GAT), .ZN(n341) );
  XNOR2_X1 U407 ( .A(n342), .B(n341), .ZN(n344) );
  XOR2_X1 U408 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n343) );
  XOR2_X1 U409 ( .A(n344), .B(n343), .Z(n349) );
  XOR2_X1 U410 ( .A(KEYINPUT46), .B(KEYINPUT108), .Z(n374) );
  XOR2_X1 U411 ( .A(KEYINPUT29), .B(KEYINPUT66), .Z(n347) );
  XNOR2_X1 U412 ( .A(KEYINPUT68), .B(KEYINPUT67), .ZN(n346) );
  XNOR2_X1 U413 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U414 ( .A(n349), .B(n348), .ZN(n360) );
  XOR2_X1 U415 ( .A(G1GAT), .B(G113GAT), .Z(n351) );
  XNOR2_X1 U416 ( .A(G29GAT), .B(G141GAT), .ZN(n350) );
  XNOR2_X1 U417 ( .A(n351), .B(n350), .ZN(n403) );
  XOR2_X1 U418 ( .A(n403), .B(n352), .Z(n354) );
  NAND2_X1 U419 ( .A1(G229GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U420 ( .A(n354), .B(n353), .ZN(n356) );
  XOR2_X1 U421 ( .A(n356), .B(n355), .Z(n358) );
  XNOR2_X1 U422 ( .A(G197GAT), .B(KEYINPUT30), .ZN(n357) );
  XNOR2_X1 U423 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U424 ( .A(n360), .B(n359), .Z(n551) );
  INV_X1 U425 ( .A(n551), .ZN(n577) );
  XOR2_X1 U426 ( .A(n361), .B(KEYINPUT33), .Z(n362) );
  XNOR2_X1 U427 ( .A(G120GAT), .B(G148GAT), .ZN(n365) );
  XNOR2_X1 U428 ( .A(n365), .B(G57GAT), .ZN(n398) );
  XOR2_X1 U429 ( .A(n398), .B(KEYINPUT32), .Z(n367) );
  NAND2_X1 U430 ( .A1(G230GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U431 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U432 ( .A(n369), .B(n368), .Z(n372) );
  XOR2_X1 U433 ( .A(G106GAT), .B(G78GAT), .Z(n410) );
  XNOR2_X1 U434 ( .A(n410), .B(n370), .ZN(n371) );
  XNOR2_X1 U435 ( .A(n372), .B(n371), .ZN(n580) );
  XOR2_X1 U436 ( .A(KEYINPUT41), .B(n580), .Z(n553) );
  INV_X1 U437 ( .A(n553), .ZN(n565) );
  NAND2_X1 U438 ( .A1(n577), .A2(n565), .ZN(n373) );
  XNOR2_X1 U439 ( .A(n374), .B(n373), .ZN(n375) );
  NOR2_X1 U440 ( .A1(n485), .A2(n375), .ZN(n376) );
  NAND2_X1 U441 ( .A1(n558), .A2(n376), .ZN(n378) );
  NOR2_X1 U442 ( .A1(n558), .A2(n473), .ZN(n379) );
  XNOR2_X1 U443 ( .A(KEYINPUT45), .B(n379), .ZN(n380) );
  NAND2_X1 U444 ( .A1(n380), .A2(n580), .ZN(n381) );
  XOR2_X1 U445 ( .A(KEYINPUT110), .B(n381), .Z(n382) );
  XOR2_X1 U446 ( .A(KEYINPUT70), .B(n577), .Z(n536) );
  NAND2_X1 U447 ( .A1(n382), .A2(n536), .ZN(n383) );
  NAND2_X1 U448 ( .A1(n384), .A2(n383), .ZN(n385) );
  XNOR2_X1 U449 ( .A(n386), .B(n385), .ZN(n531) );
  NOR2_X1 U450 ( .A1(n501), .A2(n531), .ZN(n387) );
  XNOR2_X1 U451 ( .A(KEYINPUT54), .B(n387), .ZN(n406) );
  XOR2_X1 U452 ( .A(KEYINPUT1), .B(KEYINPUT91), .Z(n389) );
  XNOR2_X1 U453 ( .A(G85GAT), .B(KEYINPUT4), .ZN(n388) );
  XNOR2_X1 U454 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U455 ( .A(n391), .B(n390), .Z(n393) );
  NAND2_X1 U456 ( .A1(G225GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U457 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U458 ( .A(n394), .B(KEYINPUT6), .Z(n397) );
  XNOR2_X1 U459 ( .A(G127GAT), .B(KEYINPUT0), .ZN(n395) );
  XNOR2_X1 U460 ( .A(n395), .B(KEYINPUT80), .ZN(n431) );
  XNOR2_X1 U461 ( .A(n431), .B(KEYINPUT5), .ZN(n396) );
  XNOR2_X1 U462 ( .A(n397), .B(n396), .ZN(n399) );
  XOR2_X1 U463 ( .A(n399), .B(n398), .Z(n405) );
  XOR2_X1 U464 ( .A(KEYINPUT2), .B(G162GAT), .Z(n401) );
  XNOR2_X1 U465 ( .A(KEYINPUT89), .B(G155GAT), .ZN(n400) );
  XNOR2_X1 U466 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U467 ( .A(KEYINPUT3), .B(n402), .Z(n422) );
  XNOR2_X1 U468 ( .A(n403), .B(n422), .ZN(n404) );
  XNOR2_X1 U469 ( .A(n405), .B(n404), .ZN(n462) );
  XOR2_X1 U470 ( .A(KEYINPUT92), .B(n462), .Z(n520) );
  INV_X1 U471 ( .A(n520), .ZN(n480) );
  NAND2_X1 U472 ( .A1(n406), .A2(n480), .ZN(n407) );
  XNOR2_X1 U473 ( .A(n407), .B(KEYINPUT64), .ZN(n450) );
  XOR2_X1 U474 ( .A(G204GAT), .B(KEYINPUT22), .Z(n409) );
  XNOR2_X1 U475 ( .A(G141GAT), .B(G148GAT), .ZN(n408) );
  XNOR2_X1 U476 ( .A(n409), .B(n408), .ZN(n411) );
  XOR2_X1 U477 ( .A(n411), .B(n410), .Z(n413) );
  XNOR2_X1 U478 ( .A(G50GAT), .B(G22GAT), .ZN(n412) );
  XNOR2_X1 U479 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U480 ( .A(KEYINPUT23), .B(KEYINPUT90), .Z(n415) );
  NAND2_X1 U481 ( .A1(G228GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U482 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U483 ( .A(n417), .B(n416), .Z(n420) );
  XNOR2_X1 U484 ( .A(n418), .B(KEYINPUT24), .ZN(n419) );
  XNOR2_X1 U485 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U486 ( .A(n422), .B(n421), .ZN(n464) );
  XOR2_X1 U487 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n424) );
  XNOR2_X1 U488 ( .A(G169GAT), .B(KEYINPUT83), .ZN(n423) );
  XNOR2_X1 U489 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U490 ( .A(KEYINPUT85), .B(G71GAT), .Z(n426) );
  XNOR2_X1 U491 ( .A(KEYINPUT20), .B(G176GAT), .ZN(n425) );
  XNOR2_X1 U492 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U493 ( .A(n428), .B(n427), .ZN(n443) );
  INV_X1 U494 ( .A(G15GAT), .ZN(n430) );
  XNOR2_X1 U495 ( .A(n430), .B(n429), .ZN(n439) );
  XOR2_X1 U496 ( .A(KEYINPUT65), .B(n431), .Z(n437) );
  XOR2_X1 U497 ( .A(G120GAT), .B(KEYINPUT86), .Z(n433) );
  XNOR2_X1 U498 ( .A(G113GAT), .B(G99GAT), .ZN(n432) );
  XNOR2_X1 U499 ( .A(n433), .B(n432), .ZN(n435) );
  XOR2_X1 U500 ( .A(G43GAT), .B(G134GAT), .Z(n434) );
  XNOR2_X1 U501 ( .A(n435), .B(n434), .ZN(n436) );
  NAND2_X1 U502 ( .A1(G227GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U503 ( .A(n441), .B(n440), .ZN(n442) );
  NAND2_X1 U504 ( .A1(n464), .A2(n533), .ZN(n444) );
  XOR2_X1 U505 ( .A(n444), .B(KEYINPUT26), .Z(n549) );
  INV_X1 U506 ( .A(n549), .ZN(n457) );
  XOR2_X1 U507 ( .A(KEYINPUT120), .B(n445), .Z(n581) );
  NOR2_X1 U508 ( .A1(n581), .A2(n473), .ZN(n449) );
  XNOR2_X1 U509 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n447) );
  NOR2_X1 U510 ( .A1(n450), .A2(n464), .ZN(n451) );
  XNOR2_X1 U511 ( .A(n451), .B(KEYINPUT55), .ZN(n567) );
  NAND2_X1 U512 ( .A1(n572), .A2(n485), .ZN(n454) );
  XOR2_X1 U513 ( .A(KEYINPUT119), .B(KEYINPUT58), .Z(n452) );
  INV_X1 U514 ( .A(KEYINPUT38), .ZN(n476) );
  INV_X1 U515 ( .A(KEYINPUT94), .ZN(n461) );
  NOR2_X1 U516 ( .A1(n533), .A2(n501), .ZN(n455) );
  NOR2_X1 U517 ( .A1(n464), .A2(n455), .ZN(n456) );
  XOR2_X1 U518 ( .A(KEYINPUT25), .B(n456), .Z(n459) );
  INV_X1 U519 ( .A(n501), .ZN(n522) );
  XOR2_X1 U520 ( .A(n522), .B(KEYINPUT27), .Z(n465) );
  NOR2_X1 U521 ( .A1(n457), .A2(n465), .ZN(n458) );
  NOR2_X1 U522 ( .A1(n459), .A2(n458), .ZN(n460) );
  XNOR2_X1 U523 ( .A(n461), .B(n460), .ZN(n463) );
  NAND2_X1 U524 ( .A1(n463), .A2(n462), .ZN(n468) );
  XOR2_X1 U525 ( .A(KEYINPUT28), .B(n464), .Z(n503) );
  INV_X1 U526 ( .A(n503), .ZN(n532) );
  OR2_X1 U527 ( .A1(n480), .A2(n465), .ZN(n530) );
  NOR2_X1 U528 ( .A1(n532), .A2(n530), .ZN(n466) );
  NAND2_X1 U529 ( .A1(n466), .A2(n533), .ZN(n467) );
  NAND2_X1 U530 ( .A1(n468), .A2(n467), .ZN(n469) );
  XNOR2_X1 U531 ( .A(n469), .B(KEYINPUT95), .ZN(n489) );
  NOR2_X1 U532 ( .A1(n489), .A2(n586), .ZN(n470) );
  XNOR2_X1 U533 ( .A(n470), .B(KEYINPUT100), .ZN(n471) );
  INV_X1 U534 ( .A(n471), .ZN(n472) );
  XNOR2_X1 U535 ( .A(KEYINPUT37), .B(n474), .ZN(n519) );
  INV_X1 U536 ( .A(n536), .ZN(n563) );
  NAND2_X1 U537 ( .A1(n580), .A2(n563), .ZN(n490) );
  NOR2_X1 U538 ( .A1(n519), .A2(n490), .ZN(n475) );
  XNOR2_X1 U539 ( .A(n476), .B(n475), .ZN(n504) );
  NOR2_X1 U540 ( .A1(n533), .A2(n504), .ZN(n479) );
  XNOR2_X1 U541 ( .A(KEYINPUT40), .B(KEYINPUT101), .ZN(n477) );
  INV_X1 U542 ( .A(G29GAT), .ZN(n484) );
  NOR2_X1 U543 ( .A1(n504), .A2(n480), .ZN(n482) );
  XNOR2_X1 U544 ( .A(KEYINPUT99), .B(KEYINPUT39), .ZN(n481) );
  XNOR2_X1 U545 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U546 ( .A(n484), .B(n483), .ZN(G1328GAT) );
  XNOR2_X1 U547 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n493) );
  XOR2_X1 U548 ( .A(KEYINPUT79), .B(KEYINPUT16), .Z(n487) );
  INV_X1 U549 ( .A(n485), .ZN(n561) );
  NAND2_X1 U550 ( .A1(n561), .A2(n586), .ZN(n486) );
  XNOR2_X1 U551 ( .A(n487), .B(n486), .ZN(n488) );
  OR2_X1 U552 ( .A1(n489), .A2(n488), .ZN(n508) );
  NOR2_X1 U553 ( .A1(n490), .A2(n508), .ZN(n491) );
  XNOR2_X1 U554 ( .A(KEYINPUT96), .B(n491), .ZN(n498) );
  NAND2_X1 U555 ( .A1(n520), .A2(n498), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n493), .B(n492), .ZN(G1324GAT) );
  XOR2_X1 U557 ( .A(G8GAT), .B(KEYINPUT97), .Z(n495) );
  NAND2_X1 U558 ( .A1(n498), .A2(n522), .ZN(n494) );
  XNOR2_X1 U559 ( .A(n495), .B(n494), .ZN(G1325GAT) );
  XOR2_X1 U560 ( .A(G15GAT), .B(KEYINPUT35), .Z(n497) );
  INV_X1 U561 ( .A(n533), .ZN(n566) );
  NAND2_X1 U562 ( .A1(n498), .A2(n566), .ZN(n496) );
  XNOR2_X1 U563 ( .A(n497), .B(n496), .ZN(G1326GAT) );
  NAND2_X1 U564 ( .A1(n498), .A2(n532), .ZN(n499) );
  XNOR2_X1 U565 ( .A(n499), .B(KEYINPUT98), .ZN(n500) );
  XNOR2_X1 U566 ( .A(G22GAT), .B(n500), .ZN(G1327GAT) );
  NOR2_X1 U567 ( .A1(n501), .A2(n504), .ZN(n502) );
  XOR2_X1 U568 ( .A(G36GAT), .B(n502), .Z(G1329GAT) );
  NOR2_X1 U569 ( .A1(n504), .A2(n503), .ZN(n505) );
  XOR2_X1 U570 ( .A(G50GAT), .B(n505), .Z(G1331GAT) );
  XNOR2_X1 U571 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n506), .B(KEYINPUT103), .ZN(n507) );
  XOR2_X1 U573 ( .A(KEYINPUT102), .B(n507), .Z(n510) );
  NAND2_X1 U574 ( .A1(n551), .A2(n565), .ZN(n518) );
  NOR2_X1 U575 ( .A1(n518), .A2(n508), .ZN(n513) );
  NAND2_X1 U576 ( .A1(n513), .A2(n520), .ZN(n509) );
  XNOR2_X1 U577 ( .A(n510), .B(n509), .ZN(G1332GAT) );
  NAND2_X1 U578 ( .A1(n522), .A2(n513), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n511), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U580 ( .A1(n566), .A2(n513), .ZN(n512) );
  XNOR2_X1 U581 ( .A(n512), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U582 ( .A(KEYINPUT104), .B(KEYINPUT43), .Z(n515) );
  NAND2_X1 U583 ( .A1(n513), .A2(n532), .ZN(n514) );
  XNOR2_X1 U584 ( .A(n515), .B(n514), .ZN(n517) );
  XOR2_X1 U585 ( .A(G78GAT), .B(KEYINPUT105), .Z(n516) );
  XNOR2_X1 U586 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NOR2_X1 U587 ( .A1(n519), .A2(n518), .ZN(n525) );
  NAND2_X1 U588 ( .A1(n520), .A2(n525), .ZN(n521) );
  XNOR2_X1 U589 ( .A(G85GAT), .B(n521), .ZN(G1336GAT) );
  NAND2_X1 U590 ( .A1(n522), .A2(n525), .ZN(n523) );
  XNOR2_X1 U591 ( .A(n523), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U592 ( .A1(n566), .A2(n525), .ZN(n524) );
  XNOR2_X1 U593 ( .A(n524), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n529) );
  XOR2_X1 U595 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n527) );
  NAND2_X1 U596 ( .A1(n525), .A2(n532), .ZN(n526) );
  XNOR2_X1 U597 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U598 ( .A(n529), .B(n528), .ZN(G1339GAT) );
  NOR2_X1 U599 ( .A1(n531), .A2(n530), .ZN(n550) );
  NOR2_X1 U600 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U601 ( .A1(n550), .A2(n534), .ZN(n535) );
  XNOR2_X1 U602 ( .A(KEYINPUT112), .B(n535), .ZN(n544) );
  NOR2_X1 U603 ( .A1(n544), .A2(n536), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n537), .B(KEYINPUT113), .ZN(n538) );
  XNOR2_X1 U605 ( .A(G113GAT), .B(n538), .ZN(G1340GAT) );
  XNOR2_X1 U606 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n540) );
  NOR2_X1 U607 ( .A1(n553), .A2(n544), .ZN(n539) );
  XNOR2_X1 U608 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  XNOR2_X1 U609 ( .A(KEYINPUT50), .B(KEYINPUT114), .ZN(n542) );
  NOR2_X1 U610 ( .A1(n558), .A2(n544), .ZN(n541) );
  XNOR2_X1 U611 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U612 ( .A(G127GAT), .B(n543), .Z(G1342GAT) );
  NOR2_X1 U613 ( .A1(n544), .A2(n561), .ZN(n548) );
  XOR2_X1 U614 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n546) );
  XNOR2_X1 U615 ( .A(G134GAT), .B(KEYINPUT116), .ZN(n545) );
  XNOR2_X1 U616 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U617 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  NAND2_X1 U618 ( .A1(n550), .A2(n549), .ZN(n560) );
  NOR2_X1 U619 ( .A1(n551), .A2(n560), .ZN(n552) );
  XOR2_X1 U620 ( .A(G141GAT), .B(n552), .Z(G1344GAT) );
  NOR2_X1 U621 ( .A1(n560), .A2(n553), .ZN(n557) );
  XOR2_X1 U622 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n555) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n554) );
  XNOR2_X1 U624 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  NOR2_X1 U626 ( .A1(n558), .A2(n560), .ZN(n559) );
  XOR2_X1 U627 ( .A(G155GAT), .B(n559), .Z(G1346GAT) );
  NOR2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U629 ( .A(G162GAT), .B(n562), .Z(G1347GAT) );
  NAND2_X1 U630 ( .A1(n563), .A2(n572), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(G169GAT), .ZN(G1348GAT) );
  XNOR2_X1 U632 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT56), .B(KEYINPUT118), .Z(n569) );
  OR2_X1 U634 ( .A1(n291), .A2(n567), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1349GAT) );
  NAND2_X1 U637 ( .A1(n586), .A2(n572), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT122), .Z(n575) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT121), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XOR2_X1 U642 ( .A(KEYINPUT59), .B(n576), .Z(n579) );
  INV_X1 U643 ( .A(n581), .ZN(n587) );
  NAND2_X1 U644 ( .A1(n577), .A2(n587), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n585) );
  XOR2_X1 U647 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n583) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT124), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  XOR2_X1 U651 ( .A(G211GAT), .B(KEYINPUT125), .Z(n589) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(G1354GAT) );
endmodule

