//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963;
  OR3_X1    g000(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n202));
  OAI21_X1  g001(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n203));
  AOI22_X1  g002(.A1(new_n202), .A2(new_n203), .B1(G29gat), .B2(G36gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT15), .ZN(new_n205));
  XOR2_X1   g004(.A(G43gat), .B(G50gat), .Z(new_n206));
  OR3_X1    g005(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n206), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT15), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n206), .A2(new_n205), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(new_n210), .A3(new_n204), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT17), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(G15gat), .B(G22gat), .Z(new_n215));
  INV_X1    g014(.A(G1gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT82), .ZN(new_n218));
  XNOR2_X1  g017(.A(G15gat), .B(G22gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT16), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n219), .B1(new_n220), .B2(G1gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n218), .A2(new_n222), .A3(G8gat), .ZN(new_n223));
  INV_X1    g022(.A(G8gat), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n217), .B(new_n221), .C1(KEYINPUT82), .C2(new_n224), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n207), .A2(new_n211), .A3(KEYINPUT17), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n214), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n223), .A2(new_n225), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(new_n212), .ZN(new_n230));
  NAND2_X1  g029(.A1(G229gat), .A2(G233gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n228), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT18), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT11), .B(G169gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n235), .B(G197gat), .ZN(new_n236));
  XOR2_X1   g035(.A(G113gat), .B(G141gat), .Z(new_n237));
  XOR2_X1   g036(.A(new_n236), .B(new_n237), .Z(new_n238));
  XOR2_X1   g037(.A(new_n238), .B(KEYINPUT12), .Z(new_n239));
  XNOR2_X1  g038(.A(new_n229), .B(new_n212), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n231), .B(KEYINPUT83), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(KEYINPUT13), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n228), .A2(KEYINPUT18), .A3(new_n230), .A4(new_n231), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n234), .A2(new_n239), .A3(new_n244), .A4(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT84), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n246), .A2(new_n247), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n239), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n234), .A2(new_n244), .A3(new_n245), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G99gat), .A2(G106gat), .ZN(new_n254));
  INV_X1    g053(.A(G85gat), .ZN(new_n255));
  INV_X1    g054(.A(G92gat), .ZN(new_n256));
  AOI22_X1  g055(.A1(KEYINPUT8), .A2(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT87), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G99gat), .B(G106gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(KEYINPUT88), .ZN(new_n261));
  NAND2_X1  g060(.A1(G85gat), .A2(G92gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(KEYINPUT7), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n259), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT89), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n259), .A2(new_n263), .ZN(new_n267));
  INV_X1    g066(.A(new_n261), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n267), .A2(KEYINPUT90), .A3(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT90), .ZN(new_n270));
  INV_X1    g069(.A(new_n263), .ZN(new_n271));
  OR2_X1    g070(.A1(new_n257), .A2(new_n258), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n258), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n270), .B1(new_n274), .B2(new_n261), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(KEYINPUT89), .A3(new_n261), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n266), .A2(new_n269), .A3(new_n275), .A4(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(KEYINPUT85), .B1(G71gat), .B2(G78gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(G57gat), .B(G64gat), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G71gat), .B(G78gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n283), .B1(new_n261), .B2(new_n274), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n267), .A2(new_n268), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n277), .A2(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(G230gat), .A2(G233gat), .ZN(new_n287));
  XOR2_X1   g086(.A(new_n287), .B(KEYINPUT94), .Z(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NOR3_X1   g088(.A1(new_n286), .A2(KEYINPUT95), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n283), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n266), .A2(new_n276), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n269), .A2(new_n275), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT91), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT91), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n277), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g095(.A(KEYINPUT10), .B(new_n291), .C1(new_n294), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT93), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT10), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n286), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n292), .A2(new_n293), .A3(KEYINPUT91), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n277), .A2(new_n295), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT93), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n303), .A2(new_n304), .A3(KEYINPUT10), .A4(new_n291), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n298), .A2(new_n300), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n290), .B1(new_n306), .B2(new_n289), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT95), .B1(new_n286), .B2(new_n289), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G120gat), .B(G148gat), .ZN(new_n310));
  INV_X1    g109(.A(G176gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n310), .B(new_n311), .ZN(new_n312));
  XOR2_X1   g111(.A(new_n312), .B(G204gat), .Z(new_n313));
  NAND2_X1  g112(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n313), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n307), .A2(new_n315), .A3(new_n308), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT4), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT1), .ZN(new_n319));
  INV_X1    g118(.A(G113gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n320), .A2(G120gat), .ZN(new_n321));
  INV_X1    g120(.A(G120gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n322), .A2(G113gat), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n319), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(G127gat), .ZN(new_n325));
  INV_X1    g124(.A(G134gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G127gat), .A2(G134gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n329), .A2(KEYINPUT67), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT67), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n331), .B1(new_n327), .B2(new_n328), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n324), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT68), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n334), .A2(new_n320), .A3(G120gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n335), .B1(new_n320), .B2(G120gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n323), .A2(new_n334), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n319), .B(new_n329), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(G155gat), .A2(G162gat), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT2), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(G155gat), .A2(G162gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  XOR2_X1   g143(.A(G141gat), .B(G148gat), .Z(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G141gat), .B(G148gat), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n343), .B1(new_n347), .B2(KEYINPUT2), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT74), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n340), .B(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n346), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n318), .B1(new_n339), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n351), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n353), .A2(KEYINPUT4), .A3(new_n333), .A4(new_n338), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n351), .A2(KEYINPUT3), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT3), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n346), .B(new_n358), .C1(new_n348), .C2(new_n350), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n339), .A3(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(KEYINPUT75), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT75), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n351), .A2(KEYINPUT3), .B1(new_n333), .B2(new_n338), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n362), .B1(new_n363), .B2(new_n359), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n355), .B(new_n356), .C1(new_n361), .C2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT5), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n366), .A2(KEYINPUT76), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n360), .A2(KEYINPUT75), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n363), .A2(new_n362), .A3(new_n359), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n367), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n371), .A2(new_n356), .A3(new_n355), .A4(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n339), .B(new_n351), .ZN(new_n375));
  INV_X1    g174(.A(new_n356), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(KEYINPUT5), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  XOR2_X1   g177(.A(G1gat), .B(G29gat), .Z(new_n379));
  XNOR2_X1  g178(.A(G57gat), .B(G85gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n381), .B(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n378), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT6), .ZN(new_n385));
  INV_X1    g184(.A(new_n377), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n386), .B1(new_n368), .B2(new_n373), .ZN(new_n387));
  INV_X1    g186(.A(new_n383), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n384), .A2(new_n385), .A3(new_n389), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n374), .A2(KEYINPUT6), .A3(new_n388), .A4(new_n377), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  XOR2_X1   g191(.A(G8gat), .B(G36gat), .Z(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(G64gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(new_n256), .ZN(new_n395));
  XNOR2_X1  g194(.A(G197gat), .B(G204gat), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT22), .ZN(new_n397));
  INV_X1    g196(.A(G211gat), .ZN(new_n398));
  INV_X1    g197(.A(G218gat), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  XOR2_X1   g200(.A(G211gat), .B(G218gat), .Z(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  NOR2_X1   g202(.A1(G169gat), .A2(G176gat), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT23), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G169gat), .A2(G176gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n411), .B1(G183gat), .B2(G190gat), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT25), .B1(new_n410), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT66), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT26), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n404), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n419));
  NOR3_X1   g218(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n418), .B(new_n419), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(G190gat), .ZN(new_n423));
  AND2_X1   g222(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n424));
  NOR2_X1   g223(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT28), .ZN(new_n427));
  XNOR2_X1  g226(.A(KEYINPUT27), .B(G183gat), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT28), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(new_n429), .A3(new_n423), .ZN(new_n430));
  NAND2_X1  g229(.A1(G183gat), .A2(G190gat), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n422), .A2(new_n427), .A3(new_n430), .A4(new_n431), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n406), .A2(new_n407), .B1(G169gat), .B2(G176gat), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT24), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT64), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT64), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n413), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n412), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n433), .B1(new_n439), .B2(KEYINPUT65), .ZN(new_n440));
  NOR2_X1   g239(.A1(G183gat), .A2(G190gat), .ZN(new_n441));
  AND2_X1   g240(.A1(G183gat), .A2(G190gat), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n441), .B1(new_n442), .B2(KEYINPUT24), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n431), .A2(new_n437), .A3(new_n434), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n437), .B1(new_n431), .B2(new_n434), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n443), .B(KEYINPUT65), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT25), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n415), .B(new_n432), .C1(new_n440), .C2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT29), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n449), .A2(new_n450), .B1(G226gat), .B2(G233gat), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n449), .A2(G226gat), .A3(G233gat), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n403), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n453), .ZN(new_n455));
  INV_X1    g254(.A(new_n403), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n455), .A2(new_n451), .A3(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n395), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n452), .A2(new_n403), .A3(new_n453), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n456), .B1(new_n455), .B2(new_n451), .ZN(new_n460));
  INV_X1    g259(.A(new_n395), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n458), .A2(new_n462), .A3(KEYINPUT30), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT30), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n459), .A2(new_n460), .A3(new_n464), .A4(new_n461), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n392), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(G227gat), .ZN(new_n468));
  INV_X1    g267(.A(G233gat), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n449), .A2(KEYINPUT69), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT65), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n474), .A2(new_n447), .A3(new_n433), .A4(new_n446), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT69), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n475), .A2(new_n476), .A3(new_n415), .A4(new_n432), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n471), .A2(new_n339), .A3(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n449), .A2(KEYINPUT69), .A3(new_n333), .A4(new_n338), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n470), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  AOI211_X1 g282(.A(new_n470), .B(new_n481), .C1(new_n478), .C2(new_n479), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n478), .A2(new_n470), .A3(new_n479), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT32), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT70), .ZN(new_n489));
  XNOR2_X1  g288(.A(G15gat), .B(G43gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(G71gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(G99gat), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT33), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n492), .B1(new_n487), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT70), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n487), .A2(new_n495), .A3(KEYINPUT32), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n489), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  OR2_X1    g296(.A1(new_n492), .A2(KEYINPUT71), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n492), .A2(KEYINPUT71), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(KEYINPUT33), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n487), .A2(KEYINPUT32), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT72), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n487), .A2(KEYINPUT72), .A3(KEYINPUT32), .A4(new_n500), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n486), .B1(new_n497), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G22gat), .B(G50gat), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n403), .B1(new_n450), .B2(new_n359), .ZN(new_n509));
  AND2_X1   g308(.A1(G228gat), .A2(G233gat), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n403), .A2(new_n450), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT78), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT3), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n403), .A2(KEYINPUT78), .A3(new_n450), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n511), .B1(new_n516), .B2(new_n353), .ZN(new_n517));
  XNOR2_X1  g316(.A(G78gat), .B(G106gat), .ZN(new_n518));
  XOR2_X1   g317(.A(new_n518), .B(KEYINPUT31), .Z(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n353), .B1(new_n512), .B2(new_n358), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n510), .B1(new_n521), .B2(new_n509), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n517), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n520), .B1(new_n517), .B2(new_n522), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n508), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n525), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n527), .A2(new_n507), .A3(new_n523), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n503), .A2(new_n504), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n489), .A2(new_n494), .A3(new_n496), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(new_n531), .A3(new_n485), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n506), .A2(new_n529), .A3(new_n532), .A4(KEYINPUT35), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n467), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n466), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n391), .A2(KEYINPUT80), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT80), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n387), .A2(new_n537), .A3(KEYINPUT6), .A4(new_n388), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n535), .B1(new_n539), .B2(new_n390), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n506), .A2(KEYINPUT81), .A3(new_n532), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT81), .B1(new_n506), .B2(new_n532), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n529), .B(new_n540), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT35), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n534), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n529), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n467), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT37), .B1(new_n454), .B2(new_n457), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT37), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n459), .A2(new_n460), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n548), .A2(new_n550), .A3(new_n395), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n551), .A2(KEYINPUT38), .ZN(new_n552));
  INV_X1    g351(.A(new_n462), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n551), .B1(new_n553), .B2(KEYINPUT38), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n539), .A2(new_n390), .A3(new_n552), .A4(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n355), .B1(new_n361), .B2(new_n364), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(new_n376), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n557), .B(KEYINPUT39), .C1(new_n376), .C2(new_n375), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT39), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n556), .A2(new_n559), .A3(new_n376), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n560), .A2(KEYINPUT79), .A3(new_n383), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT79), .B1(new_n560), .B2(new_n383), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n558), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT40), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n558), .B(KEYINPUT40), .C1(new_n561), .C2(new_n562), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n565), .A2(new_n535), .A3(new_n389), .A4(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n555), .A2(new_n567), .A3(new_n529), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT36), .ZN(new_n569));
  NOR3_X1   g368(.A1(new_n497), .A2(new_n486), .A3(new_n505), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n485), .B1(new_n530), .B2(new_n531), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n506), .A2(new_n532), .A3(KEYINPUT36), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n547), .A2(new_n568), .A3(new_n574), .ZN(new_n575));
  AOI211_X1 g374(.A(new_n253), .B(new_n317), .C1(new_n545), .C2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G134gat), .B(G162gat), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  AND2_X1   g377(.A1(G232gat), .A2(G233gat), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n303), .A2(new_n212), .B1(KEYINPUT41), .B2(new_n579), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n301), .A2(new_n302), .A3(new_n227), .A4(new_n214), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n578), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n579), .A2(KEYINPUT41), .ZN(new_n584));
  XNOR2_X1  g383(.A(G190gat), .B(G218gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n580), .A2(new_n578), .A3(new_n581), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n583), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n586), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n580), .A2(new_n578), .A3(new_n581), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n589), .B1(new_n590), .B2(new_n582), .ZN(new_n591));
  XNOR2_X1  g390(.A(G127gat), .B(G155gat), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n592), .B(KEYINPUT86), .Z(new_n593));
  INV_X1    g392(.A(G183gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT21), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n226), .B(new_n594), .C1(new_n595), .C2(new_n283), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n283), .A2(new_n595), .ZN(new_n597));
  OAI21_X1  g396(.A(G183gat), .B1(new_n597), .B2(new_n229), .ZN(new_n598));
  INV_X1    g397(.A(G231gat), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n599), .A2(new_n469), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n596), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n600), .B1(new_n596), .B2(new_n598), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n593), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n603), .ZN(new_n605));
  INV_X1    g404(.A(new_n593), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n605), .A2(new_n601), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n283), .A2(new_n595), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(new_n398), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n608), .B(new_n610), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n604), .A2(new_n607), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n611), .B1(new_n604), .B2(new_n607), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n588), .A2(new_n591), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT92), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n588), .A2(new_n591), .A3(new_n614), .A4(KEYINPUT92), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n576), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n392), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(KEYINPUT96), .B(G1gat), .Z(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(G1324gat));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n535), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(G8gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT97), .B(G8gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT16), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n620), .A2(new_n535), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT42), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT42), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT98), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT98), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n631), .A2(new_n636), .A3(new_n633), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(G1325gat));
  NOR2_X1   g437(.A1(new_n541), .A2(new_n542), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(G15gat), .B1(new_n620), .B2(new_n640), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n506), .A2(KEYINPUT36), .A3(new_n532), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT36), .B1(new_n506), .B2(new_n532), .ZN(new_n643));
  OAI21_X1  g442(.A(KEYINPUT99), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT99), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n572), .A2(new_n645), .A3(new_n573), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n620), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n641), .B1(new_n648), .B2(G15gat), .ZN(G1326gat));
  NAND2_X1  g448(.A1(new_n620), .A2(new_n546), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT43), .B(G22gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(G1327gat));
  AND2_X1   g451(.A1(new_n588), .A2(new_n591), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n653), .B1(new_n545), .B2(new_n575), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n317), .A2(new_n614), .A3(new_n253), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(G29gat), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n656), .A2(new_n657), .A3(new_n621), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT45), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n644), .A2(new_n646), .A3(new_n547), .A4(new_n568), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n545), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n588), .A2(new_n591), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT100), .B(KEYINPUT44), .Z(new_n663));
  NAND3_X1  g462(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n664), .B1(new_n665), .B2(new_n654), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n666), .A2(new_n655), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n621), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n659), .B1(new_n669), .B2(new_n657), .ZN(G1328gat));
  INV_X1    g469(.A(G36gat), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n656), .A2(new_n671), .A3(new_n535), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT101), .B(KEYINPUT46), .Z(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n667), .A2(new_n535), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n674), .B1(new_n676), .B2(new_n671), .ZN(G1329gat));
  INV_X1    g476(.A(G43gat), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n656), .A2(new_n678), .A3(new_n640), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n667), .A2(new_n647), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT103), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(G43gat), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n680), .A2(KEYINPUT103), .ZN(new_n683));
  OAI211_X1 g482(.A(KEYINPUT47), .B(new_n679), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT102), .B(KEYINPUT47), .Z(new_n685));
  AOI21_X1  g484(.A(new_n678), .B1(new_n667), .B2(new_n647), .ZN(new_n686));
  INV_X1    g485(.A(new_n679), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n684), .A2(new_n688), .ZN(G1330gat));
  INV_X1    g488(.A(KEYINPUT48), .ZN(new_n690));
  INV_X1    g489(.A(new_n663), .ZN(new_n691));
  AOI211_X1 g490(.A(new_n653), .B(new_n691), .C1(new_n545), .C2(new_n660), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n543), .A2(new_n544), .ZN(new_n693));
  INV_X1    g492(.A(new_n534), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n693), .A2(new_n575), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n665), .B1(new_n695), .B2(new_n662), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n546), .B(new_n655), .C1(new_n692), .C2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n666), .A2(KEYINPUT104), .A3(new_n546), .A4(new_n655), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n699), .A2(new_n700), .A3(G50gat), .ZN(new_n701));
  INV_X1    g500(.A(G50gat), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n656), .A2(new_n702), .A3(new_n546), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n690), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n697), .A2(G50gat), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n705), .A2(new_n690), .A3(new_n703), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT105), .B1(new_n704), .B2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT105), .ZN(new_n709));
  INV_X1    g508(.A(new_n703), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n702), .B1(new_n697), .B2(new_n698), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n710), .B1(new_n711), .B2(new_n700), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n709), .B(new_n706), .C1(new_n712), .C2(new_n690), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n708), .A2(new_n713), .ZN(G1331gat));
  INV_X1    g513(.A(new_n317), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n715), .B1(new_n545), .B2(new_n660), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n617), .A2(new_n618), .A3(new_n253), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n716), .A2(KEYINPUT106), .A3(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(KEYINPUT106), .B1(new_n716), .B2(new_n718), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n621), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(G57gat), .ZN(G1332gat));
  OAI21_X1  g523(.A(KEYINPUT107), .B1(new_n720), .B2(new_n721), .ZN(new_n725));
  INV_X1    g524(.A(new_n721), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n726), .A2(new_n727), .A3(new_n719), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n466), .B1(new_n725), .B2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n730));
  NAND2_X1  g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n730), .B1(new_n729), .B2(new_n731), .ZN(new_n733));
  OAI22_X1  g532(.A1(new_n732), .A2(new_n733), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n729), .A2(new_n731), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT108), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n737));
  NOR2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n734), .A2(new_n739), .ZN(G1333gat));
  INV_X1    g539(.A(KEYINPUT50), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n725), .A2(new_n728), .ZN(new_n742));
  INV_X1    g541(.A(new_n647), .ZN(new_n743));
  OAI21_X1  g542(.A(G71gat), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(G71gat), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n722), .A2(new_n745), .A3(new_n640), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n741), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n743), .B1(new_n725), .B2(new_n728), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n741), .B(new_n746), .C1(new_n748), .C2(new_n745), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n747), .A2(new_n750), .ZN(G1334gat));
  NOR2_X1   g550(.A1(new_n742), .A2(new_n529), .ZN(new_n752));
  XNOR2_X1  g551(.A(KEYINPUT109), .B(G78gat), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1335gat));
  AOI21_X1  g553(.A(new_n653), .B1(new_n545), .B2(new_n660), .ZN(new_n755));
  INV_X1    g554(.A(new_n614), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n253), .A2(new_n756), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(KEYINPUT110), .Z(new_n758));
  AND3_X1   g557(.A1(new_n755), .A2(KEYINPUT51), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT51), .B1(new_n755), .B2(new_n758), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n761), .A2(new_n715), .ZN(new_n762));
  AOI21_X1  g561(.A(G85gat), .B1(new_n762), .B2(new_n621), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n666), .A2(new_n317), .A3(new_n758), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT111), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n666), .A2(KEYINPUT111), .A3(new_n317), .A4(new_n758), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n769), .A2(new_n255), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n763), .B1(new_n770), .B2(new_n621), .ZN(G1336gat));
  OAI21_X1  g570(.A(G92gat), .B1(new_n764), .B2(new_n466), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n256), .B(new_n317), .C1(new_n759), .C2(new_n760), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n772), .B(new_n773), .C1(new_n466), .C2(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(new_n466), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n768), .A2(new_n535), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n776), .B1(new_n777), .B2(G92gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n775), .B1(new_n778), .B2(new_n773), .ZN(G1337gat));
  OAI21_X1  g578(.A(G99gat), .B1(new_n769), .B2(new_n743), .ZN(new_n780));
  INV_X1    g579(.A(G99gat), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n762), .A2(new_n781), .A3(new_n640), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(G1338gat));
  INV_X1    g582(.A(G106gat), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n784), .B1(new_n768), .B2(new_n546), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n317), .A2(new_n784), .A3(new_n546), .ZN(new_n786));
  XOR2_X1   g585(.A(new_n786), .B(KEYINPUT112), .Z(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(new_n759), .B2(new_n760), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(KEYINPUT53), .B1(new_n785), .B2(new_n789), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n666), .A2(new_n317), .A3(new_n546), .A4(new_n758), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT53), .B1(new_n791), .B2(G106gat), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n792), .A2(KEYINPUT113), .A3(new_n788), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT113), .B1(new_n792), .B2(new_n788), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n790), .A2(new_n795), .ZN(G1339gat));
  NOR2_X1   g595(.A1(new_n717), .A2(new_n317), .ZN(new_n797));
  INV_X1    g596(.A(new_n238), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n240), .A2(new_n243), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n231), .B1(new_n228), .B2(new_n230), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n801), .B1(new_n248), .B2(new_n249), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n317), .A2(new_n653), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n306), .A2(new_n289), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n298), .A2(new_n305), .A3(new_n288), .A4(new_n300), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n805), .A2(KEYINPUT54), .A3(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n306), .A2(new_n808), .A3(new_n289), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n807), .A2(KEYINPUT55), .A3(new_n313), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT114), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n313), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n813), .A2(new_n814), .A3(KEYINPUT55), .A4(new_n807), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  INV_X1    g616(.A(new_n807), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n817), .B1(new_n818), .B2(new_n812), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n653), .A2(new_n253), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n802), .A2(new_n821), .ZN(new_n822));
  OAI211_X1 g621(.A(KEYINPUT115), .B(new_n801), .C1(new_n248), .C2(new_n249), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n662), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n819), .A2(new_n820), .A3(new_n316), .A4(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n804), .B1(new_n816), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n797), .B1(new_n826), .B2(new_n756), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n392), .A2(new_n535), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n546), .A2(new_n570), .A3(new_n571), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n253), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n832), .A2(new_n320), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n639), .A2(new_n546), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n830), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(G113gat), .B1(new_n836), .B2(new_n253), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n834), .A2(new_n837), .ZN(G1340gat));
  NAND3_X1  g637(.A1(new_n832), .A2(new_n322), .A3(new_n317), .ZN(new_n839));
  OAI21_X1  g638(.A(G120gat), .B1(new_n836), .B2(new_n715), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(G1341gat));
  NAND2_X1  g640(.A1(new_n832), .A2(new_n614), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n325), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n830), .A2(G127gat), .A3(new_n614), .A4(new_n835), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n845), .B(new_n846), .ZN(G1342gat));
  AND3_X1   g646(.A1(new_n832), .A2(new_n326), .A3(new_n662), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT56), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(G134gat), .B1(new_n836), .B2(new_n653), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n848), .A2(new_n849), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(G1343gat));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n854), .B1(new_n827), .B2(new_n529), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n811), .A2(new_n815), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n824), .A2(new_n316), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n856), .A2(new_n857), .A3(new_n820), .A4(new_n819), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n614), .B1(new_n858), .B2(new_n804), .ZN(new_n859));
  OAI211_X1 g658(.A(KEYINPUT57), .B(new_n546), .C1(new_n859), .C2(new_n797), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n855), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  OR3_X1    g661(.A1(new_n647), .A2(KEYINPUT117), .A3(new_n829), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT117), .B1(new_n647), .B2(new_n829), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI211_X1 g664(.A(KEYINPUT118), .B(new_n854), .C1(new_n827), .C2(new_n529), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n862), .A2(new_n865), .A3(new_n833), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(G141gat), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n827), .A2(new_n529), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n647), .A2(new_n829), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OR3_X1    g670(.A1(new_n871), .A2(G141gat), .A3(new_n253), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT58), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT58), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n868), .A2(new_n875), .A3(new_n872), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(G1344gat));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n826), .A2(new_n756), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n619), .A2(KEYINPUT119), .A3(new_n253), .A4(new_n715), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT119), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n881), .B1(new_n717), .B2(new_n317), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n529), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n878), .B1(new_n884), .B2(KEYINPUT57), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n880), .A2(new_n882), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n546), .B1(new_n859), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(KEYINPUT120), .A3(new_n854), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n885), .A2(new_n860), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n715), .B1(new_n863), .B2(new_n864), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n862), .A2(new_n893), .A3(new_n866), .A4(new_n890), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n871), .A2(new_n715), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(new_n893), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n892), .B(new_n894), .C1(G148gat), .C2(new_n896), .ZN(G1345gat));
  NAND3_X1  g696(.A1(new_n862), .A2(new_n865), .A3(new_n866), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n614), .A2(G155gat), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n871), .A2(new_n756), .ZN(new_n900));
  OAI22_X1  g699(.A1(new_n898), .A2(new_n899), .B1(G155gat), .B2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n901), .B(new_n902), .ZN(G1346gat));
  INV_X1    g702(.A(G162gat), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n898), .A2(new_n904), .A3(new_n653), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n869), .A2(new_n662), .A3(new_n870), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n905), .B1(new_n904), .B2(new_n906), .ZN(G1347gat));
  INV_X1    g706(.A(new_n827), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n621), .A2(new_n466), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT123), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n908), .A2(new_n835), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(G169gat), .B1(new_n911), .B2(new_n253), .ZN(new_n912));
  INV_X1    g711(.A(G169gat), .ZN(new_n913));
  AND4_X1   g712(.A1(new_n913), .A2(new_n908), .A3(new_n831), .A4(new_n909), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n914), .A2(new_n915), .A3(new_n833), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n914), .B2(new_n833), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n912), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g719(.A(KEYINPUT124), .B(new_n912), .C1(new_n916), .C2(new_n917), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1348gat));
  AND3_X1   g721(.A1(new_n908), .A2(new_n831), .A3(new_n909), .ZN(new_n923));
  AOI21_X1  g722(.A(G176gat), .B1(new_n923), .B2(new_n317), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n911), .A2(new_n311), .A3(new_n715), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(G1349gat));
  NAND3_X1  g725(.A1(new_n923), .A2(new_n614), .A3(new_n428), .ZN(new_n927));
  OAI21_X1  g726(.A(G183gat), .B1(new_n911), .B2(new_n756), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT60), .ZN(G1350gat));
  OR2_X1    g729(.A1(new_n911), .A2(new_n653), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(G190gat), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT125), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT125), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n931), .A2(new_n934), .A3(G190gat), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n933), .A2(KEYINPUT61), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n923), .A2(new_n423), .A3(new_n662), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT61), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n932), .A2(KEYINPUT125), .A3(new_n938), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(G1351gat));
  NAND2_X1  g739(.A1(new_n910), .A2(new_n743), .ZN(new_n941));
  XOR2_X1   g740(.A(new_n941), .B(KEYINPUT126), .Z(new_n942));
  NAND3_X1  g741(.A1(new_n889), .A2(new_n833), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(G197gat), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n647), .A2(new_n621), .A3(new_n466), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n869), .A2(new_n945), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n946), .A2(G197gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n944), .B1(new_n253), .B2(new_n947), .ZN(G1352gat));
  INV_X1    g747(.A(new_n946), .ZN(new_n949));
  XNOR2_X1  g748(.A(KEYINPUT127), .B(G204gat), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n949), .A2(new_n317), .A3(new_n951), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n952), .A2(KEYINPUT62), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(KEYINPUT62), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n889), .A2(new_n317), .A3(new_n942), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n953), .B(new_n954), .C1(new_n955), .C2(new_n951), .ZN(G1353gat));
  NAND3_X1  g755(.A1(new_n949), .A2(new_n398), .A3(new_n614), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n889), .A2(new_n614), .A3(new_n942), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n958), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT63), .B1(new_n958), .B2(G211gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(G1354gat));
  NAND3_X1  g760(.A1(new_n949), .A2(new_n399), .A3(new_n662), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n889), .A2(new_n662), .A3(new_n942), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n962), .B1(new_n963), .B2(new_n399), .ZN(G1355gat));
endmodule


