

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U549 ( .A1(n524), .A2(G2104), .ZN(n893) );
  NOR2_X1 U550 ( .A1(G2104), .A2(n524), .ZN(n902) );
  BUF_X1 U551 ( .A(n720), .Z(G164) );
  XNOR2_X1 U552 ( .A(n758), .B(KEYINPUT29), .ZN(n759) );
  NOR2_X2 U553 ( .A1(G651), .A2(n639), .ZN(n656) );
  INV_X1 U554 ( .A(n519), .ZN(n895) );
  INV_X1 U555 ( .A(KEYINPUT23), .ZN(n520) );
  AND2_X1 U556 ( .A1(n978), .A2(n517), .ZN(n516) );
  OR2_X1 U557 ( .A1(n792), .A2(n803), .ZN(n517) );
  INV_X1 U558 ( .A(KEYINPUT26), .ZN(n733) );
  NAND2_X1 U559 ( .A1(n763), .A2(n762), .ZN(n776) );
  AND2_X1 U560 ( .A1(n765), .A2(n764), .ZN(n766) );
  INV_X1 U561 ( .A(G2105), .ZN(n524) );
  XNOR2_X1 U562 ( .A(n521), .B(n520), .ZN(n522) );
  NOR2_X2 U563 ( .A1(G2104), .A2(G2105), .ZN(n518) );
  XOR2_X1 U564 ( .A(KEYINPUT17), .B(n518), .Z(n531) );
  INV_X1 U565 ( .A(n531), .ZN(n519) );
  NAND2_X1 U566 ( .A1(n895), .A2(G137), .ZN(n523) );
  NAND2_X1 U567 ( .A1(G101), .A2(n893), .ZN(n521) );
  NAND2_X1 U568 ( .A1(n523), .A2(n522), .ZN(n528) );
  AND2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n899) );
  NAND2_X1 U570 ( .A1(G113), .A2(n899), .ZN(n526) );
  NAND2_X1 U571 ( .A1(G125), .A2(n902), .ZN(n525) );
  NAND2_X1 U572 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X2 U573 ( .A1(n528), .A2(n527), .ZN(G160) );
  NAND2_X1 U574 ( .A1(G102), .A2(n893), .ZN(n530) );
  NAND2_X1 U575 ( .A1(G114), .A2(n899), .ZN(n529) );
  AND2_X1 U576 ( .A1(n530), .A2(n529), .ZN(n535) );
  AND2_X1 U577 ( .A1(n531), .A2(G138), .ZN(n533) );
  INV_X1 U578 ( .A(KEYINPUT90), .ZN(n532) );
  XNOR2_X1 U579 ( .A(n533), .B(n532), .ZN(n534) );
  NAND2_X1 U580 ( .A1(n535), .A2(n534), .ZN(n537) );
  AND2_X1 U581 ( .A1(G126), .A2(n902), .ZN(n536) );
  NOR2_X1 U582 ( .A1(n537), .A2(n536), .ZN(n539) );
  INV_X1 U583 ( .A(KEYINPUT91), .ZN(n538) );
  XNOR2_X1 U584 ( .A(n539), .B(n538), .ZN(n720) );
  XOR2_X1 U585 ( .A(KEYINPUT81), .B(KEYINPUT18), .Z(n542) );
  NAND2_X1 U586 ( .A1(G123), .A2(n902), .ZN(n541) );
  XNOR2_X1 U587 ( .A(n542), .B(n541), .ZN(n549) );
  NAND2_X1 U588 ( .A1(G99), .A2(n893), .ZN(n544) );
  NAND2_X1 U589 ( .A1(G135), .A2(n895), .ZN(n543) );
  NAND2_X1 U590 ( .A1(n544), .A2(n543), .ZN(n547) );
  NAND2_X1 U591 ( .A1(n899), .A2(G111), .ZN(n545) );
  XOR2_X1 U592 ( .A(KEYINPUT82), .B(n545), .Z(n546) );
  NOR2_X1 U593 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U594 ( .A1(n549), .A2(n548), .ZN(n961) );
  XNOR2_X1 U595 ( .A(G2096), .B(n961), .ZN(n550) );
  OR2_X1 U596 ( .A1(G2100), .A2(n550), .ZN(G156) );
  INV_X1 U597 ( .A(G57), .ZN(G237) );
  INV_X1 U598 ( .A(G120), .ZN(G236) );
  INV_X1 U599 ( .A(G108), .ZN(G238) );
  NOR2_X1 U600 ( .A1(G651), .A2(G543), .ZN(n653) );
  NAND2_X1 U601 ( .A1(G88), .A2(n653), .ZN(n552) );
  XOR2_X1 U602 ( .A(KEYINPUT0), .B(G543), .Z(n639) );
  INV_X1 U603 ( .A(G651), .ZN(n553) );
  NOR2_X1 U604 ( .A1(n639), .A2(n553), .ZN(n650) );
  NAND2_X1 U605 ( .A1(G75), .A2(n650), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n552), .A2(n551), .ZN(n558) );
  NAND2_X1 U607 ( .A1(G50), .A2(n656), .ZN(n556) );
  NOR2_X1 U608 ( .A1(G543), .A2(n553), .ZN(n554) );
  XOR2_X1 U609 ( .A(KEYINPUT1), .B(n554), .Z(n652) );
  NAND2_X1 U610 ( .A1(G62), .A2(n652), .ZN(n555) );
  NAND2_X1 U611 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U612 ( .A1(n558), .A2(n557), .ZN(G166) );
  NAND2_X1 U613 ( .A1(G90), .A2(n653), .ZN(n560) );
  NAND2_X1 U614 ( .A1(G77), .A2(n650), .ZN(n559) );
  NAND2_X1 U615 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U616 ( .A(n561), .B(KEYINPUT9), .ZN(n563) );
  NAND2_X1 U617 ( .A1(G64), .A2(n652), .ZN(n562) );
  NAND2_X1 U618 ( .A1(n563), .A2(n562), .ZN(n566) );
  NAND2_X1 U619 ( .A1(n656), .A2(G52), .ZN(n564) );
  XOR2_X1 U620 ( .A(KEYINPUT66), .B(n564), .Z(n565) );
  NOR2_X1 U621 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U622 ( .A(KEYINPUT67), .B(n567), .Z(G171) );
  NAND2_X1 U623 ( .A1(G76), .A2(n650), .ZN(n571) );
  XOR2_X1 U624 ( .A(KEYINPUT4), .B(KEYINPUT77), .Z(n569) );
  NAND2_X1 U625 ( .A1(G89), .A2(n653), .ZN(n568) );
  XNOR2_X1 U626 ( .A(n569), .B(n568), .ZN(n570) );
  NAND2_X1 U627 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U628 ( .A(n572), .B(KEYINPUT78), .ZN(n573) );
  XNOR2_X1 U629 ( .A(KEYINPUT5), .B(n573), .ZN(n578) );
  NAND2_X1 U630 ( .A1(G51), .A2(n656), .ZN(n575) );
  NAND2_X1 U631 ( .A1(G63), .A2(n652), .ZN(n574) );
  NAND2_X1 U632 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U633 ( .A(KEYINPUT6), .B(n576), .Z(n577) );
  NAND2_X1 U634 ( .A1(n578), .A2(n577), .ZN(n580) );
  XOR2_X1 U635 ( .A(KEYINPUT7), .B(KEYINPUT79), .Z(n579) );
  XNOR2_X1 U636 ( .A(n580), .B(n579), .ZN(G168) );
  XOR2_X1 U637 ( .A(G168), .B(KEYINPUT8), .Z(n581) );
  XNOR2_X1 U638 ( .A(KEYINPUT80), .B(n581), .ZN(G286) );
  NAND2_X1 U639 ( .A1(G94), .A2(G452), .ZN(n582) );
  XOR2_X1 U640 ( .A(KEYINPUT68), .B(n582), .Z(G173) );
  NAND2_X1 U641 ( .A1(G7), .A2(G661), .ZN(n583) );
  XNOR2_X1 U642 ( .A(n583), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U643 ( .A(G223), .ZN(n831) );
  NAND2_X1 U644 ( .A1(n831), .A2(G567), .ZN(n584) );
  XOR2_X1 U645 ( .A(KEYINPUT11), .B(n584), .Z(G234) );
  XNOR2_X1 U646 ( .A(KEYINPUT72), .B(KEYINPUT12), .ZN(n586) );
  NAND2_X1 U647 ( .A1(n653), .A2(G81), .ZN(n585) );
  XNOR2_X1 U648 ( .A(n586), .B(n585), .ZN(n588) );
  NAND2_X1 U649 ( .A1(G68), .A2(n650), .ZN(n587) );
  NAND2_X1 U650 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U651 ( .A(KEYINPUT13), .B(n589), .Z(n592) );
  NAND2_X1 U652 ( .A1(n652), .A2(G56), .ZN(n590) );
  XOR2_X1 U653 ( .A(KEYINPUT14), .B(n590), .Z(n591) );
  NOR2_X1 U654 ( .A1(n592), .A2(n591), .ZN(n594) );
  NAND2_X1 U655 ( .A1(n656), .A2(G43), .ZN(n593) );
  NAND2_X1 U656 ( .A1(n594), .A2(n593), .ZN(n984) );
  INV_X1 U657 ( .A(G860), .ZN(n627) );
  OR2_X1 U658 ( .A1(n984), .A2(n627), .ZN(G153) );
  INV_X1 U659 ( .A(G171), .ZN(G301) );
  NAND2_X1 U660 ( .A1(G66), .A2(n652), .ZN(n601) );
  NAND2_X1 U661 ( .A1(G92), .A2(n653), .ZN(n596) );
  NAND2_X1 U662 ( .A1(G79), .A2(n650), .ZN(n595) );
  NAND2_X1 U663 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U664 ( .A1(G54), .A2(n656), .ZN(n597) );
  XNOR2_X1 U665 ( .A(KEYINPUT73), .B(n597), .ZN(n598) );
  NOR2_X1 U666 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U667 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U668 ( .A(n602), .B(KEYINPUT15), .ZN(n603) );
  XNOR2_X2 U669 ( .A(KEYINPUT74), .B(n603), .ZN(n995) );
  NOR2_X1 U670 ( .A1(G868), .A2(n995), .ZN(n604) );
  XNOR2_X1 U671 ( .A(n604), .B(KEYINPUT75), .ZN(n606) );
  NAND2_X1 U672 ( .A1(G868), .A2(G301), .ZN(n605) );
  NAND2_X1 U673 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U674 ( .A(KEYINPUT76), .B(n607), .ZN(G284) );
  NAND2_X1 U675 ( .A1(G78), .A2(n650), .ZN(n608) );
  XNOR2_X1 U676 ( .A(n608), .B(KEYINPUT70), .ZN(n610) );
  NAND2_X1 U677 ( .A1(n652), .A2(G65), .ZN(n609) );
  NAND2_X1 U678 ( .A1(n610), .A2(n609), .ZN(n613) );
  NAND2_X1 U679 ( .A1(G91), .A2(n653), .ZN(n611) );
  XNOR2_X1 U680 ( .A(KEYINPUT69), .B(n611), .ZN(n612) );
  NOR2_X1 U681 ( .A1(n613), .A2(n612), .ZN(n616) );
  NAND2_X1 U682 ( .A1(G53), .A2(n656), .ZN(n614) );
  XOR2_X1 U683 ( .A(KEYINPUT71), .B(n614), .Z(n615) );
  NAND2_X1 U684 ( .A1(n616), .A2(n615), .ZN(G299) );
  NAND2_X1 U685 ( .A1(G868), .A2(G286), .ZN(n619) );
  INV_X1 U686 ( .A(G868), .ZN(n617) );
  NAND2_X1 U687 ( .A1(G299), .A2(n617), .ZN(n618) );
  NAND2_X1 U688 ( .A1(n619), .A2(n618), .ZN(G297) );
  NAND2_X1 U689 ( .A1(n627), .A2(G559), .ZN(n620) );
  NAND2_X1 U690 ( .A1(n620), .A2(n995), .ZN(n621) );
  XNOR2_X1 U691 ( .A(n621), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U692 ( .A1(G868), .A2(n984), .ZN(n624) );
  NAND2_X1 U693 ( .A1(n995), .A2(G868), .ZN(n622) );
  NOR2_X1 U694 ( .A1(G559), .A2(n622), .ZN(n623) );
  NOR2_X1 U695 ( .A1(n624), .A2(n623), .ZN(G282) );
  XNOR2_X1 U696 ( .A(n984), .B(KEYINPUT83), .ZN(n626) );
  NAND2_X1 U697 ( .A1(n995), .A2(G559), .ZN(n625) );
  XNOR2_X1 U698 ( .A(n626), .B(n625), .ZN(n667) );
  NAND2_X1 U699 ( .A1(n627), .A2(n667), .ZN(n635) );
  NAND2_X1 U700 ( .A1(G93), .A2(n653), .ZN(n629) );
  NAND2_X1 U701 ( .A1(G80), .A2(n650), .ZN(n628) );
  NAND2_X1 U702 ( .A1(n629), .A2(n628), .ZN(n634) );
  NAND2_X1 U703 ( .A1(n656), .A2(G55), .ZN(n630) );
  XNOR2_X1 U704 ( .A(n630), .B(KEYINPUT84), .ZN(n632) );
  NAND2_X1 U705 ( .A1(G67), .A2(n652), .ZN(n631) );
  NAND2_X1 U706 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U707 ( .A1(n634), .A2(n633), .ZN(n669) );
  XOR2_X1 U708 ( .A(n635), .B(n669), .Z(G145) );
  NAND2_X1 U709 ( .A1(G49), .A2(n656), .ZN(n637) );
  NAND2_X1 U710 ( .A1(G74), .A2(G651), .ZN(n636) );
  NAND2_X1 U711 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U712 ( .A1(n652), .A2(n638), .ZN(n641) );
  NAND2_X1 U713 ( .A1(n639), .A2(G87), .ZN(n640) );
  NAND2_X1 U714 ( .A1(n641), .A2(n640), .ZN(G288) );
  NAND2_X1 U715 ( .A1(G61), .A2(n652), .ZN(n643) );
  NAND2_X1 U716 ( .A1(G86), .A2(n653), .ZN(n642) );
  NAND2_X1 U717 ( .A1(n643), .A2(n642), .ZN(n646) );
  NAND2_X1 U718 ( .A1(n650), .A2(G73), .ZN(n644) );
  XOR2_X1 U719 ( .A(KEYINPUT2), .B(n644), .Z(n645) );
  NOR2_X1 U720 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U721 ( .A(KEYINPUT85), .B(n647), .Z(n649) );
  NAND2_X1 U722 ( .A1(n656), .A2(G48), .ZN(n648) );
  NAND2_X1 U723 ( .A1(n649), .A2(n648), .ZN(G305) );
  NAND2_X1 U724 ( .A1(G72), .A2(n650), .ZN(n651) );
  XNOR2_X1 U725 ( .A(n651), .B(KEYINPUT64), .ZN(n661) );
  NAND2_X1 U726 ( .A1(G60), .A2(n652), .ZN(n655) );
  NAND2_X1 U727 ( .A1(G85), .A2(n653), .ZN(n654) );
  NAND2_X1 U728 ( .A1(n655), .A2(n654), .ZN(n659) );
  NAND2_X1 U729 ( .A1(G47), .A2(n656), .ZN(n657) );
  XNOR2_X1 U730 ( .A(KEYINPUT65), .B(n657), .ZN(n658) );
  NOR2_X1 U731 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U732 ( .A1(n661), .A2(n660), .ZN(G290) );
  XNOR2_X1 U733 ( .A(G166), .B(KEYINPUT19), .ZN(n666) );
  XNOR2_X1 U734 ( .A(n669), .B(G288), .ZN(n664) );
  XNOR2_X1 U735 ( .A(G299), .B(G305), .ZN(n662) );
  XNOR2_X1 U736 ( .A(n662), .B(G290), .ZN(n663) );
  XNOR2_X1 U737 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U738 ( .A(n666), .B(n665), .ZN(n912) );
  XNOR2_X1 U739 ( .A(n667), .B(n912), .ZN(n668) );
  NAND2_X1 U740 ( .A1(n668), .A2(G868), .ZN(n671) );
  OR2_X1 U741 ( .A1(G868), .A2(n669), .ZN(n670) );
  NAND2_X1 U742 ( .A1(n671), .A2(n670), .ZN(G295) );
  NAND2_X1 U743 ( .A1(G2078), .A2(G2084), .ZN(n673) );
  XOR2_X1 U744 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n672) );
  XNOR2_X1 U745 ( .A(n673), .B(n672), .ZN(n674) );
  NAND2_X1 U746 ( .A1(G2090), .A2(n674), .ZN(n675) );
  XNOR2_X1 U747 ( .A(KEYINPUT21), .B(n675), .ZN(n676) );
  NAND2_X1 U748 ( .A1(n676), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U749 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U750 ( .A1(G238), .A2(G236), .ZN(n677) );
  NAND2_X1 U751 ( .A1(G69), .A2(n677), .ZN(n678) );
  NOR2_X1 U752 ( .A1(n678), .A2(G237), .ZN(n679) );
  XNOR2_X1 U753 ( .A(n679), .B(KEYINPUT89), .ZN(n836) );
  NAND2_X1 U754 ( .A1(n836), .A2(G567), .ZN(n686) );
  XOR2_X1 U755 ( .A(KEYINPUT87), .B(KEYINPUT22), .Z(n681) );
  NAND2_X1 U756 ( .A1(G132), .A2(G82), .ZN(n680) );
  XNOR2_X1 U757 ( .A(n681), .B(n680), .ZN(n682) );
  NOR2_X1 U758 ( .A1(n682), .A2(G218), .ZN(n683) );
  XNOR2_X1 U759 ( .A(KEYINPUT88), .B(n683), .ZN(n684) );
  NAND2_X1 U760 ( .A1(n684), .A2(G96), .ZN(n837) );
  NAND2_X1 U761 ( .A1(n837), .A2(G2106), .ZN(n685) );
  NAND2_X1 U762 ( .A1(n686), .A2(n685), .ZN(n921) );
  NAND2_X1 U763 ( .A1(G661), .A2(G483), .ZN(n687) );
  NOR2_X1 U764 ( .A1(n921), .A2(n687), .ZN(n834) );
  NAND2_X1 U765 ( .A1(n834), .A2(G36), .ZN(G176) );
  INV_X1 U766 ( .A(G166), .ZN(G303) );
  NAND2_X1 U767 ( .A1(n893), .A2(G95), .ZN(n688) );
  XNOR2_X1 U768 ( .A(n688), .B(KEYINPUT94), .ZN(n690) );
  NAND2_X1 U769 ( .A1(G119), .A2(n902), .ZN(n689) );
  NAND2_X1 U770 ( .A1(n690), .A2(n689), .ZN(n694) );
  NAND2_X1 U771 ( .A1(G131), .A2(n895), .ZN(n692) );
  NAND2_X1 U772 ( .A1(G107), .A2(n899), .ZN(n691) );
  NAND2_X1 U773 ( .A1(n692), .A2(n691), .ZN(n693) );
  OR2_X1 U774 ( .A1(n694), .A2(n693), .ZN(n885) );
  AND2_X1 U775 ( .A1(n885), .A2(G1991), .ZN(n703) );
  NAND2_X1 U776 ( .A1(G141), .A2(n895), .ZN(n696) );
  NAND2_X1 U777 ( .A1(G129), .A2(n902), .ZN(n695) );
  NAND2_X1 U778 ( .A1(n696), .A2(n695), .ZN(n699) );
  NAND2_X1 U779 ( .A1(n893), .A2(G105), .ZN(n697) );
  XOR2_X1 U780 ( .A(KEYINPUT38), .B(n697), .Z(n698) );
  NOR2_X1 U781 ( .A1(n699), .A2(n698), .ZN(n701) );
  NAND2_X1 U782 ( .A1(n899), .A2(G117), .ZN(n700) );
  NAND2_X1 U783 ( .A1(n701), .A2(n700), .ZN(n886) );
  AND2_X1 U784 ( .A1(n886), .A2(G1996), .ZN(n702) );
  NOR2_X1 U785 ( .A1(n703), .A2(n702), .ZN(n948) );
  NOR2_X1 U786 ( .A1(G164), .A2(G1384), .ZN(n704) );
  NAND2_X1 U787 ( .A1(G160), .A2(G40), .ZN(n717) );
  NOR2_X1 U788 ( .A1(n704), .A2(n717), .ZN(n826) );
  INV_X1 U789 ( .A(n826), .ZN(n705) );
  NOR2_X1 U790 ( .A1(n948), .A2(n705), .ZN(n816) );
  INV_X1 U791 ( .A(n816), .ZN(n716) );
  XNOR2_X1 U792 ( .A(G2067), .B(KEYINPUT37), .ZN(n822) );
  NAND2_X1 U793 ( .A1(G104), .A2(n893), .ZN(n707) );
  NAND2_X1 U794 ( .A1(G140), .A2(n895), .ZN(n706) );
  NAND2_X1 U795 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U796 ( .A(KEYINPUT34), .B(n708), .ZN(n714) );
  NAND2_X1 U797 ( .A1(G116), .A2(n899), .ZN(n710) );
  NAND2_X1 U798 ( .A1(G128), .A2(n902), .ZN(n709) );
  NAND2_X1 U799 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U800 ( .A(KEYINPUT93), .B(n711), .ZN(n712) );
  XNOR2_X1 U801 ( .A(KEYINPUT35), .B(n712), .ZN(n713) );
  NOR2_X1 U802 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U803 ( .A(KEYINPUT36), .B(n715), .ZN(n892) );
  NOR2_X1 U804 ( .A1(n822), .A2(n892), .ZN(n963) );
  NAND2_X1 U805 ( .A1(n826), .A2(n963), .ZN(n820) );
  NAND2_X1 U806 ( .A1(n716), .A2(n820), .ZN(n810) );
  INV_X1 U807 ( .A(n717), .ZN(n719) );
  INV_X1 U808 ( .A(G1384), .ZN(n718) );
  NAND2_X1 U809 ( .A1(n719), .A2(n718), .ZN(n721) );
  OR2_X4 U810 ( .A1(n721), .A2(n720), .ZN(n768) );
  NOR2_X1 U811 ( .A1(G2084), .A2(n768), .ZN(n722) );
  NAND2_X1 U812 ( .A1(G8), .A2(n722), .ZN(n767) );
  NAND2_X1 U813 ( .A1(G8), .A2(n768), .ZN(n803) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n803), .ZN(n723) );
  INV_X1 U815 ( .A(n723), .ZN(n765) );
  NOR2_X1 U816 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U817 ( .A1(G8), .A2(n724), .ZN(n725) );
  XNOR2_X1 U818 ( .A(KEYINPUT30), .B(n725), .ZN(n726) );
  NOR2_X1 U819 ( .A1(G168), .A2(n726), .ZN(n730) );
  INV_X1 U820 ( .A(G1961), .ZN(n922) );
  NAND2_X1 U821 ( .A1(n768), .A2(n922), .ZN(n728) );
  INV_X1 U822 ( .A(n768), .ZN(n738) );
  XNOR2_X1 U823 ( .A(KEYINPUT25), .B(G2078), .ZN(n1006) );
  NAND2_X1 U824 ( .A1(n738), .A2(n1006), .ZN(n727) );
  NAND2_X1 U825 ( .A1(n728), .A2(n727), .ZN(n761) );
  NOR2_X1 U826 ( .A1(G171), .A2(n761), .ZN(n729) );
  NOR2_X1 U827 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U828 ( .A(KEYINPUT31), .B(n731), .Z(n774) );
  INV_X1 U829 ( .A(G1996), .ZN(n732) );
  NOR2_X2 U830 ( .A1(n768), .A2(n732), .ZN(n734) );
  XNOR2_X1 U831 ( .A(n734), .B(n733), .ZN(n736) );
  NAND2_X1 U832 ( .A1(n768), .A2(G1341), .ZN(n735) );
  NAND2_X1 U833 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X2 U834 ( .A1(n737), .A2(n984), .ZN(n744) );
  NAND2_X1 U835 ( .A1(n744), .A2(n995), .ZN(n742) );
  NOR2_X1 U836 ( .A1(G2067), .A2(n768), .ZN(n740) );
  NOR2_X1 U837 ( .A1(n738), .A2(G1348), .ZN(n739) );
  NOR2_X1 U838 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U839 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U840 ( .A(n743), .B(KEYINPUT97), .ZN(n746) );
  NOR2_X1 U841 ( .A1(n995), .A2(n744), .ZN(n745) );
  NOR2_X1 U842 ( .A1(n746), .A2(n745), .ZN(n752) );
  INV_X1 U843 ( .A(n768), .ZN(n747) );
  NAND2_X1 U844 ( .A1(n747), .A2(G2072), .ZN(n748) );
  XOR2_X1 U845 ( .A(KEYINPUT27), .B(n748), .Z(n750) );
  NAND2_X1 U846 ( .A1(G1956), .A2(n768), .ZN(n749) );
  NAND2_X1 U847 ( .A1(n750), .A2(n749), .ZN(n754) );
  NOR2_X1 U848 ( .A1(G299), .A2(n754), .ZN(n751) );
  NOR2_X1 U849 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U850 ( .A(KEYINPUT98), .B(n753), .ZN(n757) );
  NAND2_X1 U851 ( .A1(G299), .A2(n754), .ZN(n755) );
  XOR2_X1 U852 ( .A(n755), .B(KEYINPUT28), .Z(n756) );
  NOR2_X1 U853 ( .A1(n757), .A2(n756), .ZN(n760) );
  INV_X1 U854 ( .A(KEYINPUT99), .ZN(n758) );
  XNOR2_X1 U855 ( .A(n760), .B(n759), .ZN(n763) );
  NAND2_X1 U856 ( .A1(G171), .A2(n761), .ZN(n762) );
  NAND2_X1 U857 ( .A1(n774), .A2(n776), .ZN(n764) );
  NAND2_X1 U858 ( .A1(n767), .A2(n766), .ZN(n783) );
  INV_X1 U859 ( .A(G8), .ZN(n773) );
  NOR2_X1 U860 ( .A1(G1971), .A2(n803), .ZN(n770) );
  NOR2_X1 U861 ( .A1(G2090), .A2(n768), .ZN(n769) );
  NOR2_X1 U862 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U863 ( .A1(n771), .A2(G303), .ZN(n772) );
  OR2_X1 U864 ( .A1(n773), .A2(n772), .ZN(n777) );
  AND2_X1 U865 ( .A1(n774), .A2(n777), .ZN(n775) );
  NAND2_X1 U866 ( .A1(n776), .A2(n775), .ZN(n780) );
  INV_X1 U867 ( .A(n777), .ZN(n778) );
  OR2_X1 U868 ( .A1(n778), .A2(G286), .ZN(n779) );
  NAND2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U870 ( .A(n781), .B(KEYINPUT32), .ZN(n782) );
  NAND2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n795) );
  NOR2_X1 U872 ( .A1(G1976), .A2(G288), .ZN(n992) );
  NOR2_X1 U873 ( .A1(G1971), .A2(G303), .ZN(n784) );
  NOR2_X1 U874 ( .A1(n992), .A2(n784), .ZN(n785) );
  NAND2_X1 U875 ( .A1(n795), .A2(n785), .ZN(n786) );
  NAND2_X1 U876 ( .A1(G1976), .A2(G288), .ZN(n996) );
  NAND2_X1 U877 ( .A1(n786), .A2(n996), .ZN(n787) );
  XNOR2_X1 U878 ( .A(KEYINPUT100), .B(n787), .ZN(n788) );
  NOR2_X1 U879 ( .A1(n788), .A2(n803), .ZN(n789) );
  INV_X1 U880 ( .A(n789), .ZN(n791) );
  INV_X1 U881 ( .A(KEYINPUT33), .ZN(n790) );
  NAND2_X1 U882 ( .A1(n791), .A2(n790), .ZN(n793) );
  XOR2_X1 U883 ( .A(G1981), .B(G305), .Z(n978) );
  NAND2_X1 U884 ( .A1(n992), .A2(KEYINPUT33), .ZN(n792) );
  NAND2_X1 U885 ( .A1(n793), .A2(n516), .ZN(n794) );
  XNOR2_X1 U886 ( .A(KEYINPUT101), .B(n794), .ZN(n808) );
  BUF_X1 U887 ( .A(n795), .Z(n798) );
  NOR2_X1 U888 ( .A1(G2090), .A2(G303), .ZN(n796) );
  NAND2_X1 U889 ( .A1(G8), .A2(n796), .ZN(n797) );
  NAND2_X1 U890 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U891 ( .A1(n803), .A2(n799), .ZN(n806) );
  NOR2_X1 U892 ( .A1(G1981), .A2(G305), .ZN(n800) );
  XNOR2_X1 U893 ( .A(n800), .B(KEYINPUT24), .ZN(n801) );
  XNOR2_X1 U894 ( .A(n801), .B(KEYINPUT95), .ZN(n802) );
  NOR2_X1 U895 ( .A1(n803), .A2(n802), .ZN(n804) );
  XOR2_X1 U896 ( .A(KEYINPUT96), .B(n804), .Z(n805) );
  NAND2_X1 U897 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U898 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U899 ( .A1(n810), .A2(n809), .ZN(n813) );
  XNOR2_X1 U900 ( .A(KEYINPUT92), .B(G1986), .ZN(n811) );
  XNOR2_X1 U901 ( .A(n811), .B(G290), .ZN(n991) );
  NAND2_X1 U902 ( .A1(n826), .A2(n991), .ZN(n812) );
  NAND2_X1 U903 ( .A1(n813), .A2(n812), .ZN(n829) );
  NOR2_X1 U904 ( .A1(G1996), .A2(n886), .ZN(n954) );
  NOR2_X1 U905 ( .A1(G1986), .A2(G290), .ZN(n814) );
  NOR2_X1 U906 ( .A1(G1991), .A2(n885), .ZN(n960) );
  NOR2_X1 U907 ( .A1(n814), .A2(n960), .ZN(n815) );
  NOR2_X1 U908 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U909 ( .A(n817), .B(KEYINPUT102), .ZN(n818) );
  NOR2_X1 U910 ( .A1(n954), .A2(n818), .ZN(n819) );
  XNOR2_X1 U911 ( .A(KEYINPUT39), .B(n819), .ZN(n821) );
  NAND2_X1 U912 ( .A1(n821), .A2(n820), .ZN(n823) );
  NAND2_X1 U913 ( .A1(n822), .A2(n892), .ZN(n947) );
  NAND2_X1 U914 ( .A1(n823), .A2(n947), .ZN(n824) );
  XOR2_X1 U915 ( .A(KEYINPUT103), .B(n824), .Z(n825) );
  NAND2_X1 U916 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U917 ( .A(KEYINPUT104), .B(n827), .ZN(n828) );
  NAND2_X1 U918 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U919 ( .A(n830), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n831), .ZN(G217) );
  AND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n832) );
  NAND2_X1 U922 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n833) );
  XNOR2_X1 U924 ( .A(KEYINPUT106), .B(n833), .ZN(n835) );
  NAND2_X1 U925 ( .A1(n835), .A2(n834), .ZN(G188) );
  XNOR2_X1 U926 ( .A(G69), .B(KEYINPUT107), .ZN(G235) );
  INV_X1 U928 ( .A(G132), .ZN(G219) );
  INV_X1 U929 ( .A(G96), .ZN(G221) );
  INV_X1 U930 ( .A(G82), .ZN(G220) );
  NOR2_X1 U931 ( .A1(n837), .A2(n836), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U933 ( .A(G1348), .B(G2454), .ZN(n838) );
  XNOR2_X1 U934 ( .A(n838), .B(G2430), .ZN(n839) );
  XNOR2_X1 U935 ( .A(n839), .B(G1341), .ZN(n845) );
  XOR2_X1 U936 ( .A(G2443), .B(G2427), .Z(n841) );
  XNOR2_X1 U937 ( .A(G2438), .B(G2446), .ZN(n840) );
  XNOR2_X1 U938 ( .A(n841), .B(n840), .ZN(n843) );
  XOR2_X1 U939 ( .A(G2451), .B(G2435), .Z(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(n844) );
  XNOR2_X1 U941 ( .A(n845), .B(n844), .ZN(n846) );
  NAND2_X1 U942 ( .A1(n846), .A2(G14), .ZN(n847) );
  XNOR2_X1 U943 ( .A(KEYINPUT105), .B(n847), .ZN(G401) );
  XNOR2_X1 U944 ( .A(G1991), .B(G2474), .ZN(n857) );
  XOR2_X1 U945 ( .A(G1986), .B(G1961), .Z(n849) );
  XNOR2_X1 U946 ( .A(G1996), .B(G1956), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U948 ( .A(G1976), .B(G1981), .Z(n851) );
  XNOR2_X1 U949 ( .A(G1966), .B(G1971), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U951 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U952 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U954 ( .A(n857), .B(n856), .ZN(G229) );
  XOR2_X1 U955 ( .A(G2678), .B(KEYINPUT42), .Z(n859) );
  XNOR2_X1 U956 ( .A(KEYINPUT109), .B(KEYINPUT43), .ZN(n858) );
  XNOR2_X1 U957 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U958 ( .A(KEYINPUT108), .B(G2090), .Z(n861) );
  XNOR2_X1 U959 ( .A(G2067), .B(G2072), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U961 ( .A(n863), .B(n862), .Z(n865) );
  XNOR2_X1 U962 ( .A(G2096), .B(G2100), .ZN(n864) );
  XNOR2_X1 U963 ( .A(n865), .B(n864), .ZN(n867) );
  XOR2_X1 U964 ( .A(G2078), .B(G2084), .Z(n866) );
  XNOR2_X1 U965 ( .A(n867), .B(n866), .ZN(G227) );
  NAND2_X1 U966 ( .A1(G100), .A2(n893), .ZN(n869) );
  NAND2_X1 U967 ( .A1(G112), .A2(n899), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U969 ( .A(n870), .B(KEYINPUT111), .ZN(n872) );
  NAND2_X1 U970 ( .A1(G136), .A2(n895), .ZN(n871) );
  NAND2_X1 U971 ( .A1(n872), .A2(n871), .ZN(n875) );
  NAND2_X1 U972 ( .A1(n902), .A2(G124), .ZN(n873) );
  XOR2_X1 U973 ( .A(KEYINPUT44), .B(n873), .Z(n874) );
  NOR2_X1 U974 ( .A1(n875), .A2(n874), .ZN(G162) );
  XNOR2_X1 U975 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n884) );
  NAND2_X1 U976 ( .A1(G103), .A2(n893), .ZN(n877) );
  NAND2_X1 U977 ( .A1(G139), .A2(n895), .ZN(n876) );
  NAND2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n882) );
  NAND2_X1 U979 ( .A1(G115), .A2(n899), .ZN(n879) );
  NAND2_X1 U980 ( .A1(G127), .A2(n902), .ZN(n878) );
  NAND2_X1 U981 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U982 ( .A(KEYINPUT47), .B(n880), .Z(n881) );
  NOR2_X1 U983 ( .A1(n882), .A2(n881), .ZN(n949) );
  XNOR2_X1 U984 ( .A(n961), .B(n949), .ZN(n883) );
  XNOR2_X1 U985 ( .A(n884), .B(n883), .ZN(n890) );
  XNOR2_X1 U986 ( .A(G162), .B(n885), .ZN(n888) );
  XOR2_X1 U987 ( .A(G160), .B(n886), .Z(n887) );
  XNOR2_X1 U988 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U989 ( .A(n890), .B(n889), .Z(n891) );
  XNOR2_X1 U990 ( .A(n892), .B(n891), .ZN(n908) );
  NAND2_X1 U991 ( .A1(n893), .A2(G106), .ZN(n894) );
  XOR2_X1 U992 ( .A(KEYINPUT113), .B(n894), .Z(n897) );
  NAND2_X1 U993 ( .A1(n895), .A2(G142), .ZN(n896) );
  NAND2_X1 U994 ( .A1(n897), .A2(n896), .ZN(n898) );
  XNOR2_X1 U995 ( .A(n898), .B(KEYINPUT45), .ZN(n901) );
  NAND2_X1 U996 ( .A1(G118), .A2(n899), .ZN(n900) );
  NAND2_X1 U997 ( .A1(n901), .A2(n900), .ZN(n905) );
  NAND2_X1 U998 ( .A1(n902), .A2(G130), .ZN(n903) );
  XOR2_X1 U999 ( .A(KEYINPUT112), .B(n903), .Z(n904) );
  NOR2_X1 U1000 ( .A1(n905), .A2(n904), .ZN(n906) );
  XOR2_X1 U1001 ( .A(G164), .B(n906), .Z(n907) );
  XNOR2_X1 U1002 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n909), .ZN(G395) );
  XNOR2_X1 U1004 ( .A(KEYINPUT114), .B(n984), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(n910), .B(G286), .ZN(n911) );
  XNOR2_X1 U1006 ( .A(n912), .B(n911), .ZN(n914) );
  XNOR2_X1 U1007 ( .A(n995), .B(G171), .ZN(n913) );
  XNOR2_X1 U1008 ( .A(n914), .B(n913), .ZN(n915) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n915), .ZN(G397) );
  OR2_X1 U1010 ( .A1(n921), .A2(G401), .ZN(n918) );
  NOR2_X1 U1011 ( .A1(G229), .A2(G227), .ZN(n916) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n916), .ZN(n917) );
  NOR2_X1 U1013 ( .A1(n918), .A2(n917), .ZN(n920) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n919) );
  NAND2_X1 U1015 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(n921), .ZN(G319) );
  XNOR2_X1 U1018 ( .A(G5), .B(n922), .ZN(n935) );
  XNOR2_X1 U1019 ( .A(G1348), .B(KEYINPUT59), .ZN(n923) );
  XNOR2_X1 U1020 ( .A(n923), .B(G4), .ZN(n927) );
  XNOR2_X1 U1021 ( .A(G1341), .B(G19), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(G20), .B(G1956), .ZN(n924) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n930) );
  XNOR2_X1 U1025 ( .A(KEYINPUT126), .B(G1981), .ZN(n928) );
  XNOR2_X1 U1026 ( .A(G6), .B(n928), .ZN(n929) );
  NOR2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1028 ( .A(KEYINPUT60), .B(n931), .Z(n933) );
  XNOR2_X1 U1029 ( .A(G1966), .B(G21), .ZN(n932) );
  NOR2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n942) );
  XNOR2_X1 U1032 ( .A(G1971), .B(G22), .ZN(n937) );
  XNOR2_X1 U1033 ( .A(G24), .B(G1986), .ZN(n936) );
  NOR2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n939) );
  XOR2_X1 U1035 ( .A(G1976), .B(G23), .Z(n938) );
  NAND2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1037 ( .A(KEYINPUT58), .B(n940), .ZN(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1039 ( .A(KEYINPUT61), .B(n943), .Z(n944) );
  NOR2_X1 U1040 ( .A1(G16), .A2(n944), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(KEYINPUT127), .B(n945), .ZN(n946) );
  NAND2_X1 U1042 ( .A1(n946), .A2(G11), .ZN(n976) );
  NAND2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n969) );
  XOR2_X1 U1044 ( .A(G2072), .B(n949), .Z(n951) );
  XOR2_X1 U1045 ( .A(G164), .B(G2078), .Z(n950) );
  NOR2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1047 ( .A(KEYINPUT50), .B(n952), .Z(n958) );
  XOR2_X1 U1048 ( .A(G2090), .B(G162), .Z(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1050 ( .A(KEYINPUT51), .B(n955), .Z(n956) );
  XOR2_X1 U1051 ( .A(KEYINPUT116), .B(n956), .Z(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n967) );
  XOR2_X1 U1053 ( .A(G2084), .B(G160), .Z(n959) );
  NOR2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n962) );
  NAND2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n964) );
  NOR2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1057 ( .A(KEYINPUT115), .B(n965), .Z(n966) );
  NAND2_X1 U1058 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1059 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1060 ( .A(n970), .B(KEYINPUT52), .ZN(n972) );
  INV_X1 U1061 ( .A(KEYINPUT55), .ZN(n971) );
  NAND2_X1 U1062 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1063 ( .A1(G29), .A2(n973), .ZN(n974) );
  XNOR2_X1 U1064 ( .A(KEYINPUT117), .B(n974), .ZN(n975) );
  NOR2_X1 U1065 ( .A1(n976), .A2(n975), .ZN(n1005) );
  XNOR2_X1 U1066 ( .A(G16), .B(KEYINPUT56), .ZN(n977) );
  XNOR2_X1 U1067 ( .A(n977), .B(KEYINPUT122), .ZN(n1003) );
  XNOR2_X1 U1068 ( .A(G1966), .B(G168), .ZN(n979) );
  NAND2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1070 ( .A(n980), .B(KEYINPUT57), .ZN(n989) );
  XNOR2_X1 U1071 ( .A(G171), .B(G1961), .ZN(n983) );
  XNOR2_X1 U1072 ( .A(G1956), .B(KEYINPUT123), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(n981), .B(G299), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n987) );
  XOR2_X1 U1075 ( .A(G1341), .B(n984), .Z(n985) );
  XNOR2_X1 U1076 ( .A(KEYINPUT125), .B(n985), .ZN(n986) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1079 ( .A1(n991), .A2(n990), .ZN(n1001) );
  XOR2_X1 U1080 ( .A(n992), .B(KEYINPUT124), .Z(n994) );
  XNOR2_X1 U1081 ( .A(G166), .B(G1971), .ZN(n993) );
  NAND2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n999) );
  XNOR2_X1 U1083 ( .A(n995), .B(G1348), .ZN(n997) );
  NAND2_X1 U1084 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1085 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1086 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1087 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1088 ( .A1(n1005), .A2(n1004), .ZN(n1029) );
  XOR2_X1 U1089 ( .A(G2067), .B(G26), .Z(n1008) );
  XNOR2_X1 U1090 ( .A(n1006), .B(G27), .ZN(n1007) );
  NAND2_X1 U1091 ( .A1(n1008), .A2(n1007), .ZN(n1014) );
  XNOR2_X1 U1092 ( .A(G1996), .B(G32), .ZN(n1009) );
  XNOR2_X1 U1093 ( .A(n1009), .B(KEYINPUT119), .ZN(n1012) );
  XOR2_X1 U1094 ( .A(G2072), .B(KEYINPUT118), .Z(n1010) );
  XNOR2_X1 U1095 ( .A(G33), .B(n1010), .ZN(n1011) );
  NAND2_X1 U1096 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1097 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1098 ( .A(KEYINPUT120), .B(n1015), .ZN(n1016) );
  NAND2_X1 U1099 ( .A1(n1016), .A2(G28), .ZN(n1018) );
  XNOR2_X1 U1100 ( .A(G25), .B(G1991), .ZN(n1017) );
  NOR2_X1 U1101 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1102 ( .A(KEYINPUT53), .B(n1019), .Z(n1023) );
  XNOR2_X1 U1103 ( .A(KEYINPUT54), .B(G34), .ZN(n1020) );
  XNOR2_X1 U1104 ( .A(n1020), .B(KEYINPUT121), .ZN(n1021) );
  XNOR2_X1 U1105 ( .A(G2084), .B(n1021), .ZN(n1022) );
  NAND2_X1 U1106 ( .A1(n1023), .A2(n1022), .ZN(n1025) );
  XNOR2_X1 U1107 ( .A(G35), .B(G2090), .ZN(n1024) );
  NOR2_X1 U1108 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1109 ( .A(KEYINPUT55), .B(n1026), .Z(n1027) );
  NOR2_X1 U1110 ( .A1(G29), .A2(n1027), .ZN(n1028) );
  NOR2_X1 U1111 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1112 ( .A(n1030), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

