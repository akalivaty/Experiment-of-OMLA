

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U549 ( .A(n520), .B(KEYINPUT65), .ZN(n871) );
  XNOR2_X1 U550 ( .A(n687), .B(n686), .ZN(n692) );
  NOR2_X1 U551 ( .A1(n677), .A2(n998), .ZN(n683) );
  OR2_X1 U552 ( .A1(n683), .A2(n990), .ZN(n684) );
  INV_X1 U553 ( .A(KEYINPUT91), .ZN(n686) );
  INV_X1 U554 ( .A(n672), .ZN(n700) );
  INV_X1 U555 ( .A(KEYINPUT29), .ZN(n698) );
  XNOR2_X1 U556 ( .A(n699), .B(n698), .ZN(n704) );
  NAND2_X1 U557 ( .A1(n670), .A2(n756), .ZN(n672) );
  NOR2_X1 U558 ( .A1(G2104), .A2(G2105), .ZN(n513) );
  INV_X1 U559 ( .A(KEYINPUT83), .ZN(n548) );
  NOR2_X1 U560 ( .A1(G651), .A2(n641), .ZN(n636) );
  XNOR2_X1 U561 ( .A(n549), .B(n548), .ZN(n551) );
  INV_X1 U562 ( .A(KEYINPUT64), .ZN(n524) );
  XNOR2_X1 U563 ( .A(n525), .B(n524), .ZN(G160) );
  XOR2_X2 U564 ( .A(KEYINPUT17), .B(n513), .Z(n880) );
  NAND2_X1 U565 ( .A1(G137), .A2(n880), .ZN(n515) );
  INV_X1 U566 ( .A(G2105), .ZN(n516) );
  NOR2_X1 U567 ( .A1(G2104), .A2(n516), .ZN(n873) );
  NAND2_X1 U568 ( .A1(G125), .A2(n873), .ZN(n514) );
  NAND2_X1 U569 ( .A1(n515), .A2(n514), .ZN(n519) );
  AND2_X1 U570 ( .A1(n516), .A2(G2104), .ZN(n877) );
  NAND2_X1 U571 ( .A1(G101), .A2(n877), .ZN(n517) );
  XNOR2_X1 U572 ( .A(KEYINPUT23), .B(n517), .ZN(n518) );
  NOR2_X1 U573 ( .A1(n519), .A2(n518), .ZN(n523) );
  NAND2_X1 U574 ( .A1(G2105), .A2(G2104), .ZN(n520) );
  NAND2_X1 U575 ( .A1(n871), .A2(G113), .ZN(n521) );
  XNOR2_X1 U576 ( .A(n521), .B(KEYINPUT66), .ZN(n522) );
  NAND2_X1 U577 ( .A1(n523), .A2(n522), .ZN(n525) );
  AND2_X1 U578 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U579 ( .A1(G99), .A2(n877), .ZN(n534) );
  NAND2_X1 U580 ( .A1(G123), .A2(n873), .ZN(n526) );
  XNOR2_X1 U581 ( .A(n526), .B(KEYINPUT18), .ZN(n529) );
  NAND2_X1 U582 ( .A1(G135), .A2(n880), .ZN(n527) );
  XNOR2_X1 U583 ( .A(n527), .B(KEYINPUT76), .ZN(n528) );
  NAND2_X1 U584 ( .A1(n529), .A2(n528), .ZN(n532) );
  NAND2_X1 U585 ( .A1(G111), .A2(n871), .ZN(n530) );
  XNOR2_X1 U586 ( .A(KEYINPUT77), .B(n530), .ZN(n531) );
  NOR2_X1 U587 ( .A1(n532), .A2(n531), .ZN(n533) );
  NAND2_X1 U588 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U589 ( .A(n535), .B(KEYINPUT78), .ZN(n940) );
  XNOR2_X1 U590 ( .A(n940), .B(G2096), .ZN(n536) );
  OR2_X1 U591 ( .A1(G2100), .A2(n536), .ZN(G156) );
  INV_X1 U592 ( .A(G57), .ZN(G237) );
  INV_X1 U593 ( .A(G132), .ZN(G219) );
  INV_X1 U594 ( .A(G651), .ZN(n541) );
  NOR2_X1 U595 ( .A1(G543), .A2(n541), .ZN(n537) );
  XOR2_X1 U596 ( .A(KEYINPUT1), .B(n537), .Z(n640) );
  NAND2_X1 U597 ( .A1(G64), .A2(n640), .ZN(n539) );
  XOR2_X1 U598 ( .A(KEYINPUT0), .B(G543), .Z(n641) );
  NAND2_X1 U599 ( .A1(G52), .A2(n636), .ZN(n538) );
  NAND2_X1 U600 ( .A1(n539), .A2(n538), .ZN(n547) );
  NOR2_X1 U601 ( .A1(G651), .A2(G543), .ZN(n627) );
  NAND2_X1 U602 ( .A1(n627), .A2(G90), .ZN(n540) );
  XNOR2_X1 U603 ( .A(n540), .B(KEYINPUT68), .ZN(n543) );
  NOR2_X1 U604 ( .A1(n641), .A2(n541), .ZN(n630) );
  NAND2_X1 U605 ( .A1(G77), .A2(n630), .ZN(n542) );
  NAND2_X1 U606 ( .A1(n543), .A2(n542), .ZN(n545) );
  XOR2_X1 U607 ( .A(KEYINPUT9), .B(KEYINPUT69), .Z(n544) );
  XOR2_X1 U608 ( .A(n545), .B(n544), .Z(n546) );
  NOR2_X1 U609 ( .A1(n547), .A2(n546), .ZN(G171) );
  NAND2_X1 U610 ( .A1(G138), .A2(n880), .ZN(n549) );
  NAND2_X1 U611 ( .A1(n877), .A2(G102), .ZN(n550) );
  NAND2_X1 U612 ( .A1(n551), .A2(n550), .ZN(n555) );
  NAND2_X1 U613 ( .A1(G126), .A2(n873), .ZN(n553) );
  NAND2_X1 U614 ( .A1(G114), .A2(n871), .ZN(n552) );
  NAND2_X1 U615 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U616 ( .A1(n555), .A2(n554), .ZN(G164) );
  NAND2_X1 U617 ( .A1(G63), .A2(n640), .ZN(n557) );
  NAND2_X1 U618 ( .A1(G51), .A2(n636), .ZN(n556) );
  NAND2_X1 U619 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U620 ( .A(KEYINPUT6), .B(n558), .Z(n566) );
  NAND2_X1 U621 ( .A1(n630), .A2(G76), .ZN(n559) );
  XNOR2_X1 U622 ( .A(KEYINPUT73), .B(n559), .ZN(n562) );
  NAND2_X1 U623 ( .A1(n627), .A2(G89), .ZN(n560) );
  XOR2_X1 U624 ( .A(n560), .B(KEYINPUT4), .Z(n561) );
  NOR2_X1 U625 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U626 ( .A(KEYINPUT5), .B(n563), .Z(n564) );
  XNOR2_X1 U627 ( .A(KEYINPUT74), .B(n564), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U629 ( .A(KEYINPUT7), .B(n567), .ZN(G168) );
  XOR2_X1 U630 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U631 ( .A1(G7), .A2(G661), .ZN(n568) );
  XNOR2_X1 U632 ( .A(n568), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U633 ( .A(G223), .ZN(n813) );
  NAND2_X1 U634 ( .A1(n813), .A2(G567), .ZN(n569) );
  XOR2_X1 U635 ( .A(KEYINPUT11), .B(n569), .Z(G234) );
  NAND2_X1 U636 ( .A1(G56), .A2(n640), .ZN(n570) );
  XOR2_X1 U637 ( .A(KEYINPUT14), .B(n570), .Z(n577) );
  NAND2_X1 U638 ( .A1(n627), .A2(G81), .ZN(n571) );
  XOR2_X1 U639 ( .A(KEYINPUT12), .B(n571), .Z(n574) );
  NAND2_X1 U640 ( .A1(n630), .A2(G68), .ZN(n572) );
  XOR2_X1 U641 ( .A(KEYINPUT72), .B(n572), .Z(n573) );
  NOR2_X1 U642 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U643 ( .A(n575), .B(KEYINPUT13), .ZN(n576) );
  NOR2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U645 ( .A1(n636), .A2(G43), .ZN(n578) );
  NAND2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n998) );
  INV_X1 U647 ( .A(G860), .ZN(n606) );
  OR2_X1 U648 ( .A1(n998), .A2(n606), .ZN(G153) );
  INV_X1 U649 ( .A(G171), .ZN(G301) );
  NAND2_X1 U650 ( .A1(G868), .A2(G301), .ZN(n588) );
  NAND2_X1 U651 ( .A1(G66), .A2(n640), .ZN(n581) );
  NAND2_X1 U652 ( .A1(G79), .A2(n630), .ZN(n580) );
  NAND2_X1 U653 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U654 ( .A1(G54), .A2(n636), .ZN(n583) );
  NAND2_X1 U655 ( .A1(G92), .A2(n627), .ZN(n582) );
  NAND2_X1 U656 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U657 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U658 ( .A(KEYINPUT15), .B(n586), .Z(n990) );
  OR2_X1 U659 ( .A1(n990), .A2(G868), .ZN(n587) );
  NAND2_X1 U660 ( .A1(n588), .A2(n587), .ZN(G284) );
  NAND2_X1 U661 ( .A1(G91), .A2(n627), .ZN(n590) );
  NAND2_X1 U662 ( .A1(G78), .A2(n630), .ZN(n589) );
  NAND2_X1 U663 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n640), .A2(G65), .ZN(n591) );
  XOR2_X1 U665 ( .A(KEYINPUT70), .B(n591), .Z(n592) );
  NOR2_X1 U666 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U667 ( .A1(n636), .A2(G53), .ZN(n594) );
  NAND2_X1 U668 ( .A1(n595), .A2(n594), .ZN(G299) );
  INV_X1 U669 ( .A(G868), .ZN(n596) );
  NOR2_X1 U670 ( .A1(G286), .A2(n596), .ZN(n598) );
  NOR2_X1 U671 ( .A1(G868), .A2(G299), .ZN(n597) );
  NOR2_X1 U672 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U673 ( .A1(G559), .A2(n606), .ZN(n599) );
  XOR2_X1 U674 ( .A(KEYINPUT75), .B(n599), .Z(n600) );
  NAND2_X1 U675 ( .A1(n600), .A2(n990), .ZN(n601) );
  XNOR2_X1 U676 ( .A(n601), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U677 ( .A1(G868), .A2(n998), .ZN(n604) );
  NAND2_X1 U678 ( .A1(G868), .A2(n990), .ZN(n602) );
  NOR2_X1 U679 ( .A1(G559), .A2(n602), .ZN(n603) );
  NOR2_X1 U680 ( .A1(n604), .A2(n603), .ZN(G282) );
  NAND2_X1 U681 ( .A1(G559), .A2(n990), .ZN(n605) );
  XOR2_X1 U682 ( .A(n998), .B(n605), .Z(n650) );
  NAND2_X1 U683 ( .A1(n606), .A2(n650), .ZN(n613) );
  NAND2_X1 U684 ( .A1(G67), .A2(n640), .ZN(n608) );
  NAND2_X1 U685 ( .A1(G55), .A2(n636), .ZN(n607) );
  NAND2_X1 U686 ( .A1(n608), .A2(n607), .ZN(n612) );
  NAND2_X1 U687 ( .A1(G93), .A2(n627), .ZN(n610) );
  NAND2_X1 U688 ( .A1(G80), .A2(n630), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n652) );
  XOR2_X1 U691 ( .A(n613), .B(n652), .Z(G145) );
  NAND2_X1 U692 ( .A1(G88), .A2(n627), .ZN(n615) );
  NAND2_X1 U693 ( .A1(G75), .A2(n630), .ZN(n614) );
  NAND2_X1 U694 ( .A1(n615), .A2(n614), .ZN(n619) );
  NAND2_X1 U695 ( .A1(G62), .A2(n640), .ZN(n617) );
  NAND2_X1 U696 ( .A1(G50), .A2(n636), .ZN(n616) );
  NAND2_X1 U697 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U698 ( .A1(n619), .A2(n618), .ZN(G166) );
  NAND2_X1 U699 ( .A1(G61), .A2(n640), .ZN(n621) );
  NAND2_X1 U700 ( .A1(G86), .A2(n627), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U702 ( .A1(n630), .A2(G73), .ZN(n622) );
  XOR2_X1 U703 ( .A(KEYINPUT2), .B(n622), .Z(n623) );
  NOR2_X1 U704 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n636), .A2(G48), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n626), .A2(n625), .ZN(G305) );
  NAND2_X1 U707 ( .A1(G60), .A2(n640), .ZN(n629) );
  NAND2_X1 U708 ( .A1(G85), .A2(n627), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U710 ( .A1(G72), .A2(n630), .ZN(n631) );
  XNOR2_X1 U711 ( .A(KEYINPUT67), .B(n631), .ZN(n632) );
  NOR2_X1 U712 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U713 ( .A1(n636), .A2(G47), .ZN(n634) );
  NAND2_X1 U714 ( .A1(n635), .A2(n634), .ZN(G290) );
  NAND2_X1 U715 ( .A1(G49), .A2(n636), .ZN(n638) );
  NAND2_X1 U716 ( .A1(G74), .A2(G651), .ZN(n637) );
  NAND2_X1 U717 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U718 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U719 ( .A1(n641), .A2(G87), .ZN(n642) );
  NAND2_X1 U720 ( .A1(n643), .A2(n642), .ZN(G288) );
  XNOR2_X1 U721 ( .A(G166), .B(KEYINPUT19), .ZN(n644) );
  XNOR2_X1 U722 ( .A(n644), .B(KEYINPUT79), .ZN(n647) );
  INV_X1 U723 ( .A(G299), .ZN(n693) );
  XNOR2_X1 U724 ( .A(n693), .B(G305), .ZN(n645) );
  XNOR2_X1 U725 ( .A(n645), .B(G290), .ZN(n646) );
  XNOR2_X1 U726 ( .A(n647), .B(n646), .ZN(n649) );
  XNOR2_X1 U727 ( .A(G288), .B(n652), .ZN(n648) );
  XNOR2_X1 U728 ( .A(n649), .B(n648), .ZN(n886) );
  XNOR2_X1 U729 ( .A(n650), .B(n886), .ZN(n651) );
  NAND2_X1 U730 ( .A1(n651), .A2(G868), .ZN(n654) );
  OR2_X1 U731 ( .A1(G868), .A2(n652), .ZN(n653) );
  NAND2_X1 U732 ( .A1(n654), .A2(n653), .ZN(G295) );
  XOR2_X1 U733 ( .A(KEYINPUT20), .B(KEYINPUT80), .Z(n656) );
  NAND2_X1 U734 ( .A1(G2084), .A2(G2078), .ZN(n655) );
  XNOR2_X1 U735 ( .A(n656), .B(n655), .ZN(n657) );
  NAND2_X1 U736 ( .A1(n657), .A2(G2090), .ZN(n658) );
  XOR2_X1 U737 ( .A(KEYINPUT21), .B(n658), .Z(n659) );
  XNOR2_X1 U738 ( .A(KEYINPUT81), .B(n659), .ZN(n660) );
  NAND2_X1 U739 ( .A1(n660), .A2(G2072), .ZN(n661) );
  XNOR2_X1 U740 ( .A(KEYINPUT82), .B(n661), .ZN(G158) );
  XNOR2_X1 U741 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U742 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  NOR2_X1 U743 ( .A1(G219), .A2(G220), .ZN(n662) );
  XOR2_X1 U744 ( .A(KEYINPUT22), .B(n662), .Z(n663) );
  NOR2_X1 U745 ( .A1(G218), .A2(n663), .ZN(n664) );
  NAND2_X1 U746 ( .A1(G96), .A2(n664), .ZN(n819) );
  NAND2_X1 U747 ( .A1(n819), .A2(G2106), .ZN(n668) );
  NAND2_X1 U748 ( .A1(G120), .A2(G108), .ZN(n665) );
  NOR2_X1 U749 ( .A1(G237), .A2(n665), .ZN(n666) );
  NAND2_X1 U750 ( .A1(G69), .A2(n666), .ZN(n820) );
  NAND2_X1 U751 ( .A1(n820), .A2(G567), .ZN(n667) );
  NAND2_X1 U752 ( .A1(n668), .A2(n667), .ZN(n821) );
  NAND2_X1 U753 ( .A1(G661), .A2(G483), .ZN(n669) );
  NOR2_X1 U754 ( .A1(n821), .A2(n669), .ZN(n816) );
  NAND2_X1 U755 ( .A1(n816), .A2(G36), .ZN(G176) );
  INV_X1 U756 ( .A(G166), .ZN(G303) );
  INV_X1 U757 ( .A(KEYINPUT89), .ZN(n676) );
  NAND2_X1 U758 ( .A1(G40), .A2(G160), .ZN(n755) );
  INV_X1 U759 ( .A(n755), .ZN(n670) );
  NOR2_X1 U760 ( .A1(G164), .A2(G1384), .ZN(n756) );
  NAND2_X1 U761 ( .A1(n700), .A2(G1996), .ZN(n671) );
  XNOR2_X1 U762 ( .A(n671), .B(KEYINPUT26), .ZN(n674) );
  NAND2_X1 U763 ( .A1(G1341), .A2(n672), .ZN(n673) );
  NAND2_X1 U764 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U765 ( .A(n676), .B(n675), .ZN(n677) );
  NAND2_X1 U766 ( .A1(n683), .A2(n990), .ZN(n682) );
  NAND2_X1 U767 ( .A1(G1348), .A2(n672), .ZN(n679) );
  NAND2_X1 U768 ( .A1(n700), .A2(G2067), .ZN(n678) );
  NAND2_X1 U769 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U770 ( .A(KEYINPUT90), .B(n680), .ZN(n681) );
  NAND2_X1 U771 ( .A1(n682), .A2(n681), .ZN(n685) );
  NAND2_X1 U772 ( .A1(n685), .A2(n684), .ZN(n687) );
  NAND2_X1 U773 ( .A1(n700), .A2(G2072), .ZN(n688) );
  XNOR2_X1 U774 ( .A(n688), .B(KEYINPUT27), .ZN(n690) );
  AND2_X1 U775 ( .A1(G1956), .A2(n672), .ZN(n689) );
  NOR2_X1 U776 ( .A1(n690), .A2(n689), .ZN(n694) );
  NAND2_X1 U777 ( .A1(n694), .A2(n693), .ZN(n691) );
  NAND2_X1 U778 ( .A1(n692), .A2(n691), .ZN(n697) );
  NOR2_X1 U779 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U780 ( .A(n695), .B(KEYINPUT28), .Z(n696) );
  NAND2_X1 U781 ( .A1(n697), .A2(n696), .ZN(n699) );
  XOR2_X1 U782 ( .A(KEYINPUT88), .B(G1961), .Z(n968) );
  NAND2_X1 U783 ( .A1(n968), .A2(n672), .ZN(n702) );
  XNOR2_X1 U784 ( .A(KEYINPUT25), .B(G2078), .ZN(n913) );
  NAND2_X1 U785 ( .A1(n700), .A2(n913), .ZN(n701) );
  NAND2_X1 U786 ( .A1(n702), .A2(n701), .ZN(n709) );
  NAND2_X1 U787 ( .A1(n709), .A2(G171), .ZN(n703) );
  NAND2_X1 U788 ( .A1(n704), .A2(n703), .ZN(n729) );
  NAND2_X1 U789 ( .A1(G8), .A2(n672), .ZN(n786) );
  NOR2_X1 U790 ( .A1(G1966), .A2(n786), .ZN(n715) );
  NOR2_X1 U791 ( .A1(n672), .A2(G2084), .ZN(n717) );
  XNOR2_X1 U792 ( .A(n717), .B(KEYINPUT87), .ZN(n705) );
  NAND2_X1 U793 ( .A1(G8), .A2(n705), .ZN(n706) );
  NOR2_X1 U794 ( .A1(n715), .A2(n706), .ZN(n707) );
  XOR2_X1 U795 ( .A(KEYINPUT30), .B(n707), .Z(n708) );
  NOR2_X1 U796 ( .A1(G168), .A2(n708), .ZN(n711) );
  NOR2_X1 U797 ( .A1(G171), .A2(n709), .ZN(n710) );
  NOR2_X1 U798 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U799 ( .A(KEYINPUT31), .B(n712), .Z(n727) );
  NAND2_X1 U800 ( .A1(n729), .A2(n727), .ZN(n714) );
  INV_X1 U801 ( .A(KEYINPUT92), .ZN(n713) );
  XNOR2_X1 U802 ( .A(n714), .B(n713), .ZN(n716) );
  NOR2_X1 U803 ( .A1(n716), .A2(n715), .ZN(n720) );
  XOR2_X1 U804 ( .A(KEYINPUT87), .B(n717), .Z(n718) );
  NAND2_X1 U805 ( .A1(G8), .A2(n718), .ZN(n719) );
  NAND2_X1 U806 ( .A1(n720), .A2(n719), .ZN(n737) );
  INV_X1 U807 ( .A(G8), .ZN(n726) );
  NOR2_X1 U808 ( .A1(G1971), .A2(n786), .ZN(n722) );
  NOR2_X1 U809 ( .A1(G2090), .A2(n672), .ZN(n721) );
  NOR2_X1 U810 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U811 ( .A(KEYINPUT93), .B(n723), .Z(n724) );
  NAND2_X1 U812 ( .A1(n724), .A2(G303), .ZN(n725) );
  OR2_X1 U813 ( .A1(n726), .A2(n725), .ZN(n730) );
  AND2_X1 U814 ( .A1(n727), .A2(n730), .ZN(n728) );
  NAND2_X1 U815 ( .A1(n729), .A2(n728), .ZN(n734) );
  INV_X1 U816 ( .A(n730), .ZN(n732) );
  AND2_X1 U817 ( .A1(G286), .A2(G8), .ZN(n731) );
  OR2_X1 U818 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U819 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U820 ( .A(n735), .B(KEYINPUT32), .ZN(n736) );
  NAND2_X1 U821 ( .A1(n737), .A2(n736), .ZN(n780) );
  NOR2_X1 U822 ( .A1(G2090), .A2(G303), .ZN(n738) );
  NAND2_X1 U823 ( .A1(G8), .A2(n738), .ZN(n739) );
  NAND2_X1 U824 ( .A1(n780), .A2(n739), .ZN(n740) );
  AND2_X1 U825 ( .A1(n740), .A2(n786), .ZN(n745) );
  NOR2_X1 U826 ( .A1(G1981), .A2(G305), .ZN(n741) );
  XOR2_X1 U827 ( .A(n741), .B(KEYINPUT24), .Z(n742) );
  XNOR2_X1 U828 ( .A(KEYINPUT86), .B(n742), .ZN(n743) );
  NOR2_X1 U829 ( .A1(n786), .A2(n743), .ZN(n744) );
  NOR2_X1 U830 ( .A1(n745), .A2(n744), .ZN(n776) );
  NAND2_X1 U831 ( .A1(G140), .A2(n880), .ZN(n747) );
  NAND2_X1 U832 ( .A1(G104), .A2(n877), .ZN(n746) );
  NAND2_X1 U833 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U834 ( .A(KEYINPUT34), .B(n748), .ZN(n753) );
  NAND2_X1 U835 ( .A1(G128), .A2(n873), .ZN(n750) );
  NAND2_X1 U836 ( .A1(G116), .A2(n871), .ZN(n749) );
  NAND2_X1 U837 ( .A1(n750), .A2(n749), .ZN(n751) );
  XOR2_X1 U838 ( .A(KEYINPUT35), .B(n751), .Z(n752) );
  NOR2_X1 U839 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U840 ( .A(KEYINPUT36), .B(n754), .ZN(n866) );
  XNOR2_X1 U841 ( .A(G2067), .B(KEYINPUT37), .ZN(n805) );
  NOR2_X1 U842 ( .A1(n866), .A2(n805), .ZN(n937) );
  NOR2_X1 U843 ( .A1(n756), .A2(n755), .ZN(n808) );
  NAND2_X1 U844 ( .A1(n937), .A2(n808), .ZN(n757) );
  XNOR2_X1 U845 ( .A(n757), .B(KEYINPUT84), .ZN(n803) );
  NAND2_X1 U846 ( .A1(G131), .A2(n880), .ZN(n759) );
  NAND2_X1 U847 ( .A1(G95), .A2(n877), .ZN(n758) );
  NAND2_X1 U848 ( .A1(n759), .A2(n758), .ZN(n762) );
  NAND2_X1 U849 ( .A1(G119), .A2(n873), .ZN(n760) );
  XNOR2_X1 U850 ( .A(KEYINPUT85), .B(n760), .ZN(n761) );
  NOR2_X1 U851 ( .A1(n762), .A2(n761), .ZN(n764) );
  NAND2_X1 U852 ( .A1(n871), .A2(G107), .ZN(n763) );
  NAND2_X1 U853 ( .A1(n764), .A2(n763), .ZN(n861) );
  AND2_X1 U854 ( .A1(n861), .A2(G1991), .ZN(n773) );
  NAND2_X1 U855 ( .A1(G141), .A2(n880), .ZN(n766) );
  NAND2_X1 U856 ( .A1(G117), .A2(n871), .ZN(n765) );
  NAND2_X1 U857 ( .A1(n766), .A2(n765), .ZN(n769) );
  NAND2_X1 U858 ( .A1(n877), .A2(G105), .ZN(n767) );
  XOR2_X1 U859 ( .A(KEYINPUT38), .B(n767), .Z(n768) );
  NOR2_X1 U860 ( .A1(n769), .A2(n768), .ZN(n771) );
  NAND2_X1 U861 ( .A1(n873), .A2(G129), .ZN(n770) );
  NAND2_X1 U862 ( .A1(n771), .A2(n770), .ZN(n859) );
  AND2_X1 U863 ( .A1(n859), .A2(G1996), .ZN(n772) );
  NOR2_X1 U864 ( .A1(n773), .A2(n772), .ZN(n939) );
  INV_X1 U865 ( .A(n808), .ZN(n774) );
  NOR2_X1 U866 ( .A1(n939), .A2(n774), .ZN(n800) );
  INV_X1 U867 ( .A(n800), .ZN(n775) );
  NAND2_X1 U868 ( .A1(n803), .A2(n775), .ZN(n790) );
  OR2_X1 U869 ( .A1(n776), .A2(n790), .ZN(n795) );
  NOR2_X1 U870 ( .A1(G1976), .A2(G288), .ZN(n785) );
  NOR2_X1 U871 ( .A1(G1971), .A2(G303), .ZN(n777) );
  NOR2_X1 U872 ( .A1(n785), .A2(n777), .ZN(n995) );
  INV_X1 U873 ( .A(KEYINPUT33), .ZN(n778) );
  AND2_X1 U874 ( .A1(n995), .A2(n778), .ZN(n779) );
  NAND2_X1 U875 ( .A1(n780), .A2(n779), .ZN(n784) );
  INV_X1 U876 ( .A(n786), .ZN(n781) );
  NAND2_X1 U877 ( .A1(G1976), .A2(G288), .ZN(n994) );
  AND2_X1 U878 ( .A1(n781), .A2(n994), .ZN(n782) );
  OR2_X1 U879 ( .A1(KEYINPUT33), .A2(n782), .ZN(n783) );
  NAND2_X1 U880 ( .A1(n784), .A2(n783), .ZN(n789) );
  NAND2_X1 U881 ( .A1(n785), .A2(KEYINPUT33), .ZN(n787) );
  NOR2_X1 U882 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U883 ( .A1(n789), .A2(n788), .ZN(n793) );
  XOR2_X1 U884 ( .A(G1981), .B(G305), .Z(n999) );
  INV_X1 U885 ( .A(n790), .ZN(n791) );
  AND2_X1 U886 ( .A1(n999), .A2(n791), .ZN(n792) );
  NAND2_X1 U887 ( .A1(n793), .A2(n792), .ZN(n794) );
  NAND2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n797) );
  XNOR2_X1 U889 ( .A(G1986), .B(G290), .ZN(n1008) );
  NAND2_X1 U890 ( .A1(n1008), .A2(n808), .ZN(n796) );
  NAND2_X1 U891 ( .A1(n797), .A2(n796), .ZN(n811) );
  NOR2_X1 U892 ( .A1(G1996), .A2(n859), .ZN(n934) );
  NOR2_X1 U893 ( .A1(G1986), .A2(G290), .ZN(n798) );
  NOR2_X1 U894 ( .A1(G1991), .A2(n861), .ZN(n943) );
  NOR2_X1 U895 ( .A1(n798), .A2(n943), .ZN(n799) );
  NOR2_X1 U896 ( .A1(n800), .A2(n799), .ZN(n801) );
  NOR2_X1 U897 ( .A1(n934), .A2(n801), .ZN(n802) );
  XNOR2_X1 U898 ( .A(n802), .B(KEYINPUT39), .ZN(n804) );
  NAND2_X1 U899 ( .A1(n804), .A2(n803), .ZN(n806) );
  NAND2_X1 U900 ( .A1(n866), .A2(n805), .ZN(n938) );
  NAND2_X1 U901 ( .A1(n806), .A2(n938), .ZN(n807) );
  NAND2_X1 U902 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U903 ( .A(KEYINPUT94), .B(n809), .ZN(n810) );
  NAND2_X1 U904 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U905 ( .A(n812), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U906 ( .A1(G2106), .A2(n813), .ZN(G217) );
  AND2_X1 U907 ( .A1(G15), .A2(G2), .ZN(n814) );
  NAND2_X1 U908 ( .A1(G661), .A2(n814), .ZN(G259) );
  NAND2_X1 U909 ( .A1(G3), .A2(G1), .ZN(n815) );
  XNOR2_X1 U910 ( .A(KEYINPUT98), .B(n815), .ZN(n817) );
  NAND2_X1 U911 ( .A1(n817), .A2(n816), .ZN(n818) );
  XOR2_X1 U912 ( .A(KEYINPUT99), .B(n818), .Z(G188) );
  NOR2_X1 U913 ( .A1(n820), .A2(n819), .ZN(G325) );
  XOR2_X1 U914 ( .A(KEYINPUT100), .B(G325), .Z(G261) );
  XOR2_X1 U915 ( .A(G108), .B(KEYINPUT110), .Z(G238) );
  INV_X1 U917 ( .A(G120), .ZN(G236) );
  INV_X1 U918 ( .A(G96), .ZN(G221) );
  INV_X1 U919 ( .A(n821), .ZN(G319) );
  XOR2_X1 U920 ( .A(KEYINPUT101), .B(G2090), .Z(n823) );
  XNOR2_X1 U921 ( .A(G2067), .B(G2084), .ZN(n822) );
  XNOR2_X1 U922 ( .A(n823), .B(n822), .ZN(n824) );
  XOR2_X1 U923 ( .A(n824), .B(G2100), .Z(n826) );
  XNOR2_X1 U924 ( .A(G2078), .B(G2072), .ZN(n825) );
  XNOR2_X1 U925 ( .A(n826), .B(n825), .ZN(n830) );
  XOR2_X1 U926 ( .A(G2096), .B(KEYINPUT43), .Z(n828) );
  XNOR2_X1 U927 ( .A(KEYINPUT42), .B(G2678), .ZN(n827) );
  XNOR2_X1 U928 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U929 ( .A(n830), .B(n829), .Z(G227) );
  XOR2_X1 U930 ( .A(KEYINPUT41), .B(G1991), .Z(n832) );
  XNOR2_X1 U931 ( .A(G1996), .B(G1976), .ZN(n831) );
  XNOR2_X1 U932 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U933 ( .A(n833), .B(KEYINPUT103), .Z(n835) );
  XNOR2_X1 U934 ( .A(G1956), .B(G1981), .ZN(n834) );
  XNOR2_X1 U935 ( .A(n835), .B(n834), .ZN(n839) );
  XOR2_X1 U936 ( .A(G1986), .B(G1971), .Z(n837) );
  XNOR2_X1 U937 ( .A(G1966), .B(G1961), .ZN(n836) );
  XNOR2_X1 U938 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U939 ( .A(n839), .B(n838), .Z(n841) );
  XNOR2_X1 U940 ( .A(KEYINPUT102), .B(G2474), .ZN(n840) );
  XNOR2_X1 U941 ( .A(n841), .B(n840), .ZN(G229) );
  NAND2_X1 U942 ( .A1(G124), .A2(n873), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n842), .B(KEYINPUT44), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n843), .B(KEYINPUT104), .ZN(n845) );
  NAND2_X1 U945 ( .A1(G100), .A2(n877), .ZN(n844) );
  NAND2_X1 U946 ( .A1(n845), .A2(n844), .ZN(n849) );
  NAND2_X1 U947 ( .A1(G136), .A2(n880), .ZN(n847) );
  NAND2_X1 U948 ( .A1(G112), .A2(n871), .ZN(n846) );
  NAND2_X1 U949 ( .A1(n847), .A2(n846), .ZN(n848) );
  NOR2_X1 U950 ( .A1(n849), .A2(n848), .ZN(G162) );
  NAND2_X1 U951 ( .A1(G142), .A2(n880), .ZN(n851) );
  NAND2_X1 U952 ( .A1(G106), .A2(n877), .ZN(n850) );
  NAND2_X1 U953 ( .A1(n851), .A2(n850), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n852), .B(KEYINPUT45), .ZN(n858) );
  NAND2_X1 U955 ( .A1(n873), .A2(G130), .ZN(n853) );
  XOR2_X1 U956 ( .A(KEYINPUT105), .B(n853), .Z(n855) );
  NAND2_X1 U957 ( .A1(n871), .A2(G118), .ZN(n854) );
  NAND2_X1 U958 ( .A1(n855), .A2(n854), .ZN(n856) );
  XOR2_X1 U959 ( .A(KEYINPUT106), .B(n856), .Z(n857) );
  NAND2_X1 U960 ( .A1(n858), .A2(n857), .ZN(n860) );
  XOR2_X1 U961 ( .A(n860), .B(n859), .Z(n865) );
  XOR2_X1 U962 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n863) );
  XOR2_X1 U963 ( .A(G164), .B(n861), .Z(n862) );
  XNOR2_X1 U964 ( .A(n863), .B(n862), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n865), .B(n864), .ZN(n868) );
  XNOR2_X1 U966 ( .A(n866), .B(G162), .ZN(n867) );
  XNOR2_X1 U967 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U968 ( .A(n940), .B(n869), .Z(n870) );
  XNOR2_X1 U969 ( .A(G160), .B(n870), .ZN(n884) );
  NAND2_X1 U970 ( .A1(n871), .A2(G115), .ZN(n872) );
  XNOR2_X1 U971 ( .A(n872), .B(KEYINPUT108), .ZN(n875) );
  NAND2_X1 U972 ( .A1(G127), .A2(n873), .ZN(n874) );
  NAND2_X1 U973 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U974 ( .A(n876), .B(KEYINPUT47), .ZN(n879) );
  NAND2_X1 U975 ( .A1(G103), .A2(n877), .ZN(n878) );
  NAND2_X1 U976 ( .A1(n879), .A2(n878), .ZN(n883) );
  NAND2_X1 U977 ( .A1(G139), .A2(n880), .ZN(n881) );
  XNOR2_X1 U978 ( .A(KEYINPUT107), .B(n881), .ZN(n882) );
  NOR2_X1 U979 ( .A1(n883), .A2(n882), .ZN(n949) );
  XNOR2_X1 U980 ( .A(n884), .B(n949), .ZN(n885) );
  NOR2_X1 U981 ( .A1(G37), .A2(n885), .ZN(G395) );
  XOR2_X1 U982 ( .A(n886), .B(G286), .Z(n888) );
  XNOR2_X1 U983 ( .A(G171), .B(n990), .ZN(n887) );
  XNOR2_X1 U984 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U985 ( .A(n889), .B(n998), .Z(n890) );
  NOR2_X1 U986 ( .A1(G37), .A2(n890), .ZN(G397) );
  XOR2_X1 U987 ( .A(KEYINPUT95), .B(KEYINPUT97), .Z(n892) );
  XNOR2_X1 U988 ( .A(G2446), .B(G2451), .ZN(n891) );
  XNOR2_X1 U989 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U990 ( .A(n893), .B(G2430), .Z(n895) );
  XNOR2_X1 U991 ( .A(G1341), .B(G1348), .ZN(n894) );
  XNOR2_X1 U992 ( .A(n895), .B(n894), .ZN(n899) );
  XOR2_X1 U993 ( .A(G2435), .B(G2438), .Z(n897) );
  XNOR2_X1 U994 ( .A(G2454), .B(KEYINPUT96), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U996 ( .A(n899), .B(n898), .Z(n901) );
  XNOR2_X1 U997 ( .A(G2443), .B(G2427), .ZN(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n902) );
  NAND2_X1 U999 ( .A1(n902), .A2(G14), .ZN(n909) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n909), .ZN(n906) );
  NOR2_X1 U1001 ( .A1(G227), .A2(G229), .ZN(n903) );
  XOR2_X1 U1002 ( .A(KEYINPUT49), .B(n903), .Z(n904) );
  XNOR2_X1 U1003 ( .A(n904), .B(KEYINPUT109), .ZN(n905) );
  NOR2_X1 U1004 ( .A1(n906), .A2(n905), .ZN(n908) );
  NOR2_X1 U1005 ( .A1(G395), .A2(G397), .ZN(n907) );
  NAND2_X1 U1006 ( .A1(n908), .A2(n907), .ZN(G225) );
  INV_X1 U1007 ( .A(G225), .ZN(G308) );
  INV_X1 U1008 ( .A(G69), .ZN(G235) );
  INV_X1 U1009 ( .A(n909), .ZN(G401) );
  XNOR2_X1 U1010 ( .A(KEYINPUT117), .B(G29), .ZN(n931) );
  XNOR2_X1 U1011 ( .A(G25), .B(KEYINPUT114), .ZN(n910) );
  XOR2_X1 U1012 ( .A(n910), .B(G1991), .Z(n911) );
  NAND2_X1 U1013 ( .A1(n911), .A2(G28), .ZN(n912) );
  XNOR2_X1 U1014 ( .A(n912), .B(KEYINPUT115), .ZN(n922) );
  XNOR2_X1 U1015 ( .A(G27), .B(n913), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(G2072), .B(G33), .ZN(n915) );
  XNOR2_X1 U1017 ( .A(G32), .B(G1996), .ZN(n914) );
  NOR2_X1 U1018 ( .A1(n915), .A2(n914), .ZN(n916) );
  NAND2_X1 U1019 ( .A1(n917), .A2(n916), .ZN(n920) );
  XNOR2_X1 U1020 ( .A(KEYINPUT116), .B(G2067), .ZN(n918) );
  XNOR2_X1 U1021 ( .A(G26), .B(n918), .ZN(n919) );
  NOR2_X1 U1022 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1024 ( .A(n923), .B(KEYINPUT53), .ZN(n926) );
  XOR2_X1 U1025 ( .A(G2084), .B(G34), .Z(n924) );
  XNOR2_X1 U1026 ( .A(KEYINPUT54), .B(n924), .ZN(n925) );
  NAND2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n928) );
  XNOR2_X1 U1028 ( .A(G35), .B(G2090), .ZN(n927) );
  NOR2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(KEYINPUT55), .B(n929), .ZN(n930) );
  NAND2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1032 ( .A(KEYINPUT118), .B(n932), .ZN(n962) );
  XOR2_X1 U1033 ( .A(G2090), .B(G162), .Z(n933) );
  NOR2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1035 ( .A(n935), .B(KEYINPUT51), .ZN(n936) );
  NOR2_X1 U1036 ( .A1(n937), .A2(n936), .ZN(n948) );
  NAND2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n946) );
  XNOR2_X1 U1038 ( .A(G2084), .B(G160), .ZN(n941) );
  NAND2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(KEYINPUT111), .B(n944), .ZN(n945) );
  NOR2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n956) );
  XNOR2_X1 U1044 ( .A(G164), .B(G2078), .ZN(n952) );
  XNOR2_X1 U1045 ( .A(G2072), .B(n949), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(n950), .B(KEYINPUT112), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(n953), .B(KEYINPUT113), .ZN(n954) );
  XOR2_X1 U1049 ( .A(KEYINPUT50), .B(n954), .Z(n955) );
  NOR2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(KEYINPUT52), .B(n957), .ZN(n959) );
  INV_X1 U1052 ( .A(KEYINPUT55), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1054 ( .A1(n960), .A2(G29), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n1020) );
  XOR2_X1 U1056 ( .A(G1976), .B(G23), .Z(n964) );
  XOR2_X1 U1057 ( .A(G1971), .B(G22), .Z(n963) );
  NAND2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(G24), .B(G1986), .ZN(n965) );
  NOR2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1061 ( .A(KEYINPUT58), .B(n967), .Z(n987) );
  XNOR2_X1 U1062 ( .A(n968), .B(G5), .ZN(n971) );
  XNOR2_X1 U1063 ( .A(G1966), .B(KEYINPUT125), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(n969), .B(G21), .ZN(n970) );
  NAND2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n984) );
  XOR2_X1 U1066 ( .A(G1348), .B(KEYINPUT59), .Z(n972) );
  XNOR2_X1 U1067 ( .A(G4), .B(n972), .ZN(n980) );
  XNOR2_X1 U1068 ( .A(G1341), .B(G19), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(G1981), .B(G6), .ZN(n973) );
  NOR2_X1 U1070 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1071 ( .A(KEYINPUT122), .B(n975), .Z(n977) );
  XNOR2_X1 U1072 ( .A(G1956), .B(G20), .ZN(n976) );
  NOR2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1074 ( .A(n978), .B(KEYINPUT123), .ZN(n979) );
  NOR2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1076 ( .A(KEYINPUT60), .B(n981), .Z(n982) );
  XNOR2_X1 U1077 ( .A(KEYINPUT124), .B(n982), .ZN(n983) );
  NOR2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1079 ( .A(KEYINPUT126), .B(n985), .Z(n986) );
  NOR2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1081 ( .A(KEYINPUT61), .B(n988), .Z(n989) );
  NOR2_X1 U1082 ( .A1(G16), .A2(n989), .ZN(n1017) );
  XOR2_X1 U1083 ( .A(G16), .B(KEYINPUT56), .Z(n1015) );
  XNOR2_X1 U1084 ( .A(n990), .B(G1348), .ZN(n991) );
  XNOR2_X1 U1085 ( .A(n991), .B(KEYINPUT120), .ZN(n993) );
  NAND2_X1 U1086 ( .A1(G1971), .A2(G303), .ZN(n992) );
  NAND2_X1 U1087 ( .A1(n993), .A2(n992), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n1006) );
  XNOR2_X1 U1090 ( .A(n998), .B(G1341), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(G1966), .B(G168), .ZN(n1000) );
  NAND2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1093 ( .A(n1001), .B(KEYINPUT57), .ZN(n1002) );
  XNOR2_X1 U1094 ( .A(KEYINPUT119), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1013) );
  XNOR2_X1 U1097 ( .A(G1956), .B(G299), .ZN(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(G1961), .B(KEYINPUT121), .ZN(n1009) );
  XNOR2_X1 U1100 ( .A(n1009), .B(G301), .ZN(n1010) );
  NAND2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(n1018), .B(KEYINPUT127), .ZN(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1107 ( .A1(n1021), .A2(G11), .ZN(n1022) );
  XOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1022), .Z(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

