//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 1 0 0 1 1 1 1 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n849,
    new_n850, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT67), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT26), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n205), .B(new_n206), .C1(new_n204), .C2(new_n202), .ZN(new_n207));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT27), .B(G183gat), .ZN(new_n209));
  INV_X1    g008(.A(G190gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n207), .A2(new_n208), .A3(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n215), .B(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n218), .B(KEYINPUT65), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT24), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n208), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n217), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n202), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT23), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n202), .A2(KEYINPUT23), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n222), .A2(new_n225), .A3(new_n206), .A4(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT25), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n215), .A2(KEYINPUT68), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n230), .A2(new_n218), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n215), .A2(KEYINPUT68), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(new_n221), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n203), .A2(KEYINPUT23), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n206), .A2(KEYINPUT66), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n235), .B1(new_n224), .B2(new_n223), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n228), .B1(new_n206), .B2(KEYINPUT66), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n233), .A2(new_n234), .A3(new_n236), .A4(new_n237), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n229), .A2(KEYINPUT69), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT69), .B1(new_n229), .B2(new_n238), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n214), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(G120gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n242), .A2(G113gat), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT1), .B1(new_n243), .B2(KEYINPUT71), .ZN(new_n244));
  XNOR2_X1  g043(.A(G127gat), .B(G134gat), .ZN(new_n245));
  XOR2_X1   g044(.A(G113gat), .B(G120gat), .Z(new_n246));
  OAI211_X1 g045(.A(new_n244), .B(new_n245), .C1(new_n246), .C2(KEYINPUT71), .ZN(new_n247));
  INV_X1    g046(.A(new_n245), .ZN(new_n248));
  XNOR2_X1  g047(.A(G113gat), .B(G120gat), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n248), .B1(KEYINPUT1), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n241), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G227gat), .ZN(new_n254));
  INV_X1    g053(.A(G233gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n251), .B(new_n214), .C1(new_n239), .C2(new_n240), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n253), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G15gat), .B(G43gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(G71gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(G99gat), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT33), .ZN(new_n262));
  OR2_X1    g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n258), .A2(KEYINPUT32), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT73), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n258), .A2(KEYINPUT72), .A3(new_n262), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT72), .B1(new_n258), .B2(new_n262), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n261), .B1(new_n258), .B2(KEYINPUT32), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n265), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n258), .A2(new_n262), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT72), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n274), .A2(new_n270), .A3(new_n266), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n275), .A2(KEYINPUT73), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n264), .B1(new_n271), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n253), .A2(new_n257), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(new_n254), .B2(new_n255), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT34), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n264), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n269), .A2(new_n265), .A3(new_n270), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n275), .A2(KEYINPUT73), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n280), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G22gat), .B(G50gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT3), .ZN(new_n290));
  XNOR2_X1  g089(.A(G197gat), .B(G204gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(G211gat), .A2(G218gat), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n292), .A2(KEYINPUT22), .ZN(new_n293));
  NAND2_X1  g092(.A1(G211gat), .A2(G218gat), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n291), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(KEYINPUT74), .ZN(new_n297));
  AOI211_X1 g096(.A(new_n292), .B(new_n295), .C1(new_n291), .C2(KEYINPUT22), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n290), .B1(new_n299), .B2(KEYINPUT29), .ZN(new_n300));
  XOR2_X1   g099(.A(G141gat), .B(G148gat), .Z(new_n301));
  INV_X1    g100(.A(G155gat), .ZN(new_n302));
  INV_X1    g101(.A(G162gat), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT2), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G155gat), .B(G162gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n301), .A2(new_n306), .A3(new_n304), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n300), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G228gat), .A2(G233gat), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n313), .B1(new_n310), .B2(KEYINPUT3), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n311), .A2(new_n312), .A3(new_n315), .ZN(new_n316));
  AND3_X1   g115(.A1(new_n308), .A2(KEYINPUT77), .A3(new_n309), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT77), .B1(new_n308), .B2(new_n309), .ZN(new_n318));
  OR2_X1    g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n300), .A2(new_n319), .B1(new_n299), .B2(new_n314), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n316), .B1(new_n320), .B2(new_n312), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n321), .B(KEYINPUT31), .ZN(new_n322));
  XOR2_X1   g121(.A(G78gat), .B(G106gat), .Z(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n322), .A2(new_n323), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n289), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n326), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n328), .A2(new_n324), .A3(new_n288), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n281), .A2(new_n287), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT30), .ZN(new_n332));
  INV_X1    g131(.A(new_n299), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n229), .A2(new_n238), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n214), .ZN(new_n335));
  NAND2_X1  g134(.A1(G226gat), .A2(G233gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n337), .A2(KEYINPUT29), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n333), .B(new_n339), .C1(new_n241), .C2(new_n336), .ZN(new_n340));
  INV_X1    g139(.A(new_n335), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n241), .A2(new_n338), .B1(new_n341), .B2(new_n337), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n340), .B1(new_n342), .B2(new_n333), .ZN(new_n343));
  XNOR2_X1  g142(.A(G8gat), .B(G36gat), .ZN(new_n344));
  INV_X1    g143(.A(G64gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n346), .B(G92gat), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n343), .A2(KEYINPUT76), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT76), .B1(new_n343), .B2(new_n347), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n332), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT75), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n343), .A2(new_n347), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n352), .B1(new_n353), .B2(new_n332), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n343), .A2(KEYINPUT75), .A3(KEYINPUT30), .A4(new_n347), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OR2_X1    g155(.A1(new_n343), .A2(new_n347), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n351), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n251), .B1(new_n317), .B2(new_n318), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n310), .A2(new_n251), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  OAI211_X1 g162(.A(KEYINPUT78), .B(new_n251), .C1(new_n317), .C2(new_n318), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n361), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(G225gat), .A2(G233gat), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT3), .B1(new_n317), .B2(new_n318), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n369), .B(new_n251), .C1(KEYINPUT3), .C2(new_n310), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT4), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n362), .B(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n372), .A3(new_n366), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n368), .A2(KEYINPUT5), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT79), .ZN(new_n375));
  OR2_X1    g174(.A1(new_n373), .A2(KEYINPUT5), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n368), .A2(new_n377), .A3(new_n373), .A4(KEYINPUT5), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G1gat), .B(G29gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n380), .B(KEYINPUT0), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(G57gat), .ZN(new_n382));
  INV_X1    g181(.A(G85gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n382), .B(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n379), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT6), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n375), .A2(new_n384), .A3(new_n376), .A4(new_n378), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n379), .A2(KEYINPUT6), .A3(new_n385), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n358), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n392), .A2(KEYINPUT83), .ZN(new_n393));
  NOR2_X1   g192(.A1(KEYINPUT83), .A2(KEYINPUT35), .ZN(new_n394));
  NOR3_X1   g193(.A1(new_n358), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  NOR3_X1   g194(.A1(new_n331), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT84), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n331), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n281), .A2(new_n287), .A3(new_n330), .A4(KEYINPUT84), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n392), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n396), .B1(new_n400), .B2(KEYINPUT35), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT37), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n347), .B1(new_n343), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n403), .B1(new_n402), .B2(new_n343), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT38), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n339), .B1(new_n241), .B2(new_n336), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n299), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n241), .A2(new_n338), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n341), .A2(new_n337), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n409), .A3(new_n333), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n407), .A2(KEYINPUT37), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT81), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT38), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT81), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n407), .A2(new_n410), .A3(new_n414), .A4(KEYINPUT37), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n412), .A2(new_n403), .A3(new_n413), .A4(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT76), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n353), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n348), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n389), .A2(new_n416), .A3(new_n390), .A4(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT82), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n420), .A2(new_n421), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n405), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n370), .A2(new_n372), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n367), .ZN(new_n426));
  OR2_X1    g225(.A1(new_n426), .A2(KEYINPUT80), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(KEYINPUT80), .ZN(new_n428));
  OR2_X1    g227(.A1(new_n365), .A2(new_n367), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n427), .A2(new_n428), .A3(KEYINPUT39), .A4(new_n429), .ZN(new_n430));
  AND2_X1   g229(.A1(new_n427), .A2(new_n428), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n384), .B(new_n430), .C1(new_n431), .C2(KEYINPUT39), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(KEYINPUT40), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n433), .A2(new_n386), .A3(new_n358), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n424), .A2(new_n330), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT36), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n285), .A2(new_n286), .ZN(new_n437));
  AOI211_X1 g236(.A(new_n282), .B(new_n280), .C1(new_n283), .C2(new_n284), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n281), .A2(KEYINPUT36), .A3(new_n287), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OR2_X1    g240(.A1(new_n392), .A2(new_n330), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n435), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n401), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT9), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n445), .A2(G71gat), .A3(G78gat), .ZN(new_n446));
  AND2_X1   g245(.A1(G71gat), .A2(G78gat), .ZN(new_n447));
  INV_X1    g246(.A(G57gat), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n448), .A2(G64gat), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n345), .A2(G57gat), .ZN(new_n450));
  OAI22_X1  g249(.A1(new_n446), .A2(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n345), .A2(G57gat), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n448), .A2(G64gat), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n452), .A2(new_n453), .A3(KEYINPUT90), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT90), .B1(new_n452), .B2(new_n453), .ZN(new_n455));
  NOR3_X1   g254(.A1(new_n454), .A2(new_n455), .A3(new_n445), .ZN(new_n456));
  NOR2_X1   g255(.A1(G71gat), .A2(G78gat), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n447), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n451), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n461), .A2(KEYINPUT21), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n462), .B(G127gat), .ZN(new_n463));
  OR2_X1    g262(.A1(G15gat), .A2(G22gat), .ZN(new_n464));
  INV_X1    g263(.A(G1gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(G15gat), .A2(G22gat), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT88), .ZN(new_n468));
  AOI21_X1  g267(.A(G8gat), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n464), .A2(new_n466), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT16), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n471), .B1(new_n472), .B2(G1gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(new_n467), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n470), .B(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n475), .B1(KEYINPUT21), .B2(new_n461), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n463), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(G127gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n462), .B(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n476), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n483));
  XNOR2_X1  g282(.A(G155gat), .B(G183gat), .ZN(new_n484));
  XOR2_X1   g283(.A(new_n483), .B(new_n484), .Z(new_n485));
  NAND2_X1  g284(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(G231gat), .A2(G233gat), .ZN(new_n487));
  INV_X1    g286(.A(G211gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n485), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n478), .A2(new_n481), .A3(new_n490), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n486), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n489), .B1(new_n486), .B2(new_n491), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(G85gat), .A2(G92gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT7), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT7), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(G85gat), .A3(G92gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(G99gat), .A2(G106gat), .ZN(new_n500));
  INV_X1    g299(.A(G92gat), .ZN(new_n501));
  AOI22_X1  g300(.A1(KEYINPUT8), .A2(new_n500), .B1(new_n383), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(G99gat), .ZN(new_n503));
  INV_X1    g302(.A(G106gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n500), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n499), .A2(new_n502), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n506), .B1(new_n499), .B2(new_n502), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT92), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n509), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT92), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(new_n512), .A3(new_n507), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT14), .ZN(new_n515));
  INV_X1    g314(.A(G29gat), .ZN(new_n516));
  INV_X1    g315(.A(G36gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT87), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT87), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n520), .A2(new_n515), .A3(new_n516), .A4(new_n517), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n519), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  XOR2_X1   g322(.A(KEYINPUT86), .B(G29gat), .Z(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(G36gat), .ZN(new_n525));
  INV_X1    g324(.A(G50gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(G43gat), .ZN(new_n527));
  INV_X1    g326(.A(G43gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(G50gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT15), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n527), .A2(new_n529), .A3(KEYINPUT15), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n523), .A2(new_n525), .A3(new_n532), .A4(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n533), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT86), .B(G29gat), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n536), .A2(new_n517), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n535), .B(new_n518), .C1(new_n537), .C2(new_n522), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT17), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n534), .A2(new_n538), .A3(KEYINPUT17), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n514), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT93), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n511), .A2(new_n507), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(new_n539), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n514), .A2(KEYINPUT93), .A3(new_n541), .A4(new_n542), .ZN(new_n549));
  NAND2_X1  g348(.A1(G232gat), .A2(G233gat), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT41), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n545), .A2(new_n548), .A3(new_n549), .A4(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G190gat), .B(G218gat), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n554), .B(KEYINPUT94), .Z(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n543), .A2(new_n544), .B1(KEYINPUT41), .B2(new_n551), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n558), .A2(new_n555), .A3(new_n548), .A4(new_n549), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT95), .B1(new_n553), .B2(new_n556), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n551), .A2(KEYINPUT41), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT91), .ZN(new_n563));
  XOR2_X1   g362(.A(G134gat), .B(G162gat), .Z(new_n564));
  XOR2_X1   g363(.A(new_n563), .B(new_n564), .Z(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n560), .B1(new_n561), .B2(new_n566), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n557), .A2(KEYINPUT95), .A3(new_n559), .A4(new_n565), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(G230gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n570), .A2(new_n255), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT10), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n499), .A2(new_n502), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n505), .A2(KEYINPUT96), .A3(new_n500), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n506), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n576), .A2(new_n499), .A3(KEYINPUT96), .A4(new_n502), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT90), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n579), .B1(new_n449), .B2(new_n450), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n452), .A2(new_n453), .A3(KEYINPUT90), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n580), .A2(KEYINPUT9), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(new_n458), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT97), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n578), .A2(new_n583), .A3(new_n584), .A4(new_n451), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT97), .B1(new_n460), .B2(new_n546), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n578), .A2(new_n583), .A3(new_n451), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n572), .B(new_n585), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n461), .A2(KEYINPUT10), .A3(new_n547), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n571), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(new_n571), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G120gat), .B(G148gat), .ZN(new_n595));
  INV_X1    g394(.A(G176gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(G204gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n599), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n591), .A2(new_n593), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n494), .A2(new_n569), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(KEYINPUT98), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT98), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n494), .A2(new_n607), .A3(new_n569), .A4(new_n604), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n444), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n474), .B(new_n469), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n541), .A2(new_n611), .A3(new_n542), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n475), .A2(new_n539), .ZN(new_n613));
  NAND2_X1  g412(.A1(G229gat), .A2(G233gat), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT18), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n614), .B(KEYINPUT13), .Z(new_n618));
  INV_X1    g417(.A(new_n613), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n475), .A2(new_n539), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n612), .A2(new_n613), .A3(KEYINPUT18), .A4(new_n614), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n617), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT85), .ZN(new_n624));
  XNOR2_X1  g423(.A(G113gat), .B(G141gat), .ZN(new_n625));
  INV_X1    g424(.A(G197gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT11), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n625), .B(G197gat), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT11), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n628), .A2(new_n631), .A3(G169gat), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT12), .ZN(new_n634));
  AOI21_X1  g433(.A(G169gat), .B1(new_n628), .B2(new_n631), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(G169gat), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n629), .A2(new_n630), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n627), .A2(KEYINPUT11), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(KEYINPUT12), .B1(new_n640), .B2(new_n632), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n624), .B1(new_n636), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n634), .B1(new_n633), .B2(new_n635), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n640), .A2(KEYINPUT12), .A3(new_n632), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n643), .A2(KEYINPUT85), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n623), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(KEYINPUT89), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n636), .A2(new_n641), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n623), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT89), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n623), .A2(new_n646), .A3(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n648), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n610), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n391), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(new_n465), .ZN(G1324gat));
  INV_X1    g457(.A(new_n358), .ZN(new_n659));
  OR3_X1    g458(.A1(new_n655), .A2(KEYINPUT99), .A3(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT99), .B1(new_n655), .B2(new_n659), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT16), .B(G8gat), .Z(new_n662));
  NAND3_X1  g461(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT42), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n660), .A2(new_n661), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(G8gat), .ZN(new_n667));
  INV_X1    g466(.A(new_n655), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n668), .A2(KEYINPUT42), .A3(new_n358), .A4(new_n662), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n665), .A2(new_n667), .A3(new_n669), .ZN(G1325gat));
  INV_X1    g469(.A(G15gat), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n655), .A2(new_n671), .A3(new_n441), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n281), .A2(new_n287), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n668), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n672), .B1(new_n671), .B2(new_n675), .ZN(G1326gat));
  NOR2_X1   g475(.A1(new_n655), .A2(new_n330), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT43), .B(G22gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  INV_X1    g478(.A(new_n569), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n680), .B1(new_n401), .B2(new_n443), .ZN(new_n681));
  INV_X1    g480(.A(new_n654), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n494), .A2(new_n682), .A3(new_n603), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n685), .A2(new_n656), .A3(new_n524), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(KEYINPUT45), .Z(new_n687));
  NAND2_X1  g486(.A1(new_n681), .A2(KEYINPUT44), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n689), .B(new_n680), .C1(new_n401), .C2(new_n443), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n683), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT100), .B1(new_n692), .B2(new_n656), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT100), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n691), .A2(new_n694), .A3(new_n391), .A4(new_n683), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n693), .A2(new_n524), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n687), .A2(new_n696), .ZN(G1328gat));
  NOR3_X1   g496(.A1(new_n685), .A2(G36gat), .A3(new_n659), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT46), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT101), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n700), .B1(new_n692), .B2(new_n659), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n691), .A2(KEYINPUT101), .A3(new_n358), .A4(new_n683), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(G36gat), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n699), .A2(new_n703), .ZN(G1329gat));
  NOR2_X1   g503(.A1(new_n441), .A2(new_n528), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n691), .A2(new_n683), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n528), .B1(new_n685), .B2(new_n673), .ZN(new_n707));
  NAND2_X1  g506(.A1(KEYINPUT102), .A2(KEYINPUT47), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  OR2_X1    g508(.A1(KEYINPUT102), .A2(KEYINPUT47), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1330gat));
  INV_X1    g510(.A(new_n330), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n526), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n685), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n691), .A2(new_n712), .A3(new_n683), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n714), .B1(new_n715), .B2(G50gat), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT48), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n716), .A2(KEYINPUT103), .A3(new_n717), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n685), .A2(new_n713), .ZN(new_n719));
  AOI211_X1 g518(.A(new_n330), .B(new_n684), .C1(new_n688), .C2(new_n690), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n719), .B1(new_n720), .B2(new_n526), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT103), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT48), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n718), .A2(new_n723), .ZN(G1331gat));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n725));
  OR2_X1    g524(.A1(new_n492), .A2(new_n493), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(new_n680), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n727), .A2(new_n682), .A3(new_n603), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT104), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n725), .B1(new_n444), .B2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n729), .ZN(new_n731));
  OAI211_X1 g530(.A(KEYINPUT105), .B(new_n731), .C1(new_n401), .C2(new_n443), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n391), .ZN(new_n734));
  XNOR2_X1  g533(.A(KEYINPUT106), .B(G57gat), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1332gat));
  NAND2_X1  g535(.A1(new_n733), .A2(new_n358), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n738));
  XOR2_X1   g537(.A(KEYINPUT49), .B(G64gat), .Z(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n737), .B2(new_n739), .ZN(G1333gat));
  NAND3_X1  g539(.A1(new_n730), .A2(new_n674), .A3(new_n732), .ZN(new_n741));
  INV_X1    g540(.A(G71gat), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n441), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n730), .A2(G71gat), .A3(new_n744), .A4(new_n732), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n743), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT50), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n751), .B(new_n743), .C1(new_n747), .C2(new_n748), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(G1334gat));
  NAND2_X1  g552(.A1(new_n733), .A2(new_n712), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g554(.A1(new_n494), .A2(new_n654), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n680), .B(new_n756), .C1(new_n401), .C2(new_n443), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n757), .A2(KEYINPUT51), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(KEYINPUT51), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n758), .A2(new_n603), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n383), .B1(new_n760), .B2(new_n656), .ZN(new_n761));
  INV_X1    g560(.A(new_n756), .ZN(new_n762));
  AOI211_X1 g561(.A(new_n604), .B(new_n762), .C1(new_n688), .C2(new_n690), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n763), .A2(G85gat), .A3(new_n391), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT108), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n761), .A2(new_n764), .A3(KEYINPUT108), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(G1336gat));
  NOR3_X1   g568(.A1(new_n760), .A2(G92gat), .A3(new_n659), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n501), .B1(new_n763), .B2(new_n358), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT52), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n760), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n773), .A2(new_n501), .A3(new_n358), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n691), .A2(new_n603), .A3(new_n756), .ZN(new_n775));
  OAI21_X1  g574(.A(G92gat), .B1(new_n775), .B2(new_n659), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n774), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n772), .A2(new_n778), .ZN(G1337gat));
  OAI21_X1  g578(.A(G99gat), .B1(new_n775), .B2(new_n441), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n674), .A2(new_n503), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n780), .B1(new_n760), .B2(new_n781), .ZN(G1338gat));
  NOR3_X1   g581(.A1(new_n760), .A2(G106gat), .A3(new_n330), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n504), .B1(new_n763), .B2(new_n712), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT53), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n773), .A2(new_n504), .A3(new_n712), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n787));
  OAI21_X1  g586(.A(G106gat), .B1(new_n775), .B2(new_n330), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n785), .A2(new_n789), .ZN(G1339gat));
  INV_X1    g589(.A(KEYINPUT112), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT109), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n588), .A2(new_n589), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794));
  INV_X1    g593(.A(new_n571), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n588), .A2(new_n571), .A3(new_n589), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT54), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n599), .B(new_n796), .C1(new_n798), .C2(new_n590), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n792), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n591), .A2(KEYINPUT54), .A3(new_n797), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n601), .B1(new_n590), .B2(new_n794), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n802), .A2(new_n803), .A3(KEYINPUT109), .A4(KEYINPUT55), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n801), .A2(new_n602), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n799), .A2(new_n800), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n567), .A2(new_n806), .A3(new_n568), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT110), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n612), .A2(new_n613), .ZN(new_n810));
  INV_X1    g609(.A(new_n614), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI211_X1 g611(.A(KEYINPUT110), .B(new_n614), .C1(new_n612), .C2(new_n613), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OR2_X1    g613(.A1(new_n619), .A2(new_n620), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n815), .B2(new_n618), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n633), .A2(new_n635), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n650), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n805), .A2(new_n808), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(KEYINPUT111), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n603), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n654), .A2(new_n806), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n801), .A2(new_n602), .A3(new_n804), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n569), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n823), .A2(new_n807), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT111), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(new_n827), .A3(new_n818), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n820), .A2(new_n825), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n726), .ZN(new_n830));
  NOR4_X1   g629(.A1(new_n726), .A2(new_n680), .A3(new_n654), .A4(new_n603), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n791), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  AOI211_X1 g632(.A(KEYINPUT112), .B(new_n831), .C1(new_n829), .C2(new_n726), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n331), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n656), .A2(new_n358), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(G113gat), .B1(new_n838), .B2(new_n682), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT113), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n833), .A2(new_n834), .A3(new_n656), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n398), .A2(new_n399), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(new_n659), .A3(new_n842), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n682), .A2(G113gat), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n840), .B1(new_n843), .B2(new_n844), .ZN(G1340gat));
  OAI21_X1  g644(.A(G120gat), .B1(new_n838), .B2(new_n604), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n603), .A2(new_n242), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n846), .B1(new_n843), .B2(new_n847), .ZN(G1341gat));
  NOR3_X1   g647(.A1(new_n838), .A2(new_n479), .A3(new_n726), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n843), .A2(new_n726), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n849), .B1(new_n850), .B2(new_n479), .ZN(G1342gat));
  NOR3_X1   g650(.A1(new_n843), .A2(G134gat), .A3(new_n569), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT56), .ZN(new_n853));
  OAI21_X1  g652(.A(G134gat), .B1(new_n838), .B2(new_n569), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(G1343gat));
  INV_X1    g654(.A(KEYINPUT114), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n833), .A2(new_n834), .A3(new_n330), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(new_n857), .B2(KEYINPUT57), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n827), .B1(new_n826), .B2(new_n818), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n815), .A2(new_n618), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n860), .A2(new_n813), .A3(new_n812), .ZN(new_n861));
  INV_X1    g660(.A(new_n817), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n651), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NOR4_X1   g662(.A1(new_n823), .A2(new_n807), .A3(KEYINPUT111), .A4(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n494), .B1(new_n865), .B2(new_n825), .ZN(new_n866));
  OAI211_X1 g665(.A(KEYINPUT57), .B(new_n712), .C1(new_n866), .C2(new_n831), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT112), .B1(new_n866), .B2(new_n831), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n830), .A2(new_n791), .A3(new_n832), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n712), .A3(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(KEYINPUT114), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n858), .A2(new_n867), .A3(new_n872), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n441), .A2(new_n837), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n873), .A2(new_n654), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT116), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n873), .A2(new_n877), .A3(new_n654), .A4(new_n874), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n876), .A2(G141gat), .A3(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT58), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n744), .A2(new_n330), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n841), .A2(new_n659), .A3(new_n881), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n882), .A2(G141gat), .A3(new_n682), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n879), .A2(new_n880), .A3(new_n884), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n875), .A2(KEYINPUT115), .A3(G141gat), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT115), .B1(new_n875), .B2(G141gat), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n886), .A2(new_n887), .A3(new_n883), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n885), .B1(new_n888), .B2(new_n880), .ZN(G1344gat));
  NAND3_X1  g688(.A1(new_n873), .A2(new_n603), .A3(new_n874), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n890), .A2(new_n891), .A3(G148gat), .ZN(new_n892));
  XNOR2_X1  g691(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n826), .A2(KEYINPUT119), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n895), .B1(new_n823), .B2(new_n807), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n894), .A2(new_n818), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n494), .B1(new_n897), .B2(new_n825), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n654), .B1(new_n606), .B2(new_n608), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n871), .B(new_n712), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n901), .B1(new_n870), .B2(KEYINPUT57), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n603), .A3(new_n874), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n893), .B1(new_n903), .B2(G148gat), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT120), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(G148gat), .ZN(new_n907));
  AOI211_X1 g706(.A(new_n604), .B(new_n901), .C1(new_n870), .C2(KEYINPUT57), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(new_n874), .ZN(new_n909));
  OAI21_X1  g708(.A(KEYINPUT120), .B1(new_n909), .B2(new_n893), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n892), .A2(new_n906), .A3(new_n910), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n882), .A2(G148gat), .A3(new_n604), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT117), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT121), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT121), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n911), .A2(new_n916), .A3(new_n913), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(G1345gat));
  INV_X1    g717(.A(new_n882), .ZN(new_n919));
  AOI21_X1  g718(.A(G155gat), .B1(new_n919), .B2(new_n494), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n873), .A2(new_n874), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n726), .A2(new_n302), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(G1346gat));
  NAND3_X1  g722(.A1(new_n919), .A2(new_n303), .A3(new_n680), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n921), .A2(new_n680), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n924), .B1(new_n925), .B2(new_n303), .ZN(G1347gat));
  NAND2_X1  g725(.A1(new_n835), .A2(new_n656), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT122), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n835), .A2(KEYINPUT122), .A3(new_n656), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n931), .A2(new_n358), .A3(new_n842), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n637), .A3(new_n654), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n659), .A2(new_n391), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n835), .A2(new_n836), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(G169gat), .B1(new_n936), .B2(new_n682), .ZN(new_n937));
  XOR2_X1   g736(.A(new_n937), .B(KEYINPUT123), .Z(new_n938));
  NAND2_X1  g737(.A1(new_n934), .A2(new_n938), .ZN(G1348gat));
  NOR3_X1   g738(.A1(new_n936), .A2(new_n596), .A3(new_n604), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n933), .A2(new_n603), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n941), .B2(new_n596), .ZN(G1349gat));
  NAND3_X1  g741(.A1(new_n933), .A2(new_n209), .A3(new_n494), .ZN(new_n943));
  OAI21_X1  g742(.A(G183gat), .B1(new_n936), .B2(new_n726), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g745(.A(G190gat), .B1(new_n936), .B2(new_n569), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT61), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n680), .A2(new_n210), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n932), .B2(new_n949), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT124), .ZN(G1351gat));
  AND2_X1   g750(.A1(new_n931), .A2(new_n881), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n952), .A2(KEYINPUT125), .A3(new_n358), .ZN(new_n953));
  AOI21_X1  g752(.A(KEYINPUT125), .B1(new_n952), .B2(new_n358), .ZN(new_n954));
  OAI211_X1 g753(.A(new_n626), .B(new_n654), .C1(new_n953), .C2(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n902), .A2(new_n441), .A3(new_n935), .ZN(new_n956));
  OAI21_X1  g755(.A(G197gat), .B1(new_n956), .B2(new_n682), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(new_n957), .ZN(G1352gat));
  AND2_X1   g757(.A1(new_n952), .A2(new_n358), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n959), .A2(new_n598), .A3(new_n603), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(KEYINPUT62), .ZN(new_n961));
  INV_X1    g760(.A(new_n956), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n962), .A2(KEYINPUT126), .A3(new_n603), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n964), .B1(new_n956), .B2(new_n604), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n963), .A2(G204gat), .A3(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n959), .A2(new_n967), .A3(new_n598), .A4(new_n603), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n961), .A2(new_n966), .A3(new_n968), .ZN(G1353gat));
  OAI211_X1 g768(.A(new_n488), .B(new_n494), .C1(new_n953), .C2(new_n954), .ZN(new_n970));
  OAI21_X1  g769(.A(G211gat), .B1(new_n956), .B2(new_n726), .ZN(new_n971));
  XOR2_X1   g770(.A(new_n971), .B(KEYINPUT63), .Z(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(new_n972), .ZN(G1354gat));
  OAI21_X1  g772(.A(new_n680), .B1(new_n953), .B2(new_n954), .ZN(new_n974));
  INV_X1    g773(.A(G218gat), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n680), .A2(G218gat), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n976), .B(KEYINPUT127), .ZN(new_n977));
  AOI22_X1  g776(.A1(new_n974), .A2(new_n975), .B1(new_n962), .B2(new_n977), .ZN(G1355gat));
endmodule


