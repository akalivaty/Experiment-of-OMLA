//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n554, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n576, new_n577, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190,
    new_n1191, new_n1192, new_n1193;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT64), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT65), .Z(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  NAND3_X1  g033(.A1(new_n458), .A2(G101), .A3(G2104), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(KEYINPUT66), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(new_n458), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n459), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n458), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n468), .A2(new_n472), .ZN(G160));
  AOI21_X1  g048(.A(new_n458), .B1(new_n462), .B2(new_n464), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT67), .ZN(new_n476));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G112), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(new_n466), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G136), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n476), .A2(new_n481), .ZN(G162));
  NOR2_X1   g057(.A1(new_n458), .A2(G114), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n485), .B1(new_n474), .B2(G126), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n458), .A2(G138), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AND3_X1   g065(.A1(new_n469), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  AND3_X1   g066(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n492));
  AOI21_X1  g067(.A(KEYINPUT3), .B1(new_n463), .B2(G2104), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n490), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n491), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n494), .A2(KEYINPUT68), .A3(KEYINPUT4), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n487), .B1(new_n497), .B2(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n500));
  OR2_X1    g075(.A1(KEYINPUT69), .A2(G651), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT69), .A2(G651), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  OAI211_X1 g079(.A(G50), .B(G543), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  OR2_X1    g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g083(.A(G88), .B(new_n508), .C1(new_n503), .C2(new_n504), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT69), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT69), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G62), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n514), .B1(new_n506), .B2(new_n507), .ZN(new_n515));
  AND2_X1   g090(.A1(G75), .A2(G543), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n505), .A2(new_n509), .A3(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  AND2_X1   g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g097(.A(KEYINPUT6), .B1(new_n510), .B2(new_n511), .ZN(new_n523));
  INV_X1    g098(.A(new_n504), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G89), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n526), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G543), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n531), .B1(new_n523), .B2(new_n524), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT70), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n530), .B1(new_n533), .B2(G51), .ZN(G168));
  NAND2_X1  g109(.A1(new_n525), .A2(G90), .ZN(new_n535));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G64), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n522), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT71), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n513), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n508), .A2(G64), .ZN(new_n541));
  AOI21_X1  g116(.A(KEYINPUT71), .B1(new_n541), .B2(new_n536), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n535), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n543), .B1(G52), .B2(new_n533), .ZN(G171));
  NAND2_X1  g119(.A1(new_n533), .A2(G43), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT72), .B(G81), .Z(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n522), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n525), .A2(new_n546), .B1(new_n549), .B2(new_n513), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g128(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n554));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  OAI211_X1 g132(.A(G91), .B(new_n508), .C1(new_n503), .C2(new_n504), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(KEYINPUT75), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n525), .A2(new_n560), .A3(G91), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n522), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n559), .A2(new_n561), .B1(G651), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n532), .A2(G53), .A3(new_n566), .ZN(new_n567));
  OAI211_X1 g142(.A(G53), .B(G543), .C1(new_n503), .C2(new_n504), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n566), .ZN(new_n570));
  NOR2_X1   g145(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n567), .B1(new_n569), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n565), .A2(new_n573), .ZN(G299));
  INV_X1    g149(.A(G171), .ZN(G301));
  NAND2_X1  g150(.A1(new_n533), .A2(G51), .ZN(new_n576));
  INV_X1    g151(.A(new_n530), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(G286));
  NAND2_X1  g153(.A1(new_n523), .A2(new_n524), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n579), .A2(G49), .A3(G543), .ZN(new_n580));
  OAI211_X1 g155(.A(G87), .B(new_n508), .C1(new_n503), .C2(new_n504), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G288));
  NAND3_X1  g158(.A1(new_n579), .A2(G86), .A3(new_n508), .ZN(new_n584));
  OAI211_X1 g159(.A(G48), .B(G543), .C1(new_n503), .C2(new_n504), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AND2_X1   g161(.A1(G73), .A2(G543), .ZN(new_n587));
  OAI21_X1  g162(.A(G61), .B1(new_n520), .B2(new_n521), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n587), .B1(new_n588), .B2(KEYINPUT76), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n508), .A2(new_n590), .A3(G61), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n512), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n586), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G305));
  AOI22_X1  g169(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n595), .A2(new_n512), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT77), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n597), .B1(G85), .B2(new_n525), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n533), .A2(G47), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n525), .A2(G92), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT10), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n508), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G651), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n533), .A2(G54), .ZN(new_n608));
  AND2_X1   g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n601), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n601), .B1(new_n609), .B2(G868), .ZN(G321));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(G299), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(new_n612), .B2(G168), .ZN(G297));
  OAI21_X1  g189(.A(new_n613), .B1(new_n612), .B2(G168), .ZN(G280));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n609), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n609), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n619), .B(KEYINPUT78), .C1(G868), .C2(new_n551), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(KEYINPUT78), .B2(new_n619), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT79), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n480), .A2(G135), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n474), .A2(G123), .ZN(new_n625));
  OR2_X1    g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n626), .B(G2104), .C1(G111), .C2(new_n458), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(G2096), .Z(new_n629));
  NAND3_X1  g204(.A1(new_n458), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2100), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n629), .A2(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(KEYINPUT14), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT80), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n641), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(new_n649), .A3(G14), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(G401));
  INV_X1    g226(.A(KEYINPUT18), .ZN(new_n652));
  XOR2_X1   g227(.A(G2067), .B(G2678), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT81), .ZN(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(KEYINPUT17), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n652), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2072), .B(G2078), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT82), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n656), .B2(KEYINPUT18), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n659), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2096), .B(G2100), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  XOR2_X1   g242(.A(G1956), .B(G2474), .Z(new_n668));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  AND2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT20), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n668), .A2(new_n669), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n667), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n667), .B2(new_n673), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n676), .B(new_n677), .Z(new_n678));
  XNOR2_X1  g253(.A(G1991), .B(G1996), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(G229));
  NAND2_X1  g258(.A1(new_n480), .A2(G141), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n474), .A2(G129), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n458), .A2(G105), .A3(G2104), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT89), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  NAND3_X1  g264(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT26), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  AOI22_X1  g268(.A1(new_n688), .A2(new_n689), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n684), .A2(new_n685), .A3(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(G29), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n697), .B2(G32), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT27), .B(G1996), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT30), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n702), .A2(G28), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n697), .B1(new_n702), .B2(G28), .ZN(new_n704));
  AND2_X1   g279(.A1(KEYINPUT31), .A2(G11), .ZN(new_n705));
  NOR2_X1   g280(.A1(KEYINPUT31), .A2(G11), .ZN(new_n706));
  OAI22_X1  g281(.A1(new_n703), .A2(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n701), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n628), .A2(new_n697), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT92), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n699), .B2(new_n700), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT24), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n712), .A2(G34), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(G34), .ZN(new_n714));
  AOI21_X1  g289(.A(G29), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G160), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(G29), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G2084), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n697), .A2(G26), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT28), .Z(new_n720));
  NAND2_X1  g295(.A1(new_n474), .A2(G128), .ZN(new_n721));
  INV_X1    g296(.A(G140), .ZN(new_n722));
  NOR2_X1   g297(.A1(G104), .A2(G2105), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT87), .Z(new_n724));
  OAI21_X1  g299(.A(G2104), .B1(new_n458), .B2(G116), .ZN(new_n725));
  OAI221_X1 g300(.A(new_n721), .B1(new_n466), .B2(new_n722), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n720), .B1(new_n726), .B2(G29), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G2067), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n708), .A2(new_n711), .A3(new_n718), .A4(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n697), .A2(G35), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G162), .B2(new_n697), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT29), .Z(new_n732));
  INV_X1    g307(.A(G2090), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G1348), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n609), .A2(G16), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G4), .B2(G16), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n734), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  AOI211_X1 g313(.A(new_n729), .B(new_n738), .C1(new_n735), .C2(new_n737), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n732), .A2(new_n733), .ZN(new_n740));
  OAI21_X1  g315(.A(KEYINPUT90), .B1(G16), .B2(G21), .ZN(new_n741));
  NAND2_X1  g316(.A1(G168), .A2(G16), .ZN(new_n742));
  MUX2_X1   g317(.A(KEYINPUT90), .B(new_n741), .S(new_n742), .Z(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT91), .B(G1966), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n739), .B(new_n746), .C1(new_n744), .C2(new_n743), .ZN(new_n747));
  INV_X1    g322(.A(G16), .ZN(new_n748));
  NOR2_X1   g323(.A1(G171), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G5), .B2(new_n748), .ZN(new_n750));
  INV_X1    g325(.A(G1961), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(G164), .A2(G29), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G27), .B2(G29), .ZN(new_n754));
  INV_X1    g329(.A(G2078), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n697), .A2(G33), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT25), .Z(new_n760));
  INV_X1    g335(.A(G139), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n762));
  OAI221_X1 g337(.A(new_n760), .B1(new_n761), .B2(new_n466), .C1(new_n458), .C2(new_n762), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT88), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n758), .B1(new_n764), .B2(new_n697), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G2072), .ZN(new_n766));
  NOR2_X1   g341(.A1(G16), .A2(G19), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n551), .B2(G16), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(G1341), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n750), .B2(new_n751), .ZN(new_n770));
  OAI22_X1  g345(.A1(new_n768), .A2(G1341), .B1(new_n755), .B2(new_n754), .ZN(new_n771));
  NOR4_X1   g346(.A1(new_n757), .A2(new_n766), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT93), .B(KEYINPUT23), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT94), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n748), .A2(G20), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n774), .B(new_n775), .Z(new_n776));
  INV_X1    g351(.A(G299), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(new_n748), .ZN(new_n778));
  INV_X1    g353(.A(G1956), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n772), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n747), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT36), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n748), .A2(G24), .ZN(new_n785));
  INV_X1    g360(.A(G290), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(new_n748), .ZN(new_n787));
  INV_X1    g362(.A(G1986), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n697), .A2(G25), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n480), .A2(G131), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT83), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n794));
  INV_X1    g369(.A(G107), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(G2105), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n474), .B2(G119), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n790), .B1(new_n799), .B2(new_n697), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT35), .B(G1991), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT84), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n800), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n789), .A2(new_n803), .ZN(new_n804));
  MUX2_X1   g379(.A(G23), .B(G288), .S(G16), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT33), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G1976), .ZN(new_n807));
  NOR2_X1   g382(.A1(G6), .A2(G16), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n593), .B2(G16), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT32), .B(G1981), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n748), .A2(G22), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G166), .B2(new_n748), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G1971), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n811), .B1(KEYINPUT85), .B2(new_n814), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n807), .B(new_n815), .C1(KEYINPUT85), .C2(new_n814), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT86), .Z(new_n817));
  INV_X1    g392(.A(KEYINPUT34), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n804), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n816), .B(KEYINPUT86), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(KEYINPUT34), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n784), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n819), .A2(new_n784), .A3(new_n821), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n783), .B1(new_n823), .B2(new_n824), .ZN(G311));
  INV_X1    g400(.A(new_n824), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n782), .B1(new_n826), .B2(new_n822), .ZN(G150));
  NAND2_X1  g402(.A1(new_n607), .A2(new_n608), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n828), .A2(new_n616), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n533), .A2(G55), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n525), .A2(G93), .ZN(new_n833));
  NAND2_X1  g408(.A1(G80), .A2(G543), .ZN(new_n834));
  INV_X1    g409(.A(G67), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n522), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT96), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n513), .B1(new_n836), .B2(new_n837), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n833), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n832), .A2(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n841), .A2(new_n551), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n551), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n831), .B(new_n844), .Z(new_n845));
  OR2_X1    g420(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n846));
  INV_X1    g421(.A(G860), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n841), .A2(new_n847), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT37), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(G145));
  XOR2_X1   g427(.A(G160), .B(KEYINPUT97), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n628), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(G162), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n489), .B1(new_n462), .B2(new_n464), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n496), .B1(new_n856), .B2(new_n488), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n469), .A2(new_n488), .A3(new_n490), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n498), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(new_n486), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n726), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n695), .ZN(new_n862));
  INV_X1    g437(.A(new_n764), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n864), .B1(new_n763), .B2(new_n862), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n798), .B(new_n631), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n474), .A2(G130), .ZN(new_n867));
  OR2_X1    g442(.A1(G106), .A2(G2105), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n868), .B(G2104), .C1(G118), .C2(new_n458), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n870), .B1(G142), .B2(new_n480), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n866), .B(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n865), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT98), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n865), .A2(new_n872), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n873), .A2(new_n874), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n855), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(G37), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n855), .B(KEYINPUT99), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n881), .A2(new_n873), .A3(new_n876), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g459(.A1(KEYINPUT103), .A2(KEYINPUT42), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n609), .A2(G299), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n828), .A2(new_n777), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT41), .ZN(new_n889));
  OR3_X1    g464(.A1(new_n888), .A2(KEYINPUT101), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(KEYINPUT101), .B1(new_n888), .B2(new_n889), .ZN(new_n891));
  AOI21_X1  g466(.A(KEYINPUT100), .B1(new_n888), .B2(new_n889), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n888), .A2(KEYINPUT100), .A3(new_n889), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n890), .B(new_n891), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n844), .B(new_n618), .Z(new_n895));
  AND2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n888), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n885), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(G288), .B(KEYINPUT102), .ZN(new_n900));
  XNOR2_X1  g475(.A(G290), .B(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n593), .B(G166), .ZN(new_n902));
  XOR2_X1   g477(.A(new_n901), .B(new_n902), .Z(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n904), .B1(KEYINPUT103), .B2(KEYINPUT42), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n894), .A2(new_n895), .ZN(new_n906));
  INV_X1    g481(.A(new_n885), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n906), .B(new_n907), .C1(new_n895), .C2(new_n897), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n899), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n905), .B1(new_n899), .B2(new_n908), .ZN(new_n910));
  OAI21_X1  g485(.A(G868), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n612), .B1(new_n832), .B2(new_n840), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(G295));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n912), .ZN(G331));
  XOR2_X1   g489(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n915));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n916));
  XNOR2_X1  g491(.A(G286), .B(G171), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n844), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n917), .A2(new_n842), .A3(new_n843), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n894), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n919), .A2(new_n923), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n920), .A2(new_n888), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n917), .B1(new_n842), .B2(new_n843), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT105), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n903), .B1(new_n922), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n928), .B1(new_n894), .B2(new_n921), .ZN(new_n930));
  AOI21_X1  g505(.A(G37), .B1(new_n930), .B2(new_n904), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n916), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  AOI211_X1 g507(.A(new_n928), .B(new_n903), .C1(new_n894), .C2(new_n921), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n924), .A2(new_n927), .A3(new_n920), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n888), .B(new_n889), .ZN(new_n935));
  AOI22_X1  g510(.A1(new_n934), .A2(new_n935), .B1(new_n919), .B2(new_n925), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n880), .B1(new_n936), .B2(new_n904), .ZN(new_n937));
  NOR3_X1   g512(.A1(new_n933), .A2(new_n937), .A3(KEYINPUT43), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n915), .B1(new_n932), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n929), .A2(new_n931), .A3(new_n916), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT43), .B1(new_n933), .B2(new_n937), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(new_n941), .A3(KEYINPUT44), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n939), .A2(new_n942), .ZN(G397));
  INV_X1    g518(.A(KEYINPUT45), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n944), .B1(G164), .B2(G1384), .ZN(new_n945));
  INV_X1    g520(.A(G40), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n468), .A2(new_n472), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n786), .A2(new_n950), .A3(new_n788), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n950), .A2(G290), .A3(G1986), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT106), .ZN(new_n954));
  XOR2_X1   g529(.A(new_n695), .B(G1996), .Z(new_n955));
  INV_X1    g530(.A(G2067), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n726), .B(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n949), .ZN(new_n959));
  XOR2_X1   g534(.A(new_n959), .B(KEYINPUT107), .Z(new_n960));
  NAND2_X1  g535(.A1(new_n799), .A2(new_n802), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n799), .A2(new_n802), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n949), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n960), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n954), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT63), .ZN(new_n967));
  NAND3_X1  g542(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT108), .ZN(new_n969));
  NAND2_X1  g544(.A1(G303), .A2(G8), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT55), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n973));
  NAND4_X1  g548(.A1(G303), .A2(new_n973), .A3(KEYINPUT55), .A4(G8), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n969), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G1971), .ZN(new_n977));
  AOI21_X1  g552(.A(G1384), .B1(new_n859), .B2(new_n486), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n947), .B1(new_n978), .B2(KEYINPUT45), .ZN(new_n979));
  AOI211_X1 g554(.A(new_n944), .B(G1384), .C1(new_n859), .C2(new_n486), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n977), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n978), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n982), .A2(new_n733), .A3(new_n947), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n976), .B1(new_n986), .B2(G8), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n986), .A2(G8), .A3(new_n976), .ZN(new_n989));
  INV_X1    g564(.A(G8), .ZN(new_n990));
  AND4_X1   g565(.A1(G1976), .A2(new_n580), .A3(new_n581), .A4(new_n582), .ZN(new_n991));
  AOI211_X1 g566(.A(new_n990), .B(new_n991), .C1(new_n978), .C2(new_n947), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT109), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n990), .B1(new_n978), .B2(new_n947), .ZN(new_n995));
  INV_X1    g570(.A(new_n991), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(new_n998), .A3(KEYINPUT52), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n994), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G1976), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT52), .B1(G288), .B2(new_n1001), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n995), .A2(new_n996), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT49), .ZN(new_n1004));
  INV_X1    g579(.A(G1981), .ZN(new_n1005));
  AOI22_X1  g580(.A1(G48), .A2(new_n532), .B1(new_n525), .B2(G86), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n589), .A2(new_n591), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n513), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1005), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n586), .A2(new_n592), .A3(G1981), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1004), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1006), .A2(new_n1008), .A3(new_n1005), .ZN(new_n1012));
  OAI21_X1  g587(.A(G1981), .B1(new_n586), .B2(new_n592), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1012), .A2(new_n1013), .A3(KEYINPUT49), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1011), .A2(new_n995), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT110), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT110), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1011), .A2(new_n995), .A3(new_n1017), .A4(new_n1014), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1003), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n988), .A2(new_n989), .A3(new_n1000), .A4(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1384), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n860), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n948), .B1(new_n1022), .B2(KEYINPUT50), .ZN(new_n1023));
  INV_X1    g598(.A(G2084), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1023), .A2(new_n1024), .A3(new_n984), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n744), .B1(new_n979), .B2(new_n980), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n990), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(G168), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n967), .B1(new_n1020), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1003), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1031), .A2(new_n1000), .A3(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1030), .B1(new_n1033), .B2(new_n987), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n988), .A2(KEYINPUT112), .A3(new_n1000), .A4(new_n1019), .ZN(new_n1035));
  AOI211_X1 g610(.A(new_n990), .B(new_n975), .C1(new_n981), .C2(new_n985), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n1028), .A2(new_n1036), .A3(new_n967), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  OR2_X1    g613(.A1(G288), .A2(G1976), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1039), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n995), .B1(new_n1040), .B2(new_n1010), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1019), .A2(new_n1036), .A3(new_n1000), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1041), .A2(new_n1042), .A3(KEYINPUT111), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1029), .A2(new_n1038), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n568), .A2(new_n570), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n572), .B1(new_n532), .B2(G53), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT114), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n567), .B(new_n1051), .C1(new_n569), .C2(new_n572), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1050), .A2(new_n565), .A3(new_n1052), .ZN(new_n1053));
  XOR2_X1   g628(.A(KEYINPUT113), .B(KEYINPUT57), .Z(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n565), .A2(KEYINPUT57), .A3(new_n573), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n947), .B1(new_n978), .B2(new_n983), .ZN(new_n1058));
  AOI211_X1 g633(.A(KEYINPUT50), .B(G1384), .C1(new_n859), .C2(new_n486), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n779), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n978), .A2(KEYINPUT45), .ZN(new_n1061));
  XNOR2_X1  g636(.A(KEYINPUT56), .B(G2072), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n945), .A2(new_n947), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1057), .A2(new_n1060), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1057), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT117), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1057), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n978), .A2(KEYINPUT115), .A3(new_n947), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT115), .B1(new_n978), .B2(new_n947), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n956), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n735), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT116), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(KEYINPUT116), .A3(new_n1077), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1079), .A2(new_n609), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1065), .B1(new_n1073), .B2(new_n1081), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1064), .A2(KEYINPUT61), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1069), .A2(new_n1083), .A3(new_n1072), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1080), .ZN(new_n1085));
  OAI211_X1 g660(.A(KEYINPUT60), .B(new_n828), .C1(new_n1085), .C2(new_n1078), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT61), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(new_n1065), .B2(new_n1070), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT58), .B(G1341), .ZN(new_n1089));
  NOR3_X1   g664(.A1(new_n1074), .A2(new_n1075), .A3(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT118), .B(G1996), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n979), .A2(new_n980), .A3(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n551), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT59), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT59), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1095), .B(new_n551), .C1(new_n1090), .C2(new_n1092), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  AND4_X1   g672(.A1(new_n1084), .A2(new_n1086), .A3(new_n1088), .A4(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT60), .B1(new_n1085), .B2(new_n1078), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT60), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1079), .A2(new_n1080), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1099), .A2(new_n1101), .A3(new_n609), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1082), .B1(new_n1098), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1105), .A2(G2078), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n979), .A2(new_n980), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1023), .A2(new_n984), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1108), .A2(new_n1109), .B1(new_n1110), .B2(new_n751), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n948), .B1(new_n1022), .B2(new_n944), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1112), .A2(new_n755), .A3(new_n1061), .ZN(new_n1113));
  AOI21_X1  g688(.A(G171), .B1(new_n1113), .B2(new_n1105), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT122), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1112), .A2(new_n1061), .A3(new_n1106), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT121), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1111), .A2(new_n1114), .A3(new_n1115), .A4(new_n1117), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1113), .A2(new_n1105), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n751), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1116), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(G171), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1120), .B1(new_n1116), .B2(KEYINPUT121), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1115), .B1(new_n1126), .B2(new_n1114), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1104), .B1(new_n1123), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(G8), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n1131));
  NAND3_X1  g706(.A1(G286), .A2(new_n1131), .A3(G8), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT119), .B1(G168), .B2(new_n990), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT51), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1130), .B(new_n1134), .C1(KEYINPUT120), .C2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1129), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1138), .B1(new_n1027), .B2(new_n1137), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT120), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT51), .B1(new_n1027), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1136), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1111), .A2(new_n1117), .ZN(new_n1144));
  OAI21_X1  g719(.A(G171), .B1(new_n1144), .B2(new_n1119), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1113), .A2(new_n1105), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1146), .A2(G301), .A3(new_n1116), .A4(new_n1120), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1145), .A2(KEYINPUT54), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1020), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1128), .A2(new_n1143), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1047), .B(KEYINPUT123), .C1(new_n1103), .C2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT62), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1142), .A2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1136), .B(KEYINPUT62), .C1(new_n1139), .C2(new_n1141), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1020), .A2(new_n1122), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(KEYINPUT124), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT124), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1153), .A2(new_n1155), .A3(new_n1158), .A4(new_n1154), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1151), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1147), .A2(KEYINPUT54), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1126), .A2(new_n1146), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1162), .B1(new_n1163), .B2(G171), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1164), .A2(new_n1142), .A3(new_n1020), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1084), .A2(new_n1086), .A3(new_n1097), .A4(new_n1088), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1099), .A2(new_n1101), .A3(new_n609), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1165), .B(new_n1128), .C1(new_n1168), .C2(new_n1082), .ZN(new_n1169));
  AOI21_X1  g744(.A(KEYINPUT123), .B1(new_n1169), .B2(new_n1047), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n966), .B1(new_n1161), .B2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n950), .A2(G1996), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT46), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n957), .A2(new_n696), .ZN(new_n1175));
  AOI22_X1  g750(.A1(new_n1173), .A2(new_n1174), .B1(new_n949), .B2(new_n1175), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n1173), .A2(KEYINPUT125), .A3(new_n1174), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT125), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1178), .B1(new_n1172), .B2(KEYINPUT46), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1176), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  XOR2_X1   g755(.A(new_n1180), .B(KEYINPUT47), .Z(new_n1181));
  XNOR2_X1  g756(.A(new_n952), .B(KEYINPUT48), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n965), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n960), .A2(new_n962), .ZN(new_n1184));
  OR2_X1    g759(.A1(new_n726), .A2(G2067), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n950), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NOR3_X1   g761(.A1(new_n1181), .A2(new_n1183), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1171), .A2(new_n1187), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g763(.A(G319), .ZN(new_n1190));
  NOR2_X1   g764(.A1(G227), .A2(new_n1190), .ZN(new_n1191));
  XOR2_X1   g765(.A(new_n1191), .B(KEYINPUT126), .Z(new_n1192));
  NOR3_X1   g766(.A1(G229), .A2(G401), .A3(new_n1192), .ZN(new_n1193));
  OAI211_X1 g767(.A(new_n883), .B(new_n1193), .C1(new_n932), .C2(new_n938), .ZN(G225));
  INV_X1    g768(.A(G225), .ZN(G308));
endmodule


