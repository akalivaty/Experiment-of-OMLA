//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 0 1 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n786, new_n787, new_n788, new_n789, new_n791, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982;
  INV_X1    g000(.A(KEYINPUT94), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n203));
  XNOR2_X1  g002(.A(G113gat), .B(G141gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G169gat), .B(G197gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n207), .B(KEYINPUT12), .ZN(new_n208));
  XOR2_X1   g007(.A(new_n208), .B(KEYINPUT86), .Z(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G15gat), .B(G22gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT16), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n211), .B1(new_n212), .B2(G1gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT88), .ZN(new_n214));
  INV_X1    g013(.A(G15gat), .ZN(new_n215));
  INV_X1    g014(.A(G22gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G1gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(G15gat), .A2(G22gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n213), .A2(new_n214), .A3(new_n220), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n211), .B(KEYINPUT88), .C1(new_n212), .C2(G1gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(G8gat), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n213), .A2(KEYINPUT89), .ZN(new_n224));
  INV_X1    g023(.A(G8gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT89), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n211), .B(new_n226), .C1(new_n212), .C2(G1gat), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n224), .A2(new_n225), .A3(new_n220), .A4(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT17), .ZN(new_n231));
  XOR2_X1   g030(.A(G43gat), .B(G50gat), .Z(new_n232));
  INV_X1    g031(.A(KEYINPUT15), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT14), .ZN(new_n235));
  NOR3_X1   g034(.A1(new_n235), .A2(G29gat), .A3(G36gat), .ZN(new_n236));
  INV_X1    g035(.A(G29gat), .ZN(new_n237));
  INV_X1    g036(.A(G36gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G29gat), .A2(G36gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT14), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n236), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G43gat), .B(G50gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT15), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n234), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n241), .A2(new_n239), .ZN(new_n246));
  OAI211_X1 g045(.A(KEYINPUT15), .B(new_n243), .C1(new_n246), .C2(new_n236), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT87), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT87), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n231), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n250), .B1(new_n245), .B2(new_n247), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n243), .B(new_n233), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT87), .B1(new_n254), .B2(new_n242), .ZN(new_n255));
  NOR3_X1   g054(.A1(new_n253), .A2(new_n255), .A3(KEYINPUT17), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n230), .B1(new_n252), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n253), .A2(new_n255), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT90), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n223), .A2(new_n228), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n260), .B1(new_n223), .B2(new_n228), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n259), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G229gat), .A2(G233gat), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n257), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT91), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT18), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n267), .B1(new_n266), .B2(new_n268), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AND3_X1   g070(.A1(new_n257), .A2(new_n264), .A3(new_n265), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n229), .A2(KEYINPUT90), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n273), .A2(new_n261), .A3(new_n258), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT93), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT93), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n273), .A2(new_n276), .A3(new_n261), .A4(new_n258), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n275), .A2(new_n264), .A3(new_n277), .ZN(new_n278));
  XOR2_X1   g077(.A(new_n265), .B(KEYINPUT92), .Z(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT13), .ZN(new_n280));
  AOI22_X1  g079(.A1(KEYINPUT18), .A2(new_n272), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n210), .B1(new_n271), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n268), .ZN(new_n283));
  AND3_X1   g082(.A1(new_n281), .A2(new_n208), .A3(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n202), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(KEYINPUT91), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n278), .A2(new_n280), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT18), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n286), .A2(new_n287), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(new_n209), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n281), .A2(new_n208), .A3(new_n283), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n291), .A2(KEYINPUT94), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n285), .A2(new_n293), .ZN(new_n294));
  AND2_X1   g093(.A1(G227gat), .A2(G233gat), .ZN(new_n295));
  INV_X1    g094(.A(G190gat), .ZN(new_n296));
  AND2_X1   g095(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT28), .ZN(new_n300));
  OR3_X1    g099(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302));
  OAI21_X1  g101(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G183gat), .A2(G190gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT28), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n306), .B(new_n296), .C1(new_n297), .C2(new_n298), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n300), .A2(new_n304), .A3(new_n305), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n302), .B1(new_n309), .B2(G190gat), .ZN(new_n310));
  OR2_X1    g109(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n296), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT23), .ZN(new_n314));
  INV_X1    g113(.A(G169gat), .ZN(new_n315));
  INV_X1    g114(.A(G176gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT25), .B1(new_n313), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n310), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n311), .A2(G190gat), .A3(new_n309), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n321), .A2(new_n319), .A3(new_n322), .A4(KEYINPUT25), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n308), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G134gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(G113gat), .B(G120gat), .ZN(new_n327));
  NOR3_X1   g126(.A1(new_n327), .A2(KEYINPUT1), .A3(G127gat), .ZN(new_n328));
  INV_X1    g127(.A(G127gat), .ZN(new_n329));
  INV_X1    g128(.A(G120gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(G113gat), .ZN(new_n331));
  INV_X1    g130(.A(G113gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G120gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT1), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n329), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n326), .B1(new_n328), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(G127gat), .B1(new_n327), .B2(KEYINPUT1), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n334), .A2(new_n335), .A3(new_n329), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(new_n339), .A3(G134gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n321), .A2(new_n319), .A3(new_n322), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT25), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(new_n323), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n346), .A2(new_n308), .B1(new_n337), .B2(new_n340), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n295), .B1(new_n342), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G15gat), .B(G43gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n349), .B(G71gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(G99gat), .ZN(new_n351));
  INV_X1    g150(.A(G71gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n349), .B(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G99gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT64), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT64), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n351), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(KEYINPUT33), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n348), .A2(KEYINPUT32), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n325), .A2(new_n341), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n346), .A2(new_n340), .A3(new_n337), .A4(new_n308), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT32), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n364), .A2(new_n295), .B1(new_n365), .B2(KEYINPUT33), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n361), .B1(new_n366), .B2(new_n356), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT34), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n364), .A2(new_n295), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT34), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n361), .B(new_n370), .C1(new_n356), .C2(new_n366), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n368), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n369), .B1(new_n368), .B2(new_n371), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT6), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT70), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n338), .A2(new_n339), .A3(G134gat), .ZN(new_n377));
  AOI21_X1  g176(.A(G134gat), .B1(new_n338), .B2(new_n339), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n337), .A2(KEYINPUT70), .A3(new_n340), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT69), .B(G155gat), .ZN(new_n381));
  INV_X1    g180(.A(G162gat), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT2), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(G148gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(G141gat), .ZN(new_n385));
  INV_X1    g184(.A(G141gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(G148gat), .ZN(new_n387));
  OR2_X1    g186(.A1(G155gat), .A2(G162gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(G155gat), .A2(G162gat), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n385), .A2(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n383), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(KEYINPUT2), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n386), .A2(G148gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n384), .A2(G141gat), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n389), .ZN(new_n396));
  NOR2_X1   g195(.A1(G155gat), .A2(G162gat), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n396), .A2(new_n397), .A3(KEYINPUT68), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT68), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n399), .B1(new_n388), .B2(new_n389), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n395), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n391), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT3), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT3), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n391), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n379), .A2(new_n380), .A3(new_n403), .A4(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(G225gat), .A2(G233gat), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n337), .A2(new_n340), .A3(new_n401), .A4(new_n391), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n377), .A2(new_n378), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n391), .A2(new_n401), .A3(KEYINPUT71), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT71), .B1(new_n391), .B2(new_n401), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n412), .B(KEYINPUT4), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n406), .A2(new_n411), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n379), .A2(new_n380), .A3(new_n402), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n418), .A2(new_n409), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n417), .B(KEYINPUT5), .C1(new_n419), .C2(new_n407), .ZN(new_n420));
  INV_X1    g219(.A(new_n415), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n413), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n412), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n410), .ZN(new_n424));
  OR2_X1    g223(.A1(new_n409), .A2(new_n410), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n408), .A2(KEYINPUT5), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n424), .A2(new_n406), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n420), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(KEYINPUT72), .B(KEYINPUT0), .ZN(new_n429));
  XNOR2_X1  g228(.A(G1gat), .B(G29gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n429), .B(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(G57gat), .B(G85gat), .ZN(new_n432));
  XOR2_X1   g231(.A(new_n431), .B(new_n432), .Z(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n375), .B1(new_n428), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n428), .A2(new_n434), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n437), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n435), .ZN(new_n440));
  INV_X1    g239(.A(G211gat), .ZN(new_n441));
  INV_X1    g240(.A(G218gat), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g242(.A1(G211gat), .A2(G218gat), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(KEYINPUT65), .B(G211gat), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT22), .B1(new_n446), .B2(G218gat), .ZN(new_n447));
  INV_X1    g246(.A(G197gat), .ZN(new_n448));
  INV_X1    g247(.A(G204gat), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(G197gat), .A2(G204gat), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n445), .B1(new_n447), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n445), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n441), .A2(KEYINPUT65), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT65), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(G211gat), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n455), .A2(new_n457), .A3(G218gat), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT22), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OR2_X1    g259(.A1(new_n450), .A2(new_n451), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n454), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  AND2_X1   g261(.A1(new_n453), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT67), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT29), .B1(new_n346), .B2(new_n308), .ZN(new_n466));
  NAND2_X1  g265(.A1(G226gat), .A2(G233gat), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n465), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n467), .B1(new_n346), .B2(new_n308), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT29), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n325), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n470), .B1(new_n472), .B2(new_n467), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n464), .B(new_n469), .C1(new_n473), .C2(new_n465), .ZN(new_n474));
  NOR3_X1   g273(.A1(new_n473), .A2(KEYINPUT66), .A3(new_n464), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT66), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n325), .A2(new_n468), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n477), .B1(new_n466), .B2(new_n468), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n476), .B1(new_n478), .B2(new_n463), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n474), .B1(new_n475), .B2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(G8gat), .B(G36gat), .ZN(new_n481));
  INV_X1    g280(.A(G64gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(G92gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(new_n484), .ZN(new_n485));
  OR3_X1    g284(.A1(new_n480), .A2(KEYINPUT30), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n480), .A2(new_n485), .ZN(new_n487));
  INV_X1    g286(.A(new_n485), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n474), .B(new_n488), .C1(new_n475), .C2(new_n479), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n487), .A2(KEYINPUT30), .A3(new_n489), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n438), .A2(new_n440), .B1(new_n486), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT29), .B1(new_n453), .B2(new_n462), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n402), .B1(new_n492), .B2(KEYINPUT3), .ZN(new_n493));
  NAND2_X1  g292(.A1(G228gat), .A2(G233gat), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n405), .A2(new_n471), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n463), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n493), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT74), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT74), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n493), .A2(new_n497), .A3(new_n500), .A4(new_n495), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n453), .A2(new_n462), .A3(KEYINPUT73), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT73), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n504), .B(new_n445), .C1(new_n447), .C2(new_n452), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n471), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n422), .B1(new_n404), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n497), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n494), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n502), .A2(new_n509), .A3(new_n216), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT75), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  XOR2_X1   g311(.A(G78gat), .B(G106gat), .Z(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(KEYINPUT31), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(G50gat), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n502), .A2(new_n509), .A3(KEYINPUT75), .A4(new_n216), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n512), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT76), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n502), .A2(new_n509), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(G22gat), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n520), .B1(new_n522), .B2(new_n510), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n216), .B1(new_n502), .B2(new_n509), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n524), .A2(new_n519), .ZN(new_n525));
  OAI211_X1 g324(.A(KEYINPUT77), .B(new_n517), .C1(new_n523), .C2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n502), .A2(new_n216), .A3(new_n509), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n519), .B1(new_n528), .B2(new_n524), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n522), .A2(new_n520), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT77), .B1(new_n531), .B2(new_n517), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n374), .B(new_n491), .C1(new_n527), .C2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT35), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT84), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n527), .A2(new_n532), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n420), .A2(KEYINPUT82), .A3(new_n427), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT82), .B1(new_n420), .B2(new_n427), .ZN(new_n538));
  NOR3_X1   g337(.A1(new_n537), .A2(new_n538), .A3(new_n433), .ZN(new_n539));
  OAI22_X1  g338(.A1(new_n539), .A2(new_n435), .B1(new_n375), .B2(new_n437), .ZN(new_n540));
  NOR3_X1   g339(.A1(new_n372), .A2(new_n373), .A3(KEYINPUT35), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n490), .A2(new_n486), .A3(KEYINPUT78), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT78), .B1(new_n490), .B2(new_n486), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n540), .B(new_n541), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n535), .B1(new_n536), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n517), .B1(new_n523), .B2(new_n525), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT77), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(new_n526), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n540), .A2(new_n541), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n490), .A2(new_n486), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT78), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n490), .A2(new_n486), .A3(KEYINPUT78), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n549), .A2(new_n550), .A3(KEYINPUT84), .A4(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n534), .A2(new_n545), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n491), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n536), .A2(new_n558), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n374), .A2(KEYINPUT36), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n374), .A2(KEYINPUT36), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n538), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n420), .A2(new_n427), .A3(KEYINPUT82), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n434), .A3(new_n564), .ZN(new_n565));
  AOI22_X1  g364(.A1(new_n565), .A2(new_n436), .B1(new_n439), .B2(KEYINPUT6), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n473), .A2(new_n464), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT83), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n478), .A2(KEYINPUT67), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n464), .B1(new_n569), .B2(new_n469), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT37), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  OR2_X1    g370(.A1(new_n480), .A2(KEYINPUT37), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT38), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n571), .A2(new_n572), .A3(new_n573), .A4(new_n485), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n480), .A2(KEYINPUT37), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n485), .B1(new_n480), .B2(KEYINPUT37), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT38), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n566), .A2(new_n489), .A3(new_n574), .A4(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n549), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n424), .A2(new_n406), .A3(new_n425), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(new_n408), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n418), .A2(new_n407), .A3(new_n409), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT39), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT79), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n582), .A2(KEYINPUT79), .A3(KEYINPUT39), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n581), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n587), .A2(new_n433), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT39), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n580), .A2(new_n589), .A3(new_n408), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT81), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT40), .ZN(new_n592));
  AOI22_X1  g391(.A1(new_n588), .A2(new_n590), .B1(KEYINPUT80), .B2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n587), .A2(KEYINPUT80), .A3(new_n433), .A4(new_n590), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT40), .B1(new_n594), .B2(new_n591), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n565), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n596), .A2(new_n555), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n559), .B(new_n562), .C1(new_n579), .C2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n294), .B1(new_n557), .B2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G183gat), .B(G211gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT98), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT19), .ZN(new_n602));
  XOR2_X1   g401(.A(G127gat), .B(G155gat), .Z(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT20), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n602), .B(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G57gat), .B(G64gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT95), .ZN(new_n608));
  AOI21_X1  g407(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G71gat), .B(G78gat), .Z(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(new_n609), .ZN(new_n614));
  INV_X1    g413(.A(G57gat), .ZN(new_n615));
  OR2_X1    g414(.A1(KEYINPUT96), .A2(G64gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(KEYINPUT96), .A2(G64gat), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT97), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(KEYINPUT97), .B1(new_n482), .B2(G57gat), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n614), .B(new_n620), .C1(new_n618), .C2(new_n621), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n613), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT21), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT99), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n624), .A2(new_n625), .A3(new_n273), .A4(new_n261), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT21), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n613), .A2(new_n622), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n273), .B(new_n261), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT99), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n626), .A2(new_n630), .A3(G231gat), .A4(G233gat), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n623), .A2(KEYINPUT21), .ZN(new_n633));
  AOI22_X1  g432(.A1(new_n626), .A2(new_n630), .B1(G231gat), .B2(G233gat), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n633), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n626), .A2(new_n630), .ZN(new_n637));
  INV_X1    g436(.A(G231gat), .ZN(new_n638));
  INV_X1    g437(.A(G233gat), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n636), .B1(new_n640), .B2(new_n631), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n606), .B1(new_n635), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n633), .B1(new_n632), .B2(new_n634), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n640), .A2(new_n636), .A3(new_n631), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n643), .A2(new_n644), .A3(new_n605), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  OR2_X1    g445(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n647));
  NAND2_X1  g446(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n647), .A2(G85gat), .A3(G92gat), .A4(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(G85gat), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n484), .ZN(new_n651));
  NOR2_X1   g450(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n652));
  NAND2_X1  g451(.A1(G85gat), .A2(G92gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(G99gat), .A2(G106gat), .ZN(new_n654));
  AOI22_X1  g453(.A1(new_n652), .A2(new_n653), .B1(new_n654), .B2(KEYINPUT8), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n649), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G99gat), .B(G106gat), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n649), .A2(new_n655), .A3(new_n657), .A4(new_n651), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n656), .A2(KEYINPUT101), .A3(new_n658), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n662), .A2(KEYINPUT102), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(KEYINPUT102), .B1(new_n662), .B2(new_n663), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n666), .B1(new_n252), .B2(new_n256), .ZN(new_n667));
  NAND3_X1  g466(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n259), .B1(new_n664), .B2(new_n665), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(G190gat), .B(G218gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(G134gat), .B(G162gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n675));
  AOI21_X1  g474(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n670), .A2(new_n673), .ZN(new_n678));
  AND3_X1   g477(.A1(new_n674), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n677), .B1(new_n678), .B2(new_n674), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n659), .A2(new_n661), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n613), .A2(new_n622), .A3(new_n682), .ZN(new_n683));
  AOI22_X1  g482(.A1(new_n613), .A2(new_n622), .B1(new_n662), .B2(new_n663), .ZN(new_n684));
  NAND2_X1  g483(.A1(G230gat), .A2(G233gat), .ZN(new_n685));
  OR3_X1    g484(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT105), .ZN(new_n687));
  INV_X1    g486(.A(new_n685), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT10), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n689), .B1(new_n683), .B2(new_n684), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n623), .B(KEYINPUT10), .C1(new_n664), .C2(new_n665), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n688), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(G120gat), .B(G148gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT106), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(new_n316), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(new_n449), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n687), .A2(new_n692), .A3(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n686), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n696), .B1(new_n698), .B2(new_n692), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n699), .A2(KEYINPUT107), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(KEYINPUT107), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n697), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n646), .A2(new_n681), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(KEYINPUT108), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n646), .A2(new_n681), .A3(new_n705), .A4(new_n702), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n599), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n438), .A2(new_n440), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(G1gat), .ZN(G1324gat));
  INV_X1    g511(.A(new_n555), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n708), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n212), .A2(new_n225), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(KEYINPUT42), .Z(new_n718));
  NAND2_X1  g517(.A1(new_n714), .A2(G8gat), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n719), .B(KEYINPUT109), .Z(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(G1325gat));
  AOI21_X1  g520(.A(G15gat), .B1(new_n708), .B2(new_n374), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n562), .A2(new_n215), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n722), .B1(new_n708), .B2(new_n723), .ZN(G1326gat));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n536), .ZN(new_n725));
  XNOR2_X1  g524(.A(KEYINPUT43), .B(G22gat), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(G1327gat));
  INV_X1    g526(.A(new_n646), .ZN(new_n728));
  INV_X1    g527(.A(new_n681), .ZN(new_n729));
  AND4_X1   g528(.A1(new_n728), .A2(new_n599), .A3(new_n729), .A4(new_n702), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n730), .A2(new_n237), .A3(new_n710), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT45), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n557), .A2(new_n598), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n729), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT44), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n681), .B1(new_n557), .B2(new_n598), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n291), .A2(new_n292), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n728), .A2(new_n702), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n733), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n737), .A2(new_n738), .ZN(new_n745));
  AOI211_X1 g544(.A(KEYINPUT44), .B(new_n681), .C1(new_n557), .C2(new_n598), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n733), .B(new_n742), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n709), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n732), .B1(new_n748), .B2(new_n237), .ZN(G1328gat));
  NAND3_X1  g548(.A1(new_n730), .A2(new_n238), .A3(new_n713), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n750), .B(KEYINPUT46), .Z(new_n751));
  AOI21_X1  g550(.A(new_n555), .B1(new_n744), .B2(new_n747), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n751), .B1(new_n238), .B2(new_n752), .ZN(G1329gat));
  NAND2_X1  g552(.A1(new_n740), .A2(new_n742), .ZN(new_n754));
  OAI21_X1  g553(.A(G43gat), .B1(new_n754), .B2(new_n562), .ZN(new_n755));
  INV_X1    g554(.A(G43gat), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n730), .A2(new_n756), .A3(new_n374), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n755), .A2(KEYINPUT47), .A3(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n757), .ZN(new_n759));
  INV_X1    g558(.A(new_n562), .ZN(new_n760));
  INV_X1    g559(.A(new_n747), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n743), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n759), .B1(new_n762), .B2(G43gat), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n758), .B1(new_n763), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g563(.A(G50gat), .B1(new_n754), .B2(new_n549), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n549), .A2(G50gat), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT111), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n730), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n765), .A2(KEYINPUT48), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n768), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n536), .B1(new_n743), .B2(new_n761), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n771), .B2(G50gat), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n769), .B1(new_n772), .B2(KEYINPUT48), .ZN(G1331gat));
  AOI211_X1 g572(.A(new_n728), .B(new_n729), .C1(new_n557), .C2(new_n598), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n702), .A2(new_n741), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n776), .A2(new_n709), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(new_n615), .ZN(G1332gat));
  INV_X1    g577(.A(KEYINPUT112), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n555), .B(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n782));
  AND2_X1   g581(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n781), .B2(new_n782), .ZN(G1333gat));
  AND2_X1   g584(.A1(new_n774), .A2(new_n775), .ZN(new_n786));
  AOI21_X1  g585(.A(G71gat), .B1(new_n786), .B2(new_n374), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n776), .A2(new_n352), .A3(new_n562), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XOR2_X1   g588(.A(new_n789), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g589(.A1(new_n786), .A2(new_n536), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g591(.A1(new_n646), .A2(new_n741), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n700), .A2(new_n701), .ZN(new_n794));
  INV_X1    g593(.A(new_n697), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  XOR2_X1   g596(.A(new_n797), .B(KEYINPUT113), .Z(new_n798));
  NAND2_X1  g597(.A1(new_n740), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(G85gat), .B1(new_n799), .B2(new_n709), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n737), .A2(KEYINPUT51), .A3(new_n793), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT51), .B1(new_n737), .B2(new_n793), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n796), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n710), .A2(new_n650), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n800), .B1(new_n803), .B2(new_n804), .ZN(G1336gat));
  OAI21_X1  g604(.A(G92gat), .B1(new_n799), .B2(new_n780), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n780), .A2(G92gat), .A3(new_n702), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(new_n801), .B2(new_n802), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n806), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n740), .A2(new_n713), .A3(new_n798), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n737), .A2(new_n793), .ZN(new_n812));
  NOR2_X1   g611(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n813));
  OR2_X1    g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI22_X1  g615(.A1(G92gat), .A2(new_n811), .B1(new_n816), .B2(new_n808), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n810), .B1(new_n817), .B2(new_n807), .ZN(G1337gat));
  OAI21_X1  g617(.A(G99gat), .B1(new_n799), .B2(new_n562), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n374), .A2(new_n354), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n819), .B1(new_n803), .B2(new_n820), .ZN(G1338gat));
  NAND3_X1  g620(.A1(new_n740), .A2(new_n536), .A3(new_n798), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(G106gat), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n549), .A2(G106gat), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n796), .B(new_n824), .C1(new_n801), .C2(new_n802), .ZN(new_n825));
  XOR2_X1   g624(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n826));
  NAND3_X1  g625(.A1(new_n823), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n702), .B1(new_n814), .B2(new_n815), .ZN(new_n828));
  AOI22_X1  g627(.A1(new_n828), .A2(new_n824), .B1(new_n822), .B2(G106gat), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n827), .B1(new_n829), .B2(new_n830), .ZN(G1339gat));
  NOR2_X1   g630(.A1(new_n703), .A2(new_n741), .ZN(new_n832));
  INV_X1    g631(.A(new_n692), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n690), .A2(new_n691), .A3(new_n688), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n833), .A2(KEYINPUT54), .A3(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n696), .ZN(new_n836));
  XNOR2_X1  g635(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n836), .B1(new_n692), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(KEYINPUT55), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n835), .A2(new_n841), .A3(new_n838), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n697), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n257), .A2(new_n264), .ZN(new_n844));
  OAI22_X1  g643(.A1(new_n280), .A2(new_n278), .B1(new_n844), .B2(new_n265), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n207), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n292), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n729), .A2(new_n843), .A3(new_n847), .ZN(new_n848));
  AOI22_X1  g647(.A1(new_n741), .A2(new_n843), .B1(new_n796), .B2(new_n847), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n848), .B1(new_n849), .B2(new_n729), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n832), .B1(new_n850), .B2(new_n728), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n851), .A2(new_n709), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n549), .A2(new_n374), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n852), .A2(new_n853), .A3(new_n780), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(G113gat), .B1(new_n855), .B2(new_n294), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n854), .A2(new_n332), .A3(new_n741), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1340gat));
  NAND2_X1  g657(.A1(new_n854), .A2(new_n796), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g659(.A1(new_n854), .A2(new_n646), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n861), .B(G127gat), .ZN(G1342gat));
  OAI21_X1  g661(.A(G134gat), .B1(new_n855), .B2(new_n681), .ZN(new_n863));
  NOR4_X1   g662(.A1(new_n851), .A2(new_n709), .A3(new_n681), .A4(new_n713), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(new_n326), .A3(new_n853), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n865), .A2(KEYINPUT56), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(KEYINPUT56), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n863), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n868), .B(new_n869), .ZN(G1343gat));
  NAND2_X1  g669(.A1(new_n843), .A2(new_n741), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n796), .A2(new_n847), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n729), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n848), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n728), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n832), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n536), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n780), .A2(new_n710), .A3(new_n562), .ZN(new_n879));
  NOR4_X1   g678(.A1(new_n878), .A2(G141gat), .A3(new_n294), .A4(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n285), .A2(new_n843), .A3(new_n293), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n729), .B1(new_n881), .B2(new_n872), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n728), .B1(new_n882), .B2(new_n874), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n876), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n536), .A2(KEYINPUT57), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XOR2_X1   g688(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n878), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n885), .B1(new_n883), .B2(new_n876), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT119), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n889), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n879), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n741), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n880), .B1(new_n898), .B2(G141gat), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT58), .ZN(new_n900));
  INV_X1    g699(.A(new_n294), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n386), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n880), .A2(KEYINPUT58), .ZN(new_n903));
  OAI22_X1  g702(.A1(new_n899), .A2(new_n900), .B1(new_n902), .B2(new_n903), .ZN(G1344gat));
  NAND3_X1  g703(.A1(new_n895), .A2(new_n796), .A3(new_n896), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n384), .A2(KEYINPUT59), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT120), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n879), .B(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n707), .A2(new_n294), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n883), .ZN(new_n910));
  AOI21_X1  g709(.A(KEYINPUT57), .B1(new_n910), .B2(new_n536), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n851), .A2(new_n549), .A3(new_n891), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n796), .B(new_n908), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(G148gat), .ZN(new_n914));
  AOI22_X1  g713(.A1(new_n905), .A2(new_n906), .B1(new_n914), .B2(KEYINPUT59), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n878), .A2(new_n879), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n384), .A3(new_n796), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(KEYINPUT121), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n905), .A2(new_n906), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT59), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n922), .B1(new_n913), .B2(G148gat), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n920), .B(new_n917), .C1(new_n921), .C2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n919), .A2(new_n924), .ZN(G1345gat));
  NAND3_X1  g724(.A1(new_n916), .A2(new_n381), .A3(new_n646), .ZN(new_n926));
  INV_X1    g725(.A(new_n897), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n927), .A2(new_n728), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n926), .B1(new_n928), .B2(new_n381), .ZN(G1346gat));
  OAI21_X1  g728(.A(G162gat), .B1(new_n927), .B2(new_n681), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n760), .A2(new_n549), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n864), .A2(new_n382), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(G1347gat));
  NAND2_X1  g732(.A1(new_n713), .A2(new_n709), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT122), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n877), .A2(new_n853), .A3(new_n935), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n936), .A2(new_n315), .A3(new_n294), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n851), .A2(new_n710), .ZN(new_n938));
  INV_X1    g737(.A(new_n780), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n938), .A2(new_n853), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(new_n741), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n937), .B1(new_n941), .B2(new_n315), .ZN(new_n942));
  XOR2_X1   g741(.A(new_n942), .B(KEYINPUT123), .Z(G1348gat));
  NOR3_X1   g742(.A1(new_n936), .A2(new_n316), .A3(new_n702), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT124), .ZN(new_n945));
  AOI21_X1  g744(.A(G176gat), .B1(new_n940), .B2(new_n796), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n945), .A2(new_n946), .ZN(G1349gat));
  OAI211_X1 g746(.A(new_n940), .B(new_n646), .C1(new_n298), .C2(new_n297), .ZN(new_n948));
  OAI21_X1  g747(.A(G183gat), .B1(new_n936), .B2(new_n728), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n948), .A2(KEYINPUT125), .A3(new_n949), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g750(.A(G190gat), .B1(new_n936), .B2(new_n681), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT61), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n940), .A2(new_n296), .A3(new_n729), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1351gat));
  AOI21_X1  g754(.A(new_n549), .B1(new_n909), .B2(new_n883), .ZN(new_n956));
  OAI22_X1  g755(.A1(new_n878), .A2(new_n891), .B1(new_n956), .B2(KEYINPUT57), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n935), .A2(new_n562), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(G197gat), .B1(new_n959), .B2(new_n294), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n938), .A2(new_n939), .A3(new_n931), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n961), .A2(new_n448), .A3(new_n741), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(G1352gat));
  NAND2_X1  g762(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n961), .A2(new_n449), .A3(new_n796), .A4(new_n964), .ZN(new_n965));
  NOR2_X1   g764(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n965), .B(new_n966), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n957), .A2(new_n796), .A3(new_n958), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n967), .B1(new_n449), .B2(new_n968), .ZN(G1353gat));
  INV_X1    g768(.A(new_n446), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n961), .A2(new_n646), .A3(new_n970), .ZN(new_n971));
  OAI211_X1 g770(.A(new_n646), .B(new_n958), .C1(new_n911), .C2(new_n912), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(KEYINPUT127), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT127), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n957), .A2(new_n974), .A3(new_n646), .A4(new_n958), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n973), .A2(G211gat), .A3(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT63), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n976), .A2(new_n977), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n971), .B1(new_n978), .B2(new_n979), .ZN(G1354gat));
  NOR3_X1   g779(.A1(new_n959), .A2(new_n442), .A3(new_n681), .ZN(new_n981));
  AOI21_X1  g780(.A(G218gat), .B1(new_n961), .B2(new_n729), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n981), .A2(new_n982), .ZN(G1355gat));
endmodule


