//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  NAND2_X1  g000(.A1(G234), .A2(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND3_X1   g002(.A1(new_n187), .A2(G952), .A3(new_n188), .ZN(new_n189));
  AND3_X1   g003(.A1(new_n187), .A2(G902), .A3(G953), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT21), .B(G898), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n189), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  OAI21_X1  g006(.A(G214), .B1(G237), .B2(G902), .ZN(new_n193));
  XOR2_X1   g007(.A(new_n193), .B(KEYINPUT83), .Z(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(G210), .B1(G237), .B2(G902), .ZN(new_n196));
  INV_X1    g010(.A(G116), .ZN(new_n197));
  INV_X1    g011(.A(G119), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(G116), .A2(G119), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  OR2_X1    g015(.A1(KEYINPUT2), .A2(G113), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT2), .A2(G113), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(KEYINPUT67), .A3(new_n203), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT2), .A2(G113), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT2), .A2(G113), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n201), .B1(new_n205), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT68), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n204), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI211_X1 g026(.A(KEYINPUT68), .B(new_n201), .C1(new_n209), .C2(new_n205), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT69), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n205), .A2(new_n209), .ZN(new_n215));
  INV_X1    g029(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT68), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT69), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n210), .A2(new_n211), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n204), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n214), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT77), .ZN(new_n223));
  INV_X1    g037(.A(G107), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n224), .A3(G104), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT3), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n223), .A2(new_n227), .A3(new_n224), .A4(G104), .ZN(new_n228));
  INV_X1    g042(.A(G104), .ZN(new_n229));
  AOI21_X1  g043(.A(G101), .B1(new_n229), .B2(G107), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n226), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT78), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n226), .A2(KEYINPUT78), .A3(new_n228), .A4(new_n230), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT4), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n229), .A2(G107), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n226), .A2(new_n228), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n236), .B1(new_n238), .B2(G101), .ZN(new_n239));
  OAI21_X1  g053(.A(G101), .B1(new_n236), .B2(KEYINPUT79), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n240), .B1(KEYINPUT79), .B2(new_n236), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT80), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT80), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n238), .A2(new_n244), .A3(new_n241), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n235), .A2(new_n239), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n222), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT5), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(new_n198), .A3(G116), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G113), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n250), .B1(KEYINPUT5), .B2(new_n201), .ZN(new_n251));
  INV_X1    g065(.A(new_n204), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n224), .A2(G104), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(new_n237), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G101), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n235), .A2(new_n253), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n247), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(G110), .B(G122), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(KEYINPUT84), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n259), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n263), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n257), .B1(new_n222), .B2(new_n246), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n265), .B1(new_n266), .B2(new_n260), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n260), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n264), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(G143), .B(G146), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT0), .ZN(new_n271));
  INV_X1    g085(.A(G128), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  XOR2_X1   g087(.A(KEYINPUT0), .B(G128), .Z(new_n274));
  OAI21_X1  g088(.A(new_n273), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G125), .ZN(new_n276));
  OAI21_X1  g090(.A(KEYINPUT85), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  OR2_X1    g091(.A1(new_n274), .A2(new_n270), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT85), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n278), .A2(new_n273), .A3(new_n279), .A4(G125), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n272), .A2(KEYINPUT1), .ZN(new_n282));
  INV_X1    g096(.A(G143), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G146), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n272), .A2(G143), .ZN(new_n285));
  OAI22_X1  g099(.A1(new_n282), .A2(new_n284), .B1(new_n285), .B2(G146), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT65), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n288), .B1(new_n270), .B2(new_n282), .ZN(new_n289));
  INV_X1    g103(.A(G146), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G143), .ZN(new_n291));
  AND4_X1   g105(.A1(new_n288), .A2(new_n282), .A3(new_n284), .A4(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n287), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n293), .A2(G125), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n281), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n188), .A2(G224), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n295), .B(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n269), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G902), .ZN(new_n301));
  AOI211_X1 g115(.A(new_n261), .B(new_n257), .C1(new_n222), .C2(new_n246), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n260), .B(KEYINPUT8), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n253), .B1(new_n235), .B2(new_n256), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n303), .B1(new_n257), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT7), .ZN(new_n306));
  OAI22_X1  g120(.A1(new_n281), .A2(new_n294), .B1(new_n306), .B2(new_n297), .ZN(new_n307));
  INV_X1    g121(.A(new_n294), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n297), .A2(new_n306), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n308), .A2(new_n277), .A3(new_n280), .A4(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n305), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n301), .B1(new_n302), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n196), .B1(new_n300), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n196), .ZN(new_n315));
  AOI211_X1 g129(.A(new_n315), .B(new_n312), .C1(new_n269), .C2(new_n299), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n195), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n192), .B1(new_n317), .B2(KEYINPUT86), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n259), .A2(new_n261), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n319), .B1(new_n265), .B2(new_n302), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n298), .B1(new_n320), .B2(new_n264), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n315), .B1(new_n321), .B2(new_n312), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n300), .A2(new_n196), .A3(new_n313), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT86), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n325), .A3(new_n195), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n318), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT16), .ZN(new_n328));
  INV_X1    g142(.A(G140), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n329), .A3(G125), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(G125), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n276), .A2(G140), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n330), .B1(new_n333), .B2(new_n328), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n290), .ZN(new_n335));
  NOR2_X1   g149(.A1(G237), .A2(G953), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(G143), .A3(G214), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(G143), .B1(new_n336), .B2(G214), .ZN(new_n339));
  OAI211_X1 g153(.A(KEYINPUT17), .B(G131), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  OAI211_X1 g154(.A(G146), .B(new_n330), .C1(new_n333), .C2(new_n328), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n335), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT90), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G237), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(new_n188), .A3(G214), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n283), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n337), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G131), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT17), .ZN(new_n350));
  INV_X1    g164(.A(G131), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n347), .A2(new_n351), .A3(new_n337), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n349), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n335), .A2(new_n340), .A3(KEYINPUT90), .A4(new_n341), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n344), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT88), .ZN(new_n356));
  INV_X1    g170(.A(G122), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G113), .ZN(new_n358));
  INV_X1    g172(.A(G113), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G122), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n356), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n358), .A2(new_n360), .A3(new_n356), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n363), .A3(G104), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(G104), .B1(new_n362), .B2(new_n363), .ZN(new_n366));
  OAI21_X1  g180(.A(KEYINPUT89), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n366), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT89), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n364), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n348), .A2(KEYINPUT18), .A3(G131), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n333), .A2(G146), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n331), .A2(new_n332), .A3(new_n290), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(KEYINPUT18), .A2(G131), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n347), .A2(new_n337), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n372), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n355), .A2(new_n371), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n365), .A2(new_n366), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n382), .B1(new_n355), .B2(new_n378), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n301), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT91), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT91), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n386), .B(new_n301), .C1(new_n380), .C2(new_n383), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(G475), .A3(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n333), .B(KEYINPUT19), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n341), .B1(new_n389), .B2(G146), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n349), .A2(new_n352), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT87), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n349), .A2(KEYINPUT87), .A3(new_n352), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n390), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n378), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n381), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n379), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G475), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n301), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT20), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT20), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n398), .A2(new_n403), .A3(new_n400), .A4(new_n301), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n388), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(G128), .B(G143), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT13), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n283), .A2(G128), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n408), .B(G134), .C1(KEYINPUT13), .C2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(G116), .B(G122), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(new_n224), .ZN(new_n412));
  INV_X1    g226(.A(G134), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n407), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n410), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n407), .B(new_n413), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n197), .A2(KEYINPUT14), .A3(G122), .ZN(new_n417));
  INV_X1    g231(.A(new_n411), .ZN(new_n418));
  OAI211_X1 g232(.A(G107), .B(new_n417), .C1(new_n418), .C2(KEYINPUT14), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n411), .A2(new_n224), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n416), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n415), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT9), .B(G234), .ZN(new_n423));
  INV_X1    g237(.A(G217), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n423), .A2(new_n424), .A3(G953), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n422), .B(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G478), .ZN(new_n428));
  OR2_X1    g242(.A1(new_n428), .A2(KEYINPUT15), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n427), .A2(new_n301), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n429), .B1(new_n427), .B2(new_n301), .ZN(new_n432));
  OR2_X1    g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n406), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(G221), .B1(new_n423), .B2(G902), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(KEYINPUT75), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G469), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n188), .A2(G227), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(G140), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT76), .B(G110), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n441), .B(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT12), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n235), .A2(new_n256), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n282), .A2(new_n284), .A3(new_n291), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT65), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n270), .A2(new_n288), .A3(new_n282), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n286), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n256), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n447), .A2(new_n448), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n450), .B1(new_n451), .B2(new_n287), .ZN(new_n452));
  AOI22_X1  g266(.A1(new_n445), .A2(new_n449), .B1(new_n235), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT11), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n454), .B1(new_n413), .B2(G137), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n413), .A2(G137), .ZN(new_n456));
  INV_X1    g270(.A(G137), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(KEYINPUT11), .A3(G134), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n455), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n351), .A2(KEYINPUT64), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n459), .B(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n444), .B1(new_n453), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n235), .A2(new_n293), .A3(new_n256), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n293), .B1(new_n235), .B2(new_n256), .ZN(new_n466));
  OAI211_X1 g280(.A(KEYINPUT12), .B(new_n461), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n235), .A2(new_n239), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n243), .A2(new_n245), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n469), .A3(new_n275), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT10), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n464), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n452), .A2(KEYINPUT10), .A3(new_n235), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n470), .A2(new_n472), .A3(new_n462), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT81), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n452), .A2(KEYINPUT10), .A3(new_n235), .ZN(new_n476));
  AOI21_X1  g290(.A(KEYINPUT10), .B1(new_n452), .B2(new_n235), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT81), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n478), .A2(new_n479), .A3(new_n462), .A4(new_n470), .ZN(new_n480));
  AOI221_X4 g294(.A(new_n443), .B1(new_n463), .B2(new_n467), .C1(new_n475), .C2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n443), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n475), .A2(new_n480), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n478), .A2(new_n470), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n461), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n482), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n439), .B(new_n301), .C1(new_n481), .C2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n483), .A2(new_n485), .A3(new_n482), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n475), .A2(new_n480), .B1(new_n467), .B2(new_n463), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n489), .B(G469), .C1(new_n482), .C2(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n439), .A2(new_n301), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n438), .B1(new_n488), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT82), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT82), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n497), .B(new_n438), .C1(new_n488), .C2(new_n494), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n435), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n327), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n457), .A2(G134), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n351), .B1(new_n413), .B2(G137), .ZN(new_n502));
  AOI22_X1  g316(.A1(new_n459), .A2(new_n351), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT66), .B1(new_n449), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n501), .ZN(new_n505));
  INV_X1    g319(.A(new_n459), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n505), .B1(new_n506), .B2(G131), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT66), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n293), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n461), .A2(new_n275), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n504), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n222), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n507), .A2(KEYINPUT70), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT70), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n503), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n513), .A2(new_n293), .A3(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n516), .A2(new_n214), .A3(new_n221), .A4(new_n510), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT28), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT28), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n336), .A2(G210), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n522), .B(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT26), .B(G101), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n524), .B(new_n525), .ZN(new_n526));
  AND4_X1   g340(.A1(new_n512), .A2(new_n519), .A3(new_n521), .A4(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT30), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n511), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n516), .A2(KEYINPUT30), .A3(new_n510), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n222), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n526), .B1(new_n531), .B2(new_n517), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n527), .A2(KEYINPUT29), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n516), .A2(new_n510), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n222), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n519), .A2(new_n521), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n526), .A2(KEYINPUT29), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n301), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(G472), .B1(new_n533), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT32), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n531), .A2(new_n517), .A3(new_n526), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT31), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n531), .A2(KEYINPUT31), .A3(new_n517), .A4(new_n526), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n519), .A2(new_n512), .A3(new_n521), .ZN(new_n545));
  INV_X1    g359(.A(new_n526), .ZN(new_n546));
  AOI22_X1  g360(.A1(new_n543), .A2(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(G472), .A2(G902), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n540), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n543), .A2(new_n544), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n545), .A2(new_n546), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(KEYINPUT32), .A3(new_n548), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n539), .A2(new_n550), .A3(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(G119), .B(G128), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(KEYINPUT72), .ZN(new_n557));
  XOR2_X1   g371(.A(KEYINPUT24), .B(G110), .Z(new_n558));
  OAI211_X1 g372(.A(new_n272), .B(G119), .C1(KEYINPUT73), .C2(KEYINPUT23), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT23), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n560), .B1(new_n198), .B2(G128), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT73), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n562), .B1(new_n198), .B2(G128), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n559), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n557), .A2(new_n558), .B1(G110), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n335), .A2(new_n341), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI22_X1  g381(.A1(new_n557), .A2(new_n558), .B1(G110), .B2(new_n564), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n341), .A2(new_n374), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT74), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n570), .B1(new_n568), .B2(new_n569), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n567), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(KEYINPUT22), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(G137), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n567), .B(new_n576), .C1(new_n571), .C2(new_n572), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n424), .B1(G234), .B2(new_n301), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(G902), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n578), .A2(new_n301), .A3(new_n579), .ZN(new_n585));
  OR2_X1    g399(.A1(new_n585), .A2(KEYINPUT25), .ZN(new_n586));
  INV_X1    g400(.A(new_n581), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n587), .B1(new_n585), .B2(KEYINPUT25), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n584), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n555), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n500), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(G101), .ZN(G3));
  INV_X1    g407(.A(KEYINPUT93), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT33), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(KEYINPUT93), .A2(KEYINPUT33), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n427), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n426), .A2(new_n594), .A3(new_n595), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(G478), .A3(new_n301), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n428), .B1(new_n426), .B2(G902), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n406), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n317), .A2(KEYINPUT92), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT92), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n606), .B(new_n195), .C1(new_n314), .C2(new_n316), .ZN(new_n607));
  AOI211_X1 g421(.A(new_n192), .B(new_n604), .C1(new_n605), .C2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(G472), .B1(new_n547), .B2(G902), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n553), .A2(new_n548), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(new_n610), .A3(new_n589), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n611), .B1(new_n496), .B2(new_n498), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(new_n613), .B(KEYINPUT94), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT95), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT34), .B(G104), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G6));
  INV_X1    g431(.A(new_n406), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n433), .ZN(new_n619));
  AOI211_X1 g433(.A(new_n192), .B(new_n619), .C1(new_n605), .C2(new_n607), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n612), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT35), .B(G107), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT96), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n621), .B(new_n623), .ZN(G9));
  NOR2_X1   g438(.A1(new_n577), .A2(KEYINPUT36), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n573), .B(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n586), .A2(new_n588), .B1(new_n582), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(KEYINPUT97), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT97), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  AND4_X1   g447(.A1(new_n610), .A2(new_n631), .A3(new_n609), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n500), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT37), .B(G110), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G12));
  NAND2_X1  g451(.A1(new_n496), .A2(new_n498), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n555), .A2(new_n631), .A3(new_n633), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n605), .A2(new_n607), .ZN(new_n640));
  INV_X1    g454(.A(G900), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n189), .B1(new_n190), .B2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n433), .A2(new_n388), .A3(new_n405), .A4(new_n643), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n644), .A2(KEYINPUT98), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(KEYINPUT98), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n638), .A2(new_n639), .A3(new_n640), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G128), .ZN(G30));
  XOR2_X1   g463(.A(new_n642), .B(KEYINPUT39), .Z(new_n650));
  NAND2_X1  g464(.A1(new_n638), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(new_n651), .B(KEYINPUT40), .Z(new_n652));
  AND2_X1   g466(.A1(new_n324), .A2(KEYINPUT99), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n324), .A2(KEYINPUT99), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT38), .ZN(new_n655));
  OR3_X1    g469(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n655), .B1(new_n653), .B2(new_n654), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n554), .A2(new_n550), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n531), .A2(new_n517), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n526), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n518), .A2(new_n526), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n535), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n662), .A2(new_n301), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(G472), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n660), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n668), .A2(new_n630), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n431), .A2(new_n432), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n388), .B2(new_n405), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n671), .A2(new_n195), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n652), .A2(new_n659), .A3(new_n669), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G143), .ZN(G45));
  NOR2_X1   g488(.A1(new_n604), .A2(new_n642), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n638), .A2(new_n639), .A3(new_n640), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G146), .ZN(G48));
  NAND2_X1  g491(.A1(new_n483), .A2(new_n485), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n443), .B1(new_n475), .B2(new_n480), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n463), .A2(new_n467), .ZN(new_n680));
  AOI22_X1  g494(.A1(new_n678), .A2(new_n443), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(G469), .B1(new_n681), .B2(G902), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n682), .A2(new_n436), .A3(new_n487), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT100), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT101), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n682), .A2(KEYINPUT100), .A3(new_n436), .A4(new_n487), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n686), .B1(new_n685), .B2(new_n687), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n688), .A2(new_n689), .A3(new_n590), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n690), .A2(KEYINPUT102), .A3(new_n608), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n685), .A2(new_n687), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(KEYINPUT101), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n608), .A2(new_n693), .A3(new_n591), .A4(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT102), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n691), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT41), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G113), .ZN(G15));
  AND4_X1   g514(.A1(new_n591), .A2(new_n620), .A3(new_n693), .A4(new_n694), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n197), .ZN(G18));
  INV_X1    g516(.A(new_n192), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n639), .A2(new_n703), .A3(new_n434), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n606), .B1(new_n324), .B2(new_n195), .ZN(new_n705));
  INV_X1    g519(.A(new_n607), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(KEYINPUT103), .B1(new_n707), .B2(new_n692), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT103), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n640), .A2(new_n709), .A3(new_n685), .A4(new_n687), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n704), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(new_n198), .ZN(G21));
  XOR2_X1   g526(.A(KEYINPUT105), .B(G472), .Z(new_n713));
  OAI21_X1  g527(.A(new_n713), .B1(new_n547), .B2(G902), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n536), .A2(new_n546), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n551), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g530(.A(new_n548), .B(KEYINPUT104), .Z(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n714), .A2(new_n671), .A3(new_n718), .A4(new_n589), .ZN(new_n719));
  AOI211_X1 g533(.A(new_n192), .B(new_n719), .C1(new_n605), .C2(new_n607), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n693), .A3(new_n694), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G122), .ZN(G24));
  AND2_X1   g536(.A1(new_n714), .A2(new_n718), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n630), .ZN(new_n724));
  INV_X1    g538(.A(new_n675), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n727), .B1(new_n708), .B2(new_n710), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(new_n276), .ZN(G27));
  NAND3_X1  g543(.A1(new_n322), .A2(new_n195), .A3(new_n323), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n590), .A2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n436), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n483), .A2(new_n680), .ZN(new_n733));
  AOI22_X1  g547(.A1(new_n733), .A2(new_n443), .B1(new_n679), .B2(new_n485), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n492), .B1(new_n734), .B2(G469), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n732), .B1(new_n735), .B2(new_n487), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n731), .A2(KEYINPUT42), .A3(new_n675), .A4(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT42), .ZN(new_n738));
  INV_X1    g552(.A(new_n730), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n739), .A2(new_n736), .A3(new_n555), .A4(new_n589), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n738), .B1(new_n740), .B2(new_n725), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G131), .ZN(G33));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n647), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n645), .A2(new_n646), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT106), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n745), .A2(new_n731), .A3(new_n736), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G134), .ZN(G36));
  INV_X1    g563(.A(KEYINPUT46), .ZN(new_n750));
  OAI21_X1  g564(.A(G469), .B1(new_n734), .B2(KEYINPUT45), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(KEYINPUT107), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT107), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n753), .B(G469), .C1(new_n734), .C2(KEYINPUT45), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n734), .A2(KEYINPUT45), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n752), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(KEYINPUT108), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT108), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n752), .A2(new_n754), .A3(new_n758), .A4(new_n755), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n750), .B1(new_n760), .B2(new_n492), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n492), .B1(new_n757), .B2(new_n759), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT46), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n761), .A2(new_n487), .A3(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT109), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT43), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n765), .A2(KEYINPUT43), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  AOI22_X1  g582(.A1(new_n618), .A2(new_n603), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n601), .A2(new_n602), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n770), .A2(new_n406), .A3(new_n767), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n609), .A2(new_n610), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n773), .A3(new_n630), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n772), .A2(KEYINPUT44), .A3(new_n773), .A4(new_n630), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n776), .A2(new_n739), .A3(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n764), .A2(new_n778), .A3(new_n436), .A4(new_n650), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT110), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(new_n457), .ZN(G39));
  OAI21_X1  g595(.A(new_n487), .B1(new_n762), .B2(KEYINPUT46), .ZN(new_n782));
  AOI211_X1 g596(.A(new_n750), .B(new_n492), .C1(new_n757), .C2(new_n759), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n436), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT47), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT47), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n786), .B(new_n436), .C1(new_n782), .C2(new_n783), .ZN(new_n787));
  NOR4_X1   g601(.A1(new_n725), .A2(new_n555), .A3(new_n589), .A4(new_n730), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n785), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT111), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n785), .A2(KEYINPUT111), .A3(new_n787), .A4(new_n788), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G140), .ZN(G42));
  NOR2_X1   g608(.A1(G952), .A2(G953), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n648), .A2(new_n676), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n728), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n640), .A2(new_n671), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n667), .A2(new_n629), .A3(new_n643), .A4(new_n736), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(new_n799), .B2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n728), .A2(new_n798), .A3(new_n805), .A4(new_n802), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n327), .B(new_n499), .C1(new_n591), .C2(new_n634), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n619), .A2(new_n604), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n327), .A2(new_n612), .A3(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n808), .A2(new_n721), .A3(new_n810), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n811), .A2(new_n701), .A3(new_n711), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n737), .A2(new_n741), .ZN(new_n813));
  INV_X1    g627(.A(new_n604), .ZN(new_n814));
  AND4_X1   g628(.A1(new_n814), .A2(new_n736), .A3(new_n630), .A4(new_n723), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n815), .B1(new_n499), .B2(new_n639), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n739), .A2(new_n643), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n748), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n813), .B1(new_n818), .B2(KEYINPUT113), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT113), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n748), .B(new_n820), .C1(new_n816), .C2(new_n817), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n812), .A2(new_n819), .A3(new_n698), .A4(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n797), .B1(new_n807), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n708), .A2(new_n710), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n726), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n648), .A2(new_n676), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n825), .A2(new_n826), .A3(new_n803), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n805), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n799), .A2(KEYINPUT52), .A3(new_n803), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n818), .A2(KEYINPUT113), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n831), .A2(new_n742), .A3(new_n821), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n701), .A2(new_n711), .ZN(new_n833));
  INV_X1    g647(.A(new_n811), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n698), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n830), .A2(KEYINPUT53), .A3(new_n832), .A4(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n796), .B1(new_n823), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT114), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n823), .A2(new_n838), .A3(new_n836), .ZN(new_n839));
  OAI211_X1 g653(.A(KEYINPUT114), .B(new_n797), .C1(new_n807), .C2(new_n822), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n837), .B1(new_n841), .B2(new_n796), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n685), .A2(new_n687), .A3(new_n739), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT116), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n843), .B(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n189), .B1(new_n769), .B2(new_n771), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT115), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI211_X1 g662(.A(KEYINPUT115), .B(new_n189), .C1(new_n769), .C2(new_n771), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n845), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(new_n630), .A3(new_n723), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n723), .A2(new_n589), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n853), .B1(new_n848), .B2(new_n849), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n692), .A2(new_n195), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n854), .A2(new_n658), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT50), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n854), .A2(new_n658), .A3(KEYINPUT50), .A4(new_n855), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n668), .A2(new_n589), .A3(new_n189), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n845), .A2(new_n618), .A3(new_n770), .A4(new_n861), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n852), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n682), .A2(new_n487), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n438), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n865), .B1(new_n785), .B2(new_n787), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n739), .B(new_n854), .C1(new_n866), .C2(KEYINPUT117), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n866), .A2(KEYINPUT117), .ZN(new_n868));
  OAI211_X1 g682(.A(KEYINPUT51), .B(new_n863), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n845), .A2(new_n814), .A3(new_n861), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n188), .A2(G952), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(new_n824), .B2(new_n854), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT48), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n851), .A2(new_n873), .A3(new_n591), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n873), .B1(new_n851), .B2(new_n591), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n870), .B(new_n872), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n854), .A2(new_n739), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n863), .B1(new_n866), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT51), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n876), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n869), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n795), .B1(new_n842), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n437), .A2(new_n194), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n618), .A2(new_n589), .A3(new_n603), .A4(new_n884), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n885), .A2(KEYINPUT112), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n885), .A2(KEYINPUT112), .B1(new_n864), .B2(KEYINPUT49), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n864), .A2(KEYINPUT49), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n668), .A2(new_n886), .A3(new_n887), .A4(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n659), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(KEYINPUT118), .B1(new_n883), .B2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT118), .ZN(new_n892));
  INV_X1    g706(.A(new_n890), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT54), .B1(new_n839), .B2(new_n840), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n881), .A2(new_n894), .A3(new_n837), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n892), .B(new_n893), .C1(new_n895), .C2(new_n795), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n891), .A2(new_n896), .ZN(G75));
  NAND4_X1  g711(.A1(new_n839), .A2(G210), .A3(G902), .A4(new_n840), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n269), .B(new_n299), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT55), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(KEYINPUT56), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n188), .A2(G952), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n898), .A2(KEYINPUT119), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT56), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n898), .A2(KEYINPUT119), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n905), .B1(new_n909), .B2(new_n900), .ZN(G51));
  XNOR2_X1  g724(.A(new_n492), .B(KEYINPUT57), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n841), .A2(new_n796), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n911), .B1(new_n912), .B2(new_n894), .ZN(new_n913));
  INV_X1    g727(.A(new_n681), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n841), .A2(new_n301), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n760), .B(KEYINPUT120), .Z(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n903), .B1(new_n915), .B2(new_n918), .ZN(G54));
  AND2_X1   g733(.A1(KEYINPUT58), .A2(G475), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n916), .A2(new_n398), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n398), .B1(new_n916), .B2(new_n920), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n921), .A2(new_n922), .A3(new_n903), .ZN(G60));
  XOR2_X1   g737(.A(new_n600), .B(KEYINPUT121), .Z(new_n924));
  NAND2_X1  g738(.A1(G478), .A2(G902), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT59), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n924), .B(new_n926), .C1(new_n912), .C2(new_n894), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n904), .ZN(new_n928));
  INV_X1    g742(.A(new_n842), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n924), .B1(new_n929), .B2(new_n926), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n928), .A2(new_n930), .ZN(G63));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n932), .A2(KEYINPUT122), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(KEYINPUT122), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT123), .Z(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(G217), .A2(G902), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT60), .Z(new_n938));
  NAND3_X1  g752(.A1(new_n839), .A2(new_n840), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n903), .B1(new_n939), .B2(new_n580), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n839), .A2(new_n628), .A3(new_n840), .A4(new_n938), .ZN(new_n941));
  AOI211_X1 g755(.A(new_n933), .B(new_n936), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n939), .A2(new_n580), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n943), .A2(new_n904), .A3(new_n941), .ZN(new_n944));
  INV_X1    g758(.A(new_n933), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n935), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n942), .A2(new_n946), .ZN(G66));
  NAND2_X1  g761(.A1(G224), .A2(G953), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n191), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n949), .B1(new_n835), .B2(new_n188), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT124), .Z(new_n951));
  OAI211_X1 g765(.A(new_n320), .B(new_n264), .C1(G898), .C2(new_n188), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(G69));
  NAND2_X1  g767(.A1(new_n641), .A2(G953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n800), .A2(new_n590), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n764), .A2(new_n436), .A3(new_n650), .A4(new_n955), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n742), .A2(new_n748), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n779), .A2(new_n956), .A3(new_n799), .A4(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n958), .B1(new_n791), .B2(new_n792), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n954), .B1(new_n959), .B2(G953), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(KEYINPUT126), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n962), .B(new_n954), .C1(new_n959), .C2(G953), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(G227), .A2(G900), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n529), .A2(new_n530), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(new_n389), .ZN(new_n967));
  AND4_X1   g781(.A1(G953), .A2(new_n964), .A3(new_n965), .A4(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n967), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n961), .B2(new_n963), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n673), .A2(new_n799), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT62), .ZN(new_n972));
  INV_X1    g786(.A(new_n793), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n731), .A2(new_n638), .A3(new_n650), .A4(new_n809), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n779), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT125), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n972), .A2(new_n973), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n969), .A2(new_n188), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n980));
  NOR3_X1   g794(.A1(new_n970), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n968), .A2(new_n981), .ZN(G72));
  NAND2_X1  g796(.A1(new_n977), .A2(new_n835), .ZN(new_n983));
  NAND2_X1  g797(.A1(G472), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT63), .Z(new_n985));
  AOI21_X1  g799(.A(new_n662), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n823), .A2(new_n836), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT127), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n541), .A2(new_n988), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(new_n532), .Z(new_n990));
  NAND3_X1  g804(.A1(new_n987), .A2(new_n985), .A3(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n985), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n992), .B1(new_n959), .B2(new_n835), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n663), .A2(new_n531), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n991), .B(new_n904), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n986), .A2(new_n995), .ZN(G57));
endmodule


