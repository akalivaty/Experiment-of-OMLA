

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U552 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X2 U553 ( .A1(n520), .A2(G2104), .ZN(n886) );
  AND2_X2 U554 ( .A1(G2105), .A2(G2104), .ZN(n893) );
  AND2_X2 U555 ( .A1(G160), .A2(G40), .ZN(n689) );
  XNOR2_X1 U556 ( .A(n691), .B(n690), .ZN(n694) );
  NAND2_X1 U557 ( .A1(n722), .A2(G2072), .ZN(n691) );
  INV_X1 U558 ( .A(KEYINPUT27), .ZN(n690) );
  INV_X1 U559 ( .A(KEYINPUT28), .ZN(n696) );
  NOR2_X1 U560 ( .A1(n979), .A2(n712), .ZN(n697) );
  NOR2_X2 U561 ( .A1(G2105), .A2(G2104), .ZN(n519) );
  NOR2_X4 U562 ( .A1(G164), .A2(G1384), .ZN(n767) );
  NAND2_X4 U563 ( .A1(n689), .A2(n767), .ZN(n736) );
  INV_X1 U564 ( .A(KEYINPUT29), .ZN(n717) );
  XNOR2_X1 U565 ( .A(n718), .B(n717), .ZN(n726) );
  INV_X1 U566 ( .A(KEYINPUT13), .ZN(n599) );
  XNOR2_X1 U567 ( .A(n599), .B(KEYINPUT70), .ZN(n600) );
  XNOR2_X1 U568 ( .A(n601), .B(n600), .ZN(n602) );
  NAND2_X1 U569 ( .A1(G114), .A2(n893), .ZN(n521) );
  INV_X1 U570 ( .A(KEYINPUT102), .ZN(n820) );
  NAND2_X1 U571 ( .A1(n819), .A2(n818), .ZN(n821) );
  NOR2_X1 U572 ( .A1(G651), .A2(G543), .ZN(n658) );
  XOR2_X2 U573 ( .A(KEYINPUT17), .B(n519), .Z(n884) );
  NAND2_X1 U574 ( .A1(G138), .A2(n884), .ZN(n527) );
  INV_X1 U575 ( .A(G2105), .ZN(n520) );
  NOR2_X1 U576 ( .A1(G2104), .A2(n520), .ZN(n528) );
  BUF_X1 U577 ( .A(n528), .Z(n890) );
  AND2_X1 U578 ( .A1(G126), .A2(n890), .ZN(n525) );
  NAND2_X1 U579 ( .A1(n886), .A2(G102), .ZN(n523) );
  XOR2_X1 U580 ( .A(KEYINPUT85), .B(n521), .Z(n522) );
  NAND2_X1 U581 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U582 ( .A1(n525), .A2(n524), .ZN(n526) );
  AND2_X2 U583 ( .A1(n527), .A2(n526), .ZN(G164) );
  NAND2_X1 U584 ( .A1(G125), .A2(n528), .ZN(n529) );
  XNOR2_X1 U585 ( .A(n529), .B(KEYINPUT64), .ZN(n532) );
  NAND2_X1 U586 ( .A1(G101), .A2(n886), .ZN(n530) );
  XOR2_X1 U587 ( .A(KEYINPUT23), .B(n530), .Z(n531) );
  NAND2_X1 U588 ( .A1(n532), .A2(n531), .ZN(n536) );
  NAND2_X1 U589 ( .A1(G113), .A2(n893), .ZN(n534) );
  NAND2_X1 U590 ( .A1(G137), .A2(n884), .ZN(n533) );
  NAND2_X1 U591 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X2 U592 ( .A1(n536), .A2(n535), .ZN(G160) );
  INV_X1 U593 ( .A(G651), .ZN(n545) );
  XNOR2_X1 U594 ( .A(G543), .B(KEYINPUT0), .ZN(n537) );
  XNOR2_X1 U595 ( .A(n537), .B(KEYINPUT65), .ZN(n650) );
  NOR2_X1 U596 ( .A1(n545), .A2(n650), .ZN(n538) );
  XNOR2_X1 U597 ( .A(KEYINPUT66), .B(n538), .ZN(n607) );
  BUF_X1 U598 ( .A(n607), .Z(n644) );
  NAND2_X1 U599 ( .A1(n644), .A2(G76), .ZN(n542) );
  XOR2_X1 U600 ( .A(KEYINPUT73), .B(KEYINPUT4), .Z(n540) );
  NAND2_X1 U601 ( .A1(G89), .A2(n658), .ZN(n539) );
  XNOR2_X1 U602 ( .A(n540), .B(n539), .ZN(n541) );
  NAND2_X1 U603 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U604 ( .A(n543), .B(KEYINPUT74), .ZN(n544) );
  XNOR2_X1 U605 ( .A(n544), .B(KEYINPUT5), .ZN(n553) );
  XNOR2_X1 U606 ( .A(KEYINPUT76), .B(KEYINPUT6), .ZN(n551) );
  NOR2_X1 U607 ( .A1(G651), .A2(n650), .ZN(n657) );
  NAND2_X1 U608 ( .A1(n657), .A2(G51), .ZN(n549) );
  NOR2_X1 U609 ( .A1(G543), .A2(n545), .ZN(n546) );
  XOR2_X1 U610 ( .A(KEYINPUT1), .B(n546), .Z(n656) );
  NAND2_X1 U611 ( .A1(n656), .A2(G63), .ZN(n547) );
  XOR2_X1 U612 ( .A(KEYINPUT75), .B(n547), .Z(n548) );
  NAND2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U614 ( .A(n551), .B(n550), .Z(n552) );
  NAND2_X1 U615 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U616 ( .A(n554), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U617 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U618 ( .A1(n658), .A2(G88), .ZN(n561) );
  NAND2_X1 U619 ( .A1(G62), .A2(n656), .ZN(n556) );
  NAND2_X1 U620 ( .A1(G50), .A2(n657), .ZN(n555) );
  NAND2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n559) );
  NAND2_X1 U622 ( .A1(G75), .A2(n644), .ZN(n557) );
  XNOR2_X1 U623 ( .A(KEYINPUT81), .B(n557), .ZN(n558) );
  NOR2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U625 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U626 ( .A(KEYINPUT82), .B(n562), .Z(G166) );
  INV_X1 U627 ( .A(G166), .ZN(G303) );
  NAND2_X1 U628 ( .A1(G64), .A2(n656), .ZN(n564) );
  NAND2_X1 U629 ( .A1(G52), .A2(n657), .ZN(n563) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n569) );
  NAND2_X1 U631 ( .A1(G90), .A2(n658), .ZN(n566) );
  NAND2_X1 U632 ( .A1(G77), .A2(n644), .ZN(n565) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U634 ( .A(KEYINPUT9), .B(n567), .Z(n568) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(G171) );
  XOR2_X1 U636 ( .A(G2446), .B(G2451), .Z(n571) );
  XNOR2_X1 U637 ( .A(G2454), .B(KEYINPUT103), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(n578) );
  XOR2_X1 U639 ( .A(G2438), .B(G2430), .Z(n573) );
  XNOR2_X1 U640 ( .A(G2435), .B(G2443), .ZN(n572) );
  XNOR2_X1 U641 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U642 ( .A(n574), .B(G2427), .Z(n576) );
  XNOR2_X1 U643 ( .A(G1341), .B(G1348), .ZN(n575) );
  XNOR2_X1 U644 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U645 ( .A(n578), .B(n577), .ZN(n579) );
  AND2_X1 U646 ( .A1(n579), .A2(G14), .ZN(G401) );
  AND2_X1 U647 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U648 ( .A1(G123), .A2(n890), .ZN(n580) );
  XNOR2_X1 U649 ( .A(n580), .B(KEYINPUT18), .ZN(n583) );
  NAND2_X1 U650 ( .A1(G99), .A2(n886), .ZN(n581) );
  XNOR2_X1 U651 ( .A(n581), .B(KEYINPUT78), .ZN(n582) );
  NAND2_X1 U652 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U653 ( .A1(G111), .A2(n893), .ZN(n585) );
  NAND2_X1 U654 ( .A1(G135), .A2(n884), .ZN(n584) );
  NAND2_X1 U655 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U656 ( .A1(n587), .A2(n586), .ZN(n923) );
  XNOR2_X1 U657 ( .A(n923), .B(G2096), .ZN(n588) );
  XNOR2_X1 U658 ( .A(n588), .B(KEYINPUT79), .ZN(n589) );
  OR2_X1 U659 ( .A1(G2100), .A2(n589), .ZN(G156) );
  INV_X1 U660 ( .A(G57), .ZN(G237) );
  INV_X1 U661 ( .A(G132), .ZN(G219) );
  INV_X1 U662 ( .A(G82), .ZN(G220) );
  XOR2_X1 U663 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n591) );
  NAND2_X1 U664 ( .A1(G7), .A2(G661), .ZN(n590) );
  XNOR2_X1 U665 ( .A(n591), .B(n590), .ZN(G223) );
  INV_X1 U666 ( .A(G223), .ZN(n837) );
  NAND2_X1 U667 ( .A1(n837), .A2(G567), .ZN(n592) );
  XOR2_X1 U668 ( .A(KEYINPUT11), .B(n592), .Z(G234) );
  NAND2_X1 U669 ( .A1(n656), .A2(G56), .ZN(n593) );
  XNOR2_X1 U670 ( .A(n593), .B(KEYINPUT14), .ZN(n595) );
  NAND2_X1 U671 ( .A1(G43), .A2(n657), .ZN(n594) );
  NAND2_X1 U672 ( .A1(n595), .A2(n594), .ZN(n603) );
  NAND2_X1 U673 ( .A1(n658), .A2(G81), .ZN(n596) );
  XNOR2_X1 U674 ( .A(n596), .B(KEYINPUT12), .ZN(n598) );
  NAND2_X1 U675 ( .A1(G68), .A2(n607), .ZN(n597) );
  NAND2_X1 U676 ( .A1(n598), .A2(n597), .ZN(n601) );
  XOR2_X1 U677 ( .A(KEYINPUT71), .B(n604), .Z(n705) );
  NAND2_X1 U678 ( .A1(n705), .A2(G860), .ZN(G153) );
  INV_X1 U679 ( .A(G171), .ZN(G301) );
  NAND2_X1 U680 ( .A1(G868), .A2(G301), .ZN(n615) );
  NAND2_X1 U681 ( .A1(G92), .A2(n658), .ZN(n612) );
  NAND2_X1 U682 ( .A1(G66), .A2(n656), .ZN(n606) );
  NAND2_X1 U683 ( .A1(G54), .A2(n657), .ZN(n605) );
  NAND2_X1 U684 ( .A1(n606), .A2(n605), .ZN(n610) );
  NAND2_X1 U685 ( .A1(n607), .A2(G79), .ZN(n608) );
  XOR2_X1 U686 ( .A(KEYINPUT72), .B(n608), .Z(n609) );
  NOR2_X1 U687 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U688 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X2 U689 ( .A(n613), .B(KEYINPUT15), .ZN(n976) );
  INV_X1 U690 ( .A(n976), .ZN(n708) );
  INV_X1 U691 ( .A(G868), .ZN(n623) );
  NAND2_X1 U692 ( .A1(n708), .A2(n623), .ZN(n614) );
  NAND2_X1 U693 ( .A1(n615), .A2(n614), .ZN(G284) );
  NAND2_X1 U694 ( .A1(n657), .A2(G53), .ZN(n618) );
  NAND2_X1 U695 ( .A1(G65), .A2(n656), .ZN(n616) );
  XOR2_X1 U696 ( .A(KEYINPUT67), .B(n616), .Z(n617) );
  NAND2_X1 U697 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U698 ( .A1(G91), .A2(n658), .ZN(n620) );
  NAND2_X1 U699 ( .A1(G78), .A2(n644), .ZN(n619) );
  NAND2_X1 U700 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n979) );
  XOR2_X1 U702 ( .A(n979), .B(KEYINPUT68), .Z(G299) );
  NOR2_X1 U703 ( .A1(G299), .A2(G868), .ZN(n625) );
  NOR2_X1 U704 ( .A1(G286), .A2(n623), .ZN(n624) );
  NOR2_X1 U705 ( .A1(n625), .A2(n624), .ZN(G297) );
  INV_X1 U706 ( .A(G860), .ZN(n633) );
  NAND2_X1 U707 ( .A1(n633), .A2(G559), .ZN(n626) );
  NAND2_X1 U708 ( .A1(n626), .A2(n976), .ZN(n627) );
  XNOR2_X1 U709 ( .A(n627), .B(KEYINPUT16), .ZN(n628) );
  XOR2_X1 U710 ( .A(KEYINPUT77), .B(n628), .Z(G148) );
  OR2_X1 U711 ( .A1(G559), .A2(n708), .ZN(n629) );
  NAND2_X1 U712 ( .A1(n629), .A2(G868), .ZN(n631) );
  OR2_X1 U713 ( .A1(n705), .A2(G868), .ZN(n630) );
  NAND2_X1 U714 ( .A1(n631), .A2(n630), .ZN(G282) );
  NAND2_X1 U715 ( .A1(G559), .A2(n976), .ZN(n632) );
  XNOR2_X1 U716 ( .A(n632), .B(n705), .ZN(n670) );
  NAND2_X1 U717 ( .A1(n633), .A2(n670), .ZN(n641) );
  NAND2_X1 U718 ( .A1(G55), .A2(n657), .ZN(n634) );
  XNOR2_X1 U719 ( .A(n634), .B(KEYINPUT80), .ZN(n636) );
  NAND2_X1 U720 ( .A1(n656), .A2(G67), .ZN(n635) );
  NAND2_X1 U721 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U722 ( .A1(G93), .A2(n658), .ZN(n638) );
  NAND2_X1 U723 ( .A1(G80), .A2(n644), .ZN(n637) );
  NAND2_X1 U724 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U725 ( .A1(n640), .A2(n639), .ZN(n672) );
  XOR2_X1 U726 ( .A(n641), .B(n672), .Z(G145) );
  NAND2_X1 U727 ( .A1(G48), .A2(n657), .ZN(n643) );
  NAND2_X1 U728 ( .A1(G86), .A2(n658), .ZN(n642) );
  NAND2_X1 U729 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U730 ( .A1(n644), .A2(G73), .ZN(n645) );
  XOR2_X1 U731 ( .A(KEYINPUT2), .B(n645), .Z(n646) );
  NOR2_X1 U732 ( .A1(n647), .A2(n646), .ZN(n649) );
  NAND2_X1 U733 ( .A1(n656), .A2(G61), .ZN(n648) );
  NAND2_X1 U734 ( .A1(n649), .A2(n648), .ZN(G305) );
  NAND2_X1 U735 ( .A1(G49), .A2(n657), .ZN(n652) );
  NAND2_X1 U736 ( .A1(G87), .A2(n650), .ZN(n651) );
  NAND2_X1 U737 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U738 ( .A1(n656), .A2(n653), .ZN(n655) );
  NAND2_X1 U739 ( .A1(G651), .A2(G74), .ZN(n654) );
  NAND2_X1 U740 ( .A1(n655), .A2(n654), .ZN(G288) );
  AND2_X1 U741 ( .A1(n656), .A2(G60), .ZN(n662) );
  NAND2_X1 U742 ( .A1(G47), .A2(n657), .ZN(n660) );
  NAND2_X1 U743 ( .A1(G85), .A2(n658), .ZN(n659) );
  NAND2_X1 U744 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U745 ( .A1(n662), .A2(n661), .ZN(n664) );
  NAND2_X1 U746 ( .A1(G72), .A2(n644), .ZN(n663) );
  NAND2_X1 U747 ( .A1(n664), .A2(n663), .ZN(G290) );
  XNOR2_X1 U748 ( .A(G303), .B(G299), .ZN(n669) );
  XNOR2_X1 U749 ( .A(n672), .B(G305), .ZN(n667) );
  XOR2_X1 U750 ( .A(KEYINPUT19), .B(G290), .Z(n665) );
  XNOR2_X1 U751 ( .A(G288), .B(n665), .ZN(n666) );
  XNOR2_X1 U752 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U753 ( .A(n669), .B(n668), .ZN(n911) );
  XNOR2_X1 U754 ( .A(n670), .B(n911), .ZN(n671) );
  NAND2_X1 U755 ( .A1(n671), .A2(G868), .ZN(n674) );
  OR2_X1 U756 ( .A1(G868), .A2(n672), .ZN(n673) );
  NAND2_X1 U757 ( .A1(n674), .A2(n673), .ZN(G295) );
  NAND2_X1 U758 ( .A1(G2084), .A2(G2078), .ZN(n675) );
  XNOR2_X1 U759 ( .A(n675), .B(KEYINPUT20), .ZN(n676) );
  XNOR2_X1 U760 ( .A(KEYINPUT83), .B(n676), .ZN(n677) );
  NAND2_X1 U761 ( .A1(n677), .A2(G2090), .ZN(n678) );
  XNOR2_X1 U762 ( .A(KEYINPUT21), .B(n678), .ZN(n679) );
  NAND2_X1 U763 ( .A1(n679), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U764 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U765 ( .A1(G220), .A2(G219), .ZN(n680) );
  XOR2_X1 U766 ( .A(KEYINPUT22), .B(n680), .Z(n681) );
  NOR2_X1 U767 ( .A1(G218), .A2(n681), .ZN(n682) );
  NAND2_X1 U768 ( .A1(G96), .A2(n682), .ZN(n842) );
  NAND2_X1 U769 ( .A1(n842), .A2(G2106), .ZN(n686) );
  NAND2_X1 U770 ( .A1(G120), .A2(G108), .ZN(n683) );
  NOR2_X1 U771 ( .A1(G237), .A2(n683), .ZN(n684) );
  NAND2_X1 U772 ( .A1(G69), .A2(n684), .ZN(n843) );
  NAND2_X1 U773 ( .A1(n843), .A2(G567), .ZN(n685) );
  NAND2_X1 U774 ( .A1(n686), .A2(n685), .ZN(n844) );
  NAND2_X1 U775 ( .A1(G483), .A2(G661), .ZN(n687) );
  NOR2_X1 U776 ( .A1(n844), .A2(n687), .ZN(n841) );
  NAND2_X1 U777 ( .A1(n841), .A2(G36), .ZN(n688) );
  XNOR2_X1 U778 ( .A(KEYINPUT84), .B(n688), .ZN(G176) );
  XNOR2_X2 U779 ( .A(n736), .B(KEYINPUT93), .ZN(n722) );
  XOR2_X1 U780 ( .A(KEYINPUT93), .B(n736), .Z(n692) );
  NAND2_X1 U781 ( .A1(n692), .A2(G1956), .ZN(n693) );
  NAND2_X1 U782 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U783 ( .A(n695), .B(KEYINPUT95), .ZN(n712) );
  XNOR2_X1 U784 ( .A(n697), .B(n696), .ZN(n716) );
  NAND2_X1 U785 ( .A1(n736), .A2(G1348), .ZN(n699) );
  NAND2_X1 U786 ( .A1(G2067), .A2(n722), .ZN(n698) );
  NAND2_X1 U787 ( .A1(n699), .A2(n698), .ZN(n709) );
  OR2_X1 U788 ( .A1(n709), .A2(n708), .ZN(n707) );
  INV_X1 U789 ( .A(n736), .ZN(n719) );
  XNOR2_X1 U790 ( .A(G1996), .B(KEYINPUT96), .ZN(n951) );
  NAND2_X1 U791 ( .A1(n719), .A2(n951), .ZN(n700) );
  XNOR2_X1 U792 ( .A(n700), .B(KEYINPUT26), .ZN(n702) );
  NAND2_X1 U793 ( .A1(G1341), .A2(n736), .ZN(n701) );
  NAND2_X1 U794 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U795 ( .A(KEYINPUT97), .B(n703), .ZN(n704) );
  NAND2_X1 U796 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U797 ( .A1(n707), .A2(n706), .ZN(n711) );
  NAND2_X1 U798 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U799 ( .A1(n711), .A2(n710), .ZN(n714) );
  NAND2_X1 U800 ( .A1(n979), .A2(n712), .ZN(n713) );
  NAND2_X1 U801 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U802 ( .A1(n716), .A2(n715), .ZN(n718) );
  NOR2_X1 U803 ( .A1(n719), .A2(G1961), .ZN(n720) );
  XOR2_X1 U804 ( .A(KEYINPUT92), .B(n720), .Z(n724) );
  XNOR2_X1 U805 ( .A(G2078), .B(KEYINPUT25), .ZN(n721) );
  XNOR2_X1 U806 ( .A(n721), .B(KEYINPUT94), .ZN(n950) );
  NAND2_X1 U807 ( .A1(n950), .A2(n722), .ZN(n723) );
  NAND2_X1 U808 ( .A1(n724), .A2(n723), .ZN(n730) );
  NAND2_X1 U809 ( .A1(n730), .A2(G171), .ZN(n725) );
  NAND2_X1 U810 ( .A1(n726), .A2(n725), .ZN(n735) );
  NAND2_X1 U811 ( .A1(G8), .A2(n736), .ZN(n810) );
  NOR2_X1 U812 ( .A1(G1966), .A2(n810), .ZN(n749) );
  NOR2_X1 U813 ( .A1(G2084), .A2(n736), .ZN(n746) );
  NOR2_X1 U814 ( .A1(n749), .A2(n746), .ZN(n727) );
  NAND2_X1 U815 ( .A1(G8), .A2(n727), .ZN(n728) );
  XNOR2_X1 U816 ( .A(KEYINPUT30), .B(n728), .ZN(n729) );
  NOR2_X1 U817 ( .A1(G168), .A2(n729), .ZN(n732) );
  NOR2_X1 U818 ( .A1(G171), .A2(n730), .ZN(n731) );
  NOR2_X1 U819 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U820 ( .A(KEYINPUT31), .B(n733), .Z(n734) );
  NAND2_X1 U821 ( .A1(n735), .A2(n734), .ZN(n747) );
  NAND2_X1 U822 ( .A1(n747), .A2(G286), .ZN(n741) );
  NOR2_X1 U823 ( .A1(G1971), .A2(n810), .ZN(n738) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n736), .ZN(n737) );
  NOR2_X1 U825 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U826 ( .A1(G303), .A2(n739), .ZN(n740) );
  NAND2_X1 U827 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U828 ( .A(n742), .B(KEYINPUT98), .ZN(n743) );
  NAND2_X1 U829 ( .A1(n743), .A2(G8), .ZN(n745) );
  XOR2_X1 U830 ( .A(KEYINPUT99), .B(KEYINPUT32), .Z(n744) );
  XNOR2_X1 U831 ( .A(n745), .B(n744), .ZN(n753) );
  NAND2_X1 U832 ( .A1(G8), .A2(n746), .ZN(n751) );
  INV_X1 U833 ( .A(n747), .ZN(n748) );
  NOR2_X1 U834 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U835 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U836 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U837 ( .A(n754), .B(KEYINPUT100), .ZN(n809) );
  NOR2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n762) );
  NOR2_X1 U839 ( .A1(G303), .A2(G1971), .ZN(n755) );
  NOR2_X1 U840 ( .A1(n762), .A2(n755), .ZN(n985) );
  AND2_X2 U841 ( .A1(n809), .A2(n985), .ZN(n757) );
  INV_X1 U842 ( .A(KEYINPUT101), .ZN(n756) );
  XNOR2_X1 U843 ( .A(n757), .B(n756), .ZN(n760) );
  NAND2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n980) );
  INV_X1 U845 ( .A(n810), .ZN(n758) );
  NAND2_X1 U846 ( .A1(n980), .A2(n758), .ZN(n759) );
  NOR2_X1 U847 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U848 ( .A1(n761), .A2(KEYINPUT33), .ZN(n765) );
  NAND2_X1 U849 ( .A1(n762), .A2(KEYINPUT33), .ZN(n763) );
  NOR2_X1 U850 ( .A1(n763), .A2(n810), .ZN(n764) );
  NOR2_X1 U851 ( .A1(n765), .A2(n764), .ZN(n800) );
  XOR2_X1 U852 ( .A(G1981), .B(G305), .Z(n973) );
  NAND2_X1 U853 ( .A1(G160), .A2(G40), .ZN(n766) );
  NOR2_X1 U854 ( .A1(n767), .A2(n766), .ZN(n833) );
  NAND2_X1 U855 ( .A1(G105), .A2(n886), .ZN(n768) );
  XNOR2_X1 U856 ( .A(n768), .B(KEYINPUT38), .ZN(n776) );
  NAND2_X1 U857 ( .A1(n893), .A2(G117), .ZN(n769) );
  XNOR2_X1 U858 ( .A(n769), .B(KEYINPUT88), .ZN(n771) );
  NAND2_X1 U859 ( .A1(G129), .A2(n890), .ZN(n770) );
  NAND2_X1 U860 ( .A1(n771), .A2(n770), .ZN(n774) );
  NAND2_X1 U861 ( .A1(G141), .A2(n884), .ZN(n772) );
  XNOR2_X1 U862 ( .A(KEYINPUT89), .B(n772), .ZN(n773) );
  NOR2_X1 U863 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U864 ( .A1(n776), .A2(n775), .ZN(n882) );
  NAND2_X1 U865 ( .A1(G1996), .A2(n882), .ZN(n785) );
  NAND2_X1 U866 ( .A1(G95), .A2(n886), .ZN(n778) );
  NAND2_X1 U867 ( .A1(G119), .A2(n890), .ZN(n777) );
  NAND2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n781) );
  NAND2_X1 U869 ( .A1(G107), .A2(n893), .ZN(n779) );
  XNOR2_X1 U870 ( .A(KEYINPUT87), .B(n779), .ZN(n780) );
  NOR2_X1 U871 ( .A1(n781), .A2(n780), .ZN(n783) );
  NAND2_X1 U872 ( .A1(n884), .A2(G131), .ZN(n782) );
  NAND2_X1 U873 ( .A1(n783), .A2(n782), .ZN(n907) );
  NAND2_X1 U874 ( .A1(G1991), .A2(n907), .ZN(n784) );
  NAND2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n928) );
  NAND2_X1 U876 ( .A1(n833), .A2(n928), .ZN(n822) );
  XNOR2_X1 U877 ( .A(G1986), .B(G290), .ZN(n987) );
  NAND2_X1 U878 ( .A1(n833), .A2(n987), .ZN(n786) );
  NAND2_X1 U879 ( .A1(n822), .A2(n786), .ZN(n815) );
  INV_X1 U880 ( .A(n815), .ZN(n787) );
  AND2_X1 U881 ( .A1(n973), .A2(n787), .ZN(n798) );
  XNOR2_X1 U882 ( .A(G2067), .B(KEYINPUT37), .ZN(n788) );
  XNOR2_X1 U883 ( .A(n788), .B(KEYINPUT86), .ZN(n830) );
  NAND2_X1 U884 ( .A1(G104), .A2(n886), .ZN(n790) );
  NAND2_X1 U885 ( .A1(G140), .A2(n884), .ZN(n789) );
  NAND2_X1 U886 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U887 ( .A(KEYINPUT34), .B(n791), .ZN(n796) );
  NAND2_X1 U888 ( .A1(G116), .A2(n893), .ZN(n793) );
  NAND2_X1 U889 ( .A1(G128), .A2(n890), .ZN(n792) );
  NAND2_X1 U890 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U891 ( .A(KEYINPUT35), .B(n794), .Z(n795) );
  NOR2_X1 U892 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U893 ( .A(KEYINPUT36), .B(n797), .ZN(n898) );
  NOR2_X1 U894 ( .A1(n830), .A2(n898), .ZN(n940) );
  NAND2_X1 U895 ( .A1(n833), .A2(n940), .ZN(n828) );
  AND2_X1 U896 ( .A1(n798), .A2(n828), .ZN(n799) );
  NAND2_X1 U897 ( .A1(n800), .A2(n799), .ZN(n819) );
  INV_X1 U898 ( .A(n828), .ZN(n817) );
  NOR2_X1 U899 ( .A1(G303), .A2(G2090), .ZN(n801) );
  NAND2_X1 U900 ( .A1(G8), .A2(n801), .ZN(n807) );
  NOR2_X1 U901 ( .A1(G1981), .A2(G305), .ZN(n802) );
  XOR2_X1 U902 ( .A(n802), .B(KEYINPUT24), .Z(n803) );
  XNOR2_X1 U903 ( .A(KEYINPUT90), .B(n803), .ZN(n804) );
  NOR2_X1 U904 ( .A1(n810), .A2(n804), .ZN(n805) );
  XOR2_X1 U905 ( .A(KEYINPUT91), .B(n805), .Z(n811) );
  INV_X1 U906 ( .A(n811), .ZN(n806) );
  AND2_X1 U907 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U908 ( .A1(n809), .A2(n808), .ZN(n813) );
  OR2_X1 U909 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U910 ( .A1(n813), .A2(n812), .ZN(n814) );
  OR2_X1 U911 ( .A1(n815), .A2(n814), .ZN(n816) );
  OR2_X1 U912 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U913 ( .A(n821), .B(n820), .ZN(n835) );
  NOR2_X1 U914 ( .A1(G1996), .A2(n882), .ZN(n932) );
  INV_X1 U915 ( .A(n822), .ZN(n825) );
  NOR2_X1 U916 ( .A1(G1991), .A2(n907), .ZN(n924) );
  NOR2_X1 U917 ( .A1(G1986), .A2(G290), .ZN(n823) );
  NOR2_X1 U918 ( .A1(n924), .A2(n823), .ZN(n824) );
  NOR2_X1 U919 ( .A1(n825), .A2(n824), .ZN(n826) );
  NOR2_X1 U920 ( .A1(n932), .A2(n826), .ZN(n827) );
  XNOR2_X1 U921 ( .A(KEYINPUT39), .B(n827), .ZN(n829) );
  NAND2_X1 U922 ( .A1(n829), .A2(n828), .ZN(n831) );
  NAND2_X1 U923 ( .A1(n830), .A2(n898), .ZN(n929) );
  NAND2_X1 U924 ( .A1(n831), .A2(n929), .ZN(n832) );
  NAND2_X1 U925 ( .A1(n833), .A2(n832), .ZN(n834) );
  NAND2_X1 U926 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U927 ( .A(n836), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n837), .ZN(G217) );
  NAND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n838) );
  XOR2_X1 U930 ( .A(KEYINPUT104), .B(n838), .Z(n839) );
  NAND2_X1 U931 ( .A1(G661), .A2(n839), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U933 ( .A1(n841), .A2(n840), .ZN(G188) );
  XNOR2_X1 U934 ( .A(G108), .B(KEYINPUT117), .ZN(G238) );
  INV_X1 U936 ( .A(G120), .ZN(G236) );
  INV_X1 U937 ( .A(G96), .ZN(G221) );
  NOR2_X1 U938 ( .A1(n843), .A2(n842), .ZN(G325) );
  INV_X1 U939 ( .A(G325), .ZN(G261) );
  INV_X1 U940 ( .A(n844), .ZN(G319) );
  XOR2_X1 U941 ( .A(KEYINPUT41), .B(G1961), .Z(n846) );
  XNOR2_X1 U942 ( .A(G1986), .B(G1981), .ZN(n845) );
  XNOR2_X1 U943 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U944 ( .A(n847), .B(KEYINPUT106), .Z(n849) );
  XNOR2_X1 U945 ( .A(G1996), .B(G1991), .ZN(n848) );
  XNOR2_X1 U946 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U947 ( .A(G1956), .B(G1966), .Z(n851) );
  XNOR2_X1 U948 ( .A(G1976), .B(G1971), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U950 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U951 ( .A(KEYINPUT107), .B(G2474), .ZN(n854) );
  XNOR2_X1 U952 ( .A(n855), .B(n854), .ZN(G229) );
  XOR2_X1 U953 ( .A(G2678), .B(G2084), .Z(n857) );
  XNOR2_X1 U954 ( .A(G2078), .B(G2072), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U956 ( .A(n858), .B(G2100), .Z(n860) );
  XNOR2_X1 U957 ( .A(G2067), .B(G2090), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U959 ( .A(G2096), .B(KEYINPUT105), .Z(n862) );
  XNOR2_X1 U960 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U962 ( .A(n864), .B(n863), .Z(G227) );
  NAND2_X1 U963 ( .A1(G112), .A2(n893), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n865), .B(KEYINPUT108), .ZN(n872) );
  NAND2_X1 U965 ( .A1(G100), .A2(n886), .ZN(n867) );
  NAND2_X1 U966 ( .A1(G136), .A2(n884), .ZN(n866) );
  NAND2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n870) );
  NAND2_X1 U968 ( .A1(n890), .A2(G124), .ZN(n868) );
  XOR2_X1 U969 ( .A(KEYINPUT44), .B(n868), .Z(n869) );
  NOR2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n871) );
  NAND2_X1 U971 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U972 ( .A(KEYINPUT109), .B(n873), .ZN(G162) );
  NAND2_X1 U973 ( .A1(G103), .A2(n886), .ZN(n875) );
  NAND2_X1 U974 ( .A1(G139), .A2(n884), .ZN(n874) );
  NAND2_X1 U975 ( .A1(n875), .A2(n874), .ZN(n880) );
  NAND2_X1 U976 ( .A1(G115), .A2(n893), .ZN(n877) );
  NAND2_X1 U977 ( .A1(G127), .A2(n890), .ZN(n876) );
  NAND2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U979 ( .A(KEYINPUT47), .B(n878), .Z(n879) );
  NOR2_X1 U980 ( .A1(n880), .A2(n879), .ZN(n935) );
  XOR2_X1 U981 ( .A(G164), .B(n935), .Z(n881) );
  XNOR2_X1 U982 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U983 ( .A(G162), .B(n883), .ZN(n900) );
  NAND2_X1 U984 ( .A1(n884), .A2(G142), .ZN(n885) );
  XOR2_X1 U985 ( .A(KEYINPUT111), .B(n885), .Z(n888) );
  NAND2_X1 U986 ( .A1(n886), .A2(G106), .ZN(n887) );
  NAND2_X1 U987 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U988 ( .A(n889), .B(KEYINPUT45), .ZN(n892) );
  NAND2_X1 U989 ( .A1(G130), .A2(n890), .ZN(n891) );
  NAND2_X1 U990 ( .A1(n892), .A2(n891), .ZN(n896) );
  NAND2_X1 U991 ( .A1(n893), .A2(G118), .ZN(n894) );
  XOR2_X1 U992 ( .A(KEYINPUT110), .B(n894), .Z(n895) );
  NOR2_X1 U993 ( .A1(n896), .A2(n895), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n909) );
  XOR2_X1 U996 ( .A(KEYINPUT112), .B(KEYINPUT46), .Z(n902) );
  XNOR2_X1 U997 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U999 ( .A(n903), .B(KEYINPUT48), .Z(n905) );
  XNOR2_X1 U1000 ( .A(G160), .B(n923), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n910), .ZN(G395) );
  XOR2_X1 U1005 ( .A(n911), .B(G286), .Z(n913) );
  XNOR2_X1 U1006 ( .A(n976), .B(n705), .ZN(n912) );
  XNOR2_X1 U1007 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1008 ( .A(n914), .B(G171), .ZN(n915) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n915), .ZN(G397) );
  NOR2_X1 U1010 ( .A1(G229), .A2(G227), .ZN(n916) );
  XNOR2_X1 U1011 ( .A(KEYINPUT49), .B(n916), .ZN(n917) );
  NOR2_X1 U1012 ( .A1(G401), .A2(n917), .ZN(n918) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n918), .ZN(n921) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(KEYINPUT115), .B(n919), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1017 ( .A(KEYINPUT116), .B(n922), .ZN(G308) );
  INV_X1 U1018 ( .A(G308), .ZN(G225) );
  INV_X1 U1019 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1020 ( .A(G160), .B(G2084), .ZN(n926) );
  NOR2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(n930) );
  NAND2_X1 U1024 ( .A1(n930), .A2(n929), .ZN(n944) );
  XOR2_X1 U1025 ( .A(G2090), .B(G162), .Z(n931) );
  NOR2_X1 U1026 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1027 ( .A(KEYINPUT51), .B(n933), .Z(n934) );
  XNOR2_X1 U1028 ( .A(KEYINPUT118), .B(n934), .ZN(n942) );
  XOR2_X1 U1029 ( .A(G2072), .B(n935), .Z(n937) );
  XOR2_X1 U1030 ( .A(G164), .B(G2078), .Z(n936) );
  NOR2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1032 ( .A(KEYINPUT50), .B(n938), .Z(n939) );
  NOR2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1034 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1035 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1036 ( .A(KEYINPUT52), .B(n945), .ZN(n946) );
  INV_X1 U1037 ( .A(KEYINPUT55), .ZN(n969) );
  NAND2_X1 U1038 ( .A1(n946), .A2(n969), .ZN(n947) );
  NAND2_X1 U1039 ( .A1(n947), .A2(G29), .ZN(n1029) );
  XNOR2_X1 U1040 ( .A(KEYINPUT54), .B(G34), .ZN(n948) );
  XNOR2_X1 U1041 ( .A(n948), .B(KEYINPUT121), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(G2084), .B(n949), .ZN(n967) );
  XNOR2_X1 U1043 ( .A(G2090), .B(G35), .ZN(n965) );
  XNOR2_X1 U1044 ( .A(n950), .B(G27), .ZN(n953) );
  XOR2_X1 U1045 ( .A(G32), .B(n951), .Z(n952) );
  NAND2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(n954), .B(KEYINPUT120), .ZN(n962) );
  XNOR2_X1 U1048 ( .A(G25), .B(G1991), .ZN(n955) );
  XNOR2_X1 U1049 ( .A(n955), .B(KEYINPUT119), .ZN(n960) );
  XOR2_X1 U1050 ( .A(G2072), .B(G33), .Z(n956) );
  NAND2_X1 U1051 ( .A1(n956), .A2(G28), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(G26), .B(G2067), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(KEYINPUT53), .B(n963), .ZN(n964) );
  NOR2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1058 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1059 ( .A(n969), .B(n968), .ZN(n971) );
  INV_X1 U1060 ( .A(G29), .ZN(n970) );
  NAND2_X1 U1061 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1062 ( .A1(G11), .A2(n972), .ZN(n1027) );
  XNOR2_X1 U1063 ( .A(G16), .B(KEYINPUT56), .ZN(n995) );
  XNOR2_X1 U1064 ( .A(G1966), .B(G168), .ZN(n974) );
  NAND2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1066 ( .A(n975), .B(KEYINPUT57), .ZN(n993) );
  XNOR2_X1 U1067 ( .A(n976), .B(G1348), .ZN(n978) );
  XNOR2_X1 U1068 ( .A(G171), .B(G1961), .ZN(n977) );
  NAND2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n991) );
  XNOR2_X1 U1070 ( .A(n705), .B(G1341), .ZN(n989) );
  XNOR2_X1 U1071 ( .A(G1956), .B(n979), .ZN(n981) );
  NAND2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n983) );
  AND2_X1 U1073 ( .A1(G303), .A2(G1971), .ZN(n982) );
  NOR2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1078 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1079 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1080 ( .A1(n995), .A2(n994), .ZN(n1025) );
  INV_X1 U1081 ( .A(G16), .ZN(n1023) );
  XNOR2_X1 U1082 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n1021) );
  XNOR2_X1 U1083 ( .A(G1348), .B(KEYINPUT59), .ZN(n996) );
  XNOR2_X1 U1084 ( .A(n996), .B(G4), .ZN(n1000) );
  XNOR2_X1 U1085 ( .A(G1981), .B(G6), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(G1956), .B(G20), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1003) );
  XOR2_X1 U1089 ( .A(KEYINPUT123), .B(G1341), .Z(n1001) );
  XNOR2_X1 U1090 ( .A(G19), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(KEYINPUT60), .B(n1004), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(n1005), .B(KEYINPUT124), .ZN(n1019) );
  XOR2_X1 U1094 ( .A(G1966), .B(G21), .Z(n1014) );
  XOR2_X1 U1095 ( .A(G1976), .B(G23), .Z(n1008) );
  XOR2_X1 U1096 ( .A(G24), .B(KEYINPUT126), .Z(n1006) );
  XNOR2_X1 U1097 ( .A(n1006), .B(G1986), .ZN(n1007) );
  NAND2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1011) );
  XOR2_X1 U1099 ( .A(KEYINPUT125), .B(G1971), .Z(n1009) );
  XNOR2_X1 U1100 ( .A(G22), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1102 ( .A(KEYINPUT58), .B(n1012), .ZN(n1013) );
  NAND2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(KEYINPUT122), .B(G1961), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(G5), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1108 ( .A(n1021), .B(n1020), .ZN(n1022) );
  NAND2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1112 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1030), .Z(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

