

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799;

  XNOR2_X2 U374 ( .A(n509), .B(n510), .ZN(n684) );
  XNOR2_X2 U375 ( .A(n371), .B(n370), .ZN(n510) );
  AND2_X2 U376 ( .A1(n463), .A2(n412), .ZN(n410) );
  XNOR2_X2 U377 ( .A(n475), .B(n474), .ZN(n508) );
  NOR2_X1 U378 ( .A1(G953), .A2(G237), .ZN(n551) );
  NAND2_X1 U379 ( .A1(n421), .A2(n650), .ZN(n423) );
  INV_X2 U380 ( .A(KEYINPUT64), .ZN(n476) );
  XNOR2_X1 U381 ( .A(n532), .B(KEYINPUT31), .ZN(n659) );
  XNOR2_X1 U382 ( .A(n606), .B(KEYINPUT40), .ZN(n420) );
  AND2_X2 U383 ( .A1(n406), .A2(n405), .ZN(n375) );
  XNOR2_X2 U384 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n473) );
  XNOR2_X2 U385 ( .A(G107), .B(G104), .ZN(n475) );
  XNOR2_X2 U386 ( .A(G110), .B(KEYINPUT81), .ZN(n474) );
  XNOR2_X2 U387 ( .A(G113), .B(KEYINPUT75), .ZN(n501) );
  XNOR2_X1 U388 ( .A(n563), .B(KEYINPUT22), .ZN(n588) );
  INV_X1 U389 ( .A(KEYINPUT2), .ZN(n387) );
  AND2_X1 U390 ( .A1(n791), .A2(n386), .ZN(n727) );
  NAND2_X1 U391 ( .A1(n400), .A2(n398), .ZN(n428) );
  XNOR2_X1 U392 ( .A(n566), .B(KEYINPUT104), .ZN(n672) );
  INV_X1 U393 ( .A(n588), .ZN(n353) );
  AND2_X1 U394 ( .A1(n449), .A2(n448), .ZN(n447) );
  OR2_X1 U395 ( .A1(n655), .A2(G902), .ZN(n506) );
  XNOR2_X1 U396 ( .A(n372), .B(G134), .ZN(n535) );
  XNOR2_X1 U397 ( .A(n501), .B(KEYINPUT3), .ZN(n371) );
  XNOR2_X2 U398 ( .A(G143), .B(G128), .ZN(n372) );
  XNOR2_X1 U399 ( .A(KEYINPUT16), .B(G122), .ZN(n507) );
  XNOR2_X1 U400 ( .A(G119), .B(G116), .ZN(n370) );
  XNOR2_X1 U401 ( .A(KEYINPUT15), .B(G902), .ZN(n594) );
  XNOR2_X2 U402 ( .A(n558), .B(KEYINPUT101), .ZN(n781) );
  OR2_X1 U403 ( .A1(n572), .A2(n573), .ZN(n558) );
  BUF_X1 U404 ( .A(n508), .Z(n354) );
  AND2_X1 U405 ( .A1(n455), .A2(n470), .ZN(n669) );
  XNOR2_X2 U406 ( .A(n629), .B(n413), .ZN(n414) );
  NAND2_X2 U407 ( .A1(n411), .A2(n409), .ZN(n629) );
  NAND2_X1 U408 ( .A1(n415), .A2(n658), .ZN(n593) );
  INV_X1 U409 ( .A(KEYINPUT98), .ZN(n450) );
  INV_X1 U410 ( .A(n564), .ZN(n453) );
  INV_X1 U411 ( .A(n460), .ZN(n422) );
  XNOR2_X1 U412 ( .A(n610), .B(n357), .ZN(n578) );
  NAND2_X1 U413 ( .A1(n435), .A2(n434), .ZN(n433) );
  AND2_X1 U414 ( .A1(n403), .A2(n401), .ZN(n400) );
  NOR2_X1 U415 ( .A1(n593), .A2(n366), .ZN(n403) );
  NAND2_X1 U416 ( .A1(n399), .A2(KEYINPUT72), .ZN(n398) );
  NOR2_X1 U417 ( .A1(n451), .A2(n443), .ZN(n442) );
  NAND2_X1 U418 ( .A1(n453), .A2(n444), .ZN(n443) );
  XNOR2_X1 U419 ( .A(n391), .B(n390), .ZN(n534) );
  INV_X1 U420 ( .A(KEYINPUT8), .ZN(n390) );
  NOR2_X1 U421 ( .A1(n376), .A2(n460), .ZN(n404) );
  NAND2_X1 U422 ( .A1(n594), .A2(n407), .ZN(n405) );
  NOR2_X1 U423 ( .A1(n640), .A2(n639), .ZN(n424) );
  OR2_X1 U424 ( .A1(n705), .A2(G902), .ZN(n367) );
  NAND2_X1 U425 ( .A1(n453), .A2(n452), .ZN(n738) );
  XNOR2_X1 U426 ( .A(KEYINPUT69), .B(KEYINPUT0), .ZN(n530) );
  XNOR2_X1 U427 ( .A(G128), .B(G119), .ZN(n483) );
  AND2_X1 U428 ( .A1(n534), .A2(G221), .ZN(n486) );
  XNOR2_X1 U429 ( .A(G110), .B(KEYINPUT23), .ZN(n484) );
  INV_X1 U430 ( .A(KEYINPUT10), .ZN(n482) );
  NOR2_X1 U431 ( .A1(n627), .A2(n607), .ZN(n605) );
  OR2_X1 U432 ( .A1(n580), .A2(n579), .ZN(n582) );
  BUF_X1 U433 ( .A(n564), .Z(n729) );
  BUF_X1 U434 ( .A(n737), .Z(n395) );
  AND2_X1 U435 ( .A1(n621), .A2(n559), .ZN(n438) );
  NAND2_X1 U436 ( .A1(n437), .A2(n436), .ZN(n417) );
  OR2_X1 U437 ( .A1(n621), .A2(n559), .ZN(n436) );
  NAND2_X1 U438 ( .A1(n659), .A2(n438), .ZN(n437) );
  AND2_X1 U439 ( .A1(n669), .A2(n438), .ZN(n416) );
  NOR2_X1 U440 ( .A1(KEYINPUT44), .A2(KEYINPUT72), .ZN(n402) );
  NOR2_X1 U441 ( .A1(n730), .A2(n450), .ZN(n444) );
  INV_X1 U442 ( .A(n466), .ZN(n462) );
  INV_X1 U443 ( .A(KEYINPUT88), .ZN(n407) );
  NOR2_X1 U444 ( .A1(G902), .A2(G237), .ZN(n519) );
  XNOR2_X1 U445 ( .A(n369), .B(KEYINPUT92), .ZN(n521) );
  OR2_X1 U446 ( .A1(n523), .A2(n520), .ZN(n369) );
  INV_X1 U447 ( .A(G210), .ZN(n520) );
  XOR2_X1 U448 ( .A(KEYINPUT5), .B(KEYINPUT97), .Z(n499) );
  XNOR2_X1 U449 ( .A(n535), .B(n472), .ZN(n497) );
  XNOR2_X1 U450 ( .A(KEYINPUT4), .B(G131), .ZN(n472) );
  XNOR2_X1 U451 ( .A(G143), .B(G128), .ZN(n397) );
  NAND2_X1 U452 ( .A1(G237), .A2(G234), .ZN(n524) );
  XNOR2_X1 U453 ( .A(n578), .B(KEYINPUT86), .ZN(n579) );
  NAND2_X1 U454 ( .A1(n446), .A2(n450), .ZN(n445) );
  OR2_X1 U455 ( .A1(n451), .A2(n738), .ZN(n446) );
  NAND2_X1 U456 ( .A1(n521), .A2(n651), .ZN(n466) );
  OR2_X1 U457 ( .A1(n710), .A2(n464), .ZN(n463) );
  NAND2_X1 U458 ( .A1(n465), .A2(n594), .ZN(n464) );
  INV_X1 U459 ( .A(n521), .ZN(n465) );
  INV_X1 U460 ( .A(G902), .ZN(n555) );
  XNOR2_X1 U461 ( .A(G116), .B(G107), .ZN(n537) );
  XOR2_X1 U462 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n548) );
  XNOR2_X1 U463 ( .A(G122), .B(G104), .ZN(n547) );
  XNOR2_X1 U464 ( .A(G143), .B(G113), .ZN(n545) );
  XOR2_X1 U465 ( .A(G140), .B(G131), .Z(n546) );
  NAND2_X1 U466 ( .A1(n458), .A2(KEYINPUT66), .ZN(n457) );
  INV_X1 U467 ( .A(n727), .ZN(n385) );
  INV_X1 U468 ( .A(G953), .ZN(n768) );
  NOR2_X1 U469 ( .A1(n737), .A2(n738), .ZN(n419) );
  INV_X1 U470 ( .A(n578), .ZN(n645) );
  INV_X1 U471 ( .A(KEYINPUT19), .ZN(n413) );
  XNOR2_X1 U472 ( .A(n602), .B(KEYINPUT82), .ZN(n627) );
  XNOR2_X1 U473 ( .A(n599), .B(KEYINPUT106), .ZN(n425) );
  INV_X1 U474 ( .A(KEYINPUT95), .ZN(n533) );
  BUF_X1 U475 ( .A(n792), .Z(n396) );
  XNOR2_X1 U476 ( .A(n487), .B(n439), .ZN(n693) );
  XNOR2_X1 U477 ( .A(n486), .B(n469), .ZN(n487) );
  XNOR2_X1 U478 ( .A(n358), .B(n483), .ZN(n440) );
  NOR2_X1 U479 ( .A1(n396), .A2(G952), .ZN(n715) );
  INV_X1 U480 ( .A(KEYINPUT35), .ZN(n456) );
  NAND2_X1 U481 ( .A1(n353), .A2(n356), .ZN(n585) );
  BUF_X1 U482 ( .A(n659), .Z(n662) );
  NAND2_X1 U483 ( .A1(n353), .A2(n471), .ZN(n566) );
  NOR2_X1 U484 ( .A1(n601), .A2(n609), .ZN(n355) );
  XOR2_X1 U485 ( .A(n582), .B(n581), .Z(n356) );
  XOR2_X1 U486 ( .A(KEYINPUT103), .B(KEYINPUT6), .Z(n357) );
  INV_X1 U487 ( .A(n730), .ZN(n452) );
  XOR2_X1 U488 ( .A(G137), .B(G140), .Z(n358) );
  OR2_X1 U489 ( .A1(n598), .A2(n529), .ZN(n359) );
  INV_X1 U490 ( .A(KEYINPUT91), .ZN(n412) );
  AND2_X1 U491 ( .A1(n463), .A2(n466), .ZN(n360) );
  AND2_X1 U492 ( .A1(n459), .A2(n457), .ZN(n361) );
  OR2_X1 U493 ( .A1(n462), .A2(n468), .ZN(n362) );
  XNOR2_X1 U494 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n363) );
  OR2_X1 U495 ( .A1(n594), .A2(n407), .ZN(n364) );
  XOR2_X1 U496 ( .A(n655), .B(n654), .Z(n365) );
  AND2_X1 U497 ( .A1(KEYINPUT72), .A2(KEYINPUT44), .ZN(n366) );
  XNOR2_X2 U498 ( .A(n367), .B(n480), .ZN(n613) );
  XNOR2_X1 U499 ( .A(n790), .B(n368), .ZN(n705) );
  XNOR2_X1 U500 ( .A(n478), .B(n496), .ZN(n368) );
  XNOR2_X1 U501 ( .A(n497), .B(n358), .ZN(n790) );
  NAND2_X1 U502 ( .A1(n792), .A2(G234), .ZN(n391) );
  NAND2_X1 U503 ( .A1(n792), .A2(G224), .ZN(n514) );
  XNOR2_X2 U504 ( .A(n476), .B(G953), .ZN(n792) );
  XNOR2_X1 U505 ( .A(n454), .B(n482), .ZN(n788) );
  XNOR2_X1 U506 ( .A(n788), .B(n440), .ZN(n439) );
  NAND2_X1 U507 ( .A1(n382), .A2(n381), .ZN(n373) );
  NAND2_X1 U508 ( .A1(n382), .A2(n381), .ZN(n380) );
  INV_X1 U509 ( .A(n394), .ZN(n619) );
  AND2_X1 U510 ( .A1(n791), .A2(KEYINPUT66), .ZN(n383) );
  BUF_X1 U511 ( .A(n718), .Z(n374) );
  NAND2_X1 U512 ( .A1(n384), .A2(n383), .ZN(n381) );
  XNOR2_X1 U513 ( .A(n424), .B(KEYINPUT48), .ZN(n421) );
  INV_X2 U514 ( .A(n423), .ZN(n791) );
  NAND2_X1 U515 ( .A1(n423), .A2(n422), .ZN(n459) );
  NOR2_X1 U516 ( .A1(n718), .A2(n364), .ZN(n376) );
  NAND2_X1 U517 ( .A1(n652), .A2(n461), .ZN(n460) );
  OR2_X1 U518 ( .A1(n718), .A2(n364), .ZN(n377) );
  AND2_X2 U519 ( .A1(n380), .A2(n385), .ZN(n378) );
  AND2_X1 U520 ( .A1(n373), .A2(n385), .ZN(n709) );
  BUF_X1 U521 ( .A(n414), .Z(n394) );
  AND2_X2 U522 ( .A1(n379), .A2(n361), .ZN(n382) );
  NAND2_X1 U523 ( .A1(n375), .A2(n404), .ZN(n379) );
  NAND2_X1 U524 ( .A1(n375), .A2(n377), .ZN(n384) );
  NOR2_X1 U525 ( .A1(n374), .A2(n387), .ZN(n386) );
  NOR2_X1 U526 ( .A1(n388), .A2(n362), .ZN(n426) );
  INV_X1 U527 ( .A(n467), .ZN(n388) );
  NAND2_X1 U528 ( .A1(n389), .A2(n433), .ZN(n567) );
  NOR2_X1 U529 ( .A1(n417), .A2(n416), .ZN(n389) );
  NAND2_X1 U530 ( .A1(n426), .A2(n463), .ZN(n408) );
  NAND2_X1 U531 ( .A1(n414), .A2(n359), .ZN(n531) );
  XNOR2_X1 U532 ( .A(n392), .B(n430), .ZN(n429) );
  NAND2_X1 U533 ( .A1(n591), .A2(n592), .ZN(n392) );
  XNOR2_X1 U534 ( .A(n684), .B(n393), .ZN(n710) );
  XNOR2_X1 U535 ( .A(n517), .B(n518), .ZN(n393) );
  XNOR2_X1 U536 ( .A(n397), .B(n454), .ZN(n516) );
  INV_X1 U537 ( .A(n418), .ZN(n399) );
  NAND2_X1 U538 ( .A1(n418), .A2(n402), .ZN(n401) );
  XNOR2_X2 U539 ( .A(n577), .B(n456), .ZN(n418) );
  NAND2_X1 U540 ( .A1(n718), .A2(n407), .ZN(n406) );
  NAND2_X1 U541 ( .A1(n408), .A2(KEYINPUT91), .ZN(n411) );
  NAND2_X1 U542 ( .A1(n426), .A2(n410), .ZN(n409) );
  XNOR2_X1 U543 ( .A(n415), .B(G119), .ZN(G21) );
  XNOR2_X2 U544 ( .A(n585), .B(n584), .ZN(n415) );
  NAND2_X1 U545 ( .A1(n589), .A2(n418), .ZN(n590) );
  XNOR2_X1 U546 ( .A(n418), .B(G122), .ZN(G24) );
  NAND2_X1 U547 ( .A1(n578), .A2(n419), .ZN(n569) );
  XNOR2_X2 U548 ( .A(n613), .B(n481), .ZN(n737) );
  NAND2_X1 U549 ( .A1(n420), .A2(n799), .ZN(n617) );
  XNOR2_X1 U550 ( .A(n420), .B(G131), .ZN(G33) );
  NAND2_X1 U551 ( .A1(n355), .A2(n425), .ZN(n602) );
  NOR2_X2 U552 ( .A1(n738), .A2(n613), .ZN(n599) );
  XNOR2_X2 U553 ( .A(n427), .B(n363), .ZN(n718) );
  NAND2_X1 U554 ( .A1(n429), .A2(n428), .ZN(n427) );
  INV_X1 U555 ( .A(KEYINPUT90), .ZN(n430) );
  XNOR2_X1 U556 ( .A(n562), .B(n533), .ZN(n455) );
  XNOR2_X1 U557 ( .A(n431), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U558 ( .A1(n432), .A2(n657), .ZN(n431) );
  XNOR2_X1 U559 ( .A(n656), .B(n365), .ZN(n432) );
  NOR2_X1 U560 ( .A1(n669), .A2(n559), .ZN(n434) );
  INV_X1 U561 ( .A(n659), .ZN(n435) );
  NAND2_X1 U562 ( .A1(n442), .A2(n441), .ZN(n449) );
  INV_X1 U563 ( .A(n737), .ZN(n441) );
  NAND2_X1 U564 ( .A1(n447), .A2(n445), .ZN(n745) );
  NAND2_X1 U565 ( .A1(n737), .A2(n450), .ZN(n448) );
  INV_X1 U566 ( .A(n732), .ZN(n451) );
  XNOR2_X2 U567 ( .A(G146), .B(G125), .ZN(n454) );
  NAND2_X1 U568 ( .A1(n455), .A2(n766), .ZN(n571) );
  INV_X1 U569 ( .A(n652), .ZN(n458) );
  INV_X1 U570 ( .A(KEYINPUT66), .ZN(n461) );
  NAND2_X1 U571 ( .A1(n360), .A2(n467), .ZN(n603) );
  NAND2_X1 U572 ( .A1(n710), .A2(n521), .ZN(n467) );
  INV_X1 U573 ( .A(n749), .ZN(n468) );
  XOR2_X1 U574 ( .A(n485), .B(n484), .Z(n469) );
  AND2_X1 U575 ( .A1(n599), .A2(n610), .ZN(n470) );
  AND2_X1 U576 ( .A1(n565), .A2(n395), .ZN(n471) );
  XNOR2_X1 U577 ( .A(n492), .B(n491), .ZN(n564) );
  INV_X1 U578 ( .A(n715), .ZN(n657) );
  XNOR2_X1 U579 ( .A(n473), .B(G101), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n515), .B(G146), .ZN(n496) );
  NAND2_X1 U581 ( .A1(n792), .A2(G227), .ZN(n477) );
  XNOR2_X1 U582 ( .A(n354), .B(n477), .ZN(n478) );
  XNOR2_X1 U583 ( .A(KEYINPUT74), .B(G469), .ZN(n479) );
  XNOR2_X1 U584 ( .A(n479), .B(KEYINPUT73), .ZN(n480) );
  XNOR2_X1 U585 ( .A(KEYINPUT68), .B(KEYINPUT1), .ZN(n481) );
  XOR2_X1 U586 ( .A(KEYINPUT24), .B(KEYINPUT76), .Z(n485) );
  NAND2_X1 U587 ( .A1(n693), .A2(n555), .ZN(n492) );
  NAND2_X1 U588 ( .A1(n594), .A2(G234), .ZN(n488) );
  XNOR2_X1 U589 ( .A(n488), .B(KEYINPUT20), .ZN(n489) );
  XNOR2_X1 U590 ( .A(KEYINPUT96), .B(n489), .ZN(n493) );
  NAND2_X1 U591 ( .A1(G217), .A2(n493), .ZN(n490) );
  XNOR2_X1 U592 ( .A(KEYINPUT25), .B(n490), .ZN(n491) );
  AND2_X1 U593 ( .A1(n493), .A2(G221), .ZN(n495) );
  INV_X1 U594 ( .A(KEYINPUT21), .ZN(n494) );
  XNOR2_X1 U595 ( .A(n495), .B(n494), .ZN(n730) );
  XNOR2_X1 U596 ( .A(n497), .B(n496), .ZN(n504) );
  NAND2_X1 U597 ( .A1(n551), .A2(G210), .ZN(n498) );
  XNOR2_X1 U598 ( .A(n498), .B(G137), .ZN(n500) );
  XNOR2_X1 U599 ( .A(n500), .B(n499), .ZN(n502) );
  XNOR2_X1 U600 ( .A(n502), .B(n510), .ZN(n503) );
  XNOR2_X1 U601 ( .A(n504), .B(n503), .ZN(n655) );
  INV_X1 U602 ( .A(G472), .ZN(n505) );
  XNOR2_X2 U603 ( .A(n506), .B(n505), .ZN(n610) );
  INV_X1 U604 ( .A(n610), .ZN(n732) );
  XNOR2_X1 U605 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U606 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n512) );
  XNOR2_X1 U607 ( .A(KEYINPUT83), .B(KEYINPUT4), .ZN(n511) );
  XNOR2_X1 U608 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U609 ( .A(n514), .B(n513), .ZN(n518) );
  XNOR2_X1 U610 ( .A(n515), .B(n516), .ZN(n517) );
  INV_X1 U611 ( .A(n594), .ZN(n651) );
  XNOR2_X1 U612 ( .A(n519), .B(KEYINPUT80), .ZN(n523) );
  INV_X1 U613 ( .A(G214), .ZN(n522) );
  OR2_X1 U614 ( .A1(n523), .A2(n522), .ZN(n749) );
  XOR2_X1 U615 ( .A(KEYINPUT79), .B(KEYINPUT14), .Z(n525) );
  XNOR2_X1 U616 ( .A(n525), .B(n524), .ZN(n527) );
  NAND2_X1 U617 ( .A1(n527), .A2(G952), .ZN(n526) );
  XOR2_X1 U618 ( .A(KEYINPUT93), .B(n526), .Z(n764) );
  NOR2_X1 U619 ( .A1(n764), .A2(G953), .ZN(n598) );
  NAND2_X1 U620 ( .A1(G902), .A2(n527), .ZN(n595) );
  OR2_X1 U621 ( .A1(G898), .A2(n768), .ZN(n528) );
  XNOR2_X1 U622 ( .A(KEYINPUT94), .B(n528), .ZN(n687) );
  NOR2_X1 U623 ( .A1(n595), .A2(n687), .ZN(n529) );
  XNOR2_X2 U624 ( .A(n531), .B(n530), .ZN(n562) );
  NAND2_X1 U625 ( .A1(n562), .A2(n745), .ZN(n532) );
  NAND2_X1 U626 ( .A1(G217), .A2(n534), .ZN(n536) );
  XNOR2_X1 U627 ( .A(n535), .B(n536), .ZN(n543) );
  XNOR2_X1 U628 ( .A(n537), .B(KEYINPUT7), .ZN(n541) );
  XOR2_X1 U629 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n539) );
  XNOR2_X1 U630 ( .A(G122), .B(KEYINPUT9), .ZN(n538) );
  XNOR2_X1 U631 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U632 ( .A(n541), .B(n540), .Z(n542) );
  XNOR2_X1 U633 ( .A(n543), .B(n542), .ZN(n675) );
  NAND2_X1 U634 ( .A1(n675), .A2(n555), .ZN(n544) );
  XNOR2_X1 U635 ( .A(n544), .B(G478), .ZN(n572) );
  XNOR2_X1 U636 ( .A(n546), .B(n545), .ZN(n550) );
  XNOR2_X1 U637 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U638 ( .A(n550), .B(n549), .Z(n554) );
  NAND2_X1 U639 ( .A1(n551), .A2(G214), .ZN(n552) );
  XNOR2_X1 U640 ( .A(n788), .B(n552), .ZN(n553) );
  XNOR2_X1 U641 ( .A(n554), .B(n553), .ZN(n698) );
  NAND2_X1 U642 ( .A1(n698), .A2(n555), .ZN(n557) );
  XOR2_X1 U643 ( .A(KEYINPUT13), .B(G475), .Z(n556) );
  XNOR2_X1 U644 ( .A(n557), .B(n556), .ZN(n560) );
  INV_X1 U645 ( .A(n560), .ZN(n573) );
  AND2_X1 U646 ( .A1(n572), .A2(n573), .ZN(n775) );
  OR2_X1 U647 ( .A1(n781), .A2(n775), .ZN(n621) );
  INV_X1 U648 ( .A(n621), .ZN(n754) );
  INV_X1 U649 ( .A(KEYINPUT102), .ZN(n559) );
  OR2_X1 U650 ( .A1(n572), .A2(n560), .ZN(n752) );
  NOR2_X1 U651 ( .A1(n752), .A2(n730), .ZN(n561) );
  NAND2_X1 U652 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U653 ( .A1(n578), .A2(n729), .ZN(n565) );
  NAND2_X1 U654 ( .A1(n567), .A2(n672), .ZN(n568) );
  XNOR2_X1 U655 ( .A(n568), .B(KEYINPUT105), .ZN(n592) );
  XNOR2_X1 U656 ( .A(n569), .B(KEYINPUT33), .ZN(n766) );
  INV_X1 U657 ( .A(KEYINPUT34), .ZN(n570) );
  XNOR2_X1 U658 ( .A(n571), .B(n570), .ZN(n576) );
  INV_X1 U659 ( .A(n572), .ZN(n574) );
  OR2_X1 U660 ( .A1(n574), .A2(n573), .ZN(n625) );
  XOR2_X1 U661 ( .A(KEYINPUT84), .B(n625), .Z(n575) );
  NAND2_X1 U662 ( .A1(n576), .A2(n575), .ZN(n577) );
  INV_X1 U663 ( .A(n737), .ZN(n736) );
  NAND2_X1 U664 ( .A1(n736), .A2(n729), .ZN(n580) );
  INV_X1 U665 ( .A(KEYINPUT85), .ZN(n581) );
  INV_X1 U666 ( .A(KEYINPUT67), .ZN(n583) );
  XNOR2_X1 U667 ( .A(n583), .B(KEYINPUT32), .ZN(n584) );
  NAND2_X1 U668 ( .A1(n729), .A2(n610), .ZN(n586) );
  OR2_X1 U669 ( .A1(n586), .A2(n736), .ZN(n587) );
  OR2_X1 U670 ( .A1(n588), .A2(n587), .ZN(n658) );
  INV_X1 U671 ( .A(n593), .ZN(n589) );
  NAND2_X1 U672 ( .A1(n590), .A2(KEYINPUT44), .ZN(n591) );
  OR2_X1 U673 ( .A1(n595), .A2(n396), .ZN(n596) );
  NOR2_X1 U674 ( .A1(G900), .A2(n596), .ZN(n597) );
  NOR2_X1 U675 ( .A1(n598), .A2(n597), .ZN(n609) );
  NAND2_X1 U676 ( .A1(n732), .A2(n749), .ZN(n600) );
  XNOR2_X1 U677 ( .A(n600), .B(KEYINPUT30), .ZN(n601) );
  XOR2_X1 U678 ( .A(KEYINPUT38), .B(n603), .Z(n607) );
  XNOR2_X1 U679 ( .A(KEYINPUT39), .B(KEYINPUT77), .ZN(n604) );
  XNOR2_X1 U680 ( .A(n605), .B(n604), .ZN(n641) );
  NAND2_X1 U681 ( .A1(n641), .A2(n781), .ZN(n606) );
  INV_X1 U682 ( .A(n607), .ZN(n750) );
  NAND2_X1 U683 ( .A1(n750), .A2(n749), .ZN(n753) );
  NOR2_X1 U684 ( .A1(n752), .A2(n753), .ZN(n608) );
  XOR2_X1 U685 ( .A(KEYINPUT41), .B(n608), .Z(n767) );
  NOR2_X1 U686 ( .A1(n730), .A2(n609), .ZN(n642) );
  NAND2_X1 U687 ( .A1(n729), .A2(n642), .ZN(n611) );
  NOR2_X1 U688 ( .A1(n611), .A2(n610), .ZN(n612) );
  XOR2_X1 U689 ( .A(KEYINPUT28), .B(n612), .Z(n614) );
  NOR2_X1 U690 ( .A1(n614), .A2(n613), .ZN(n618) );
  NAND2_X1 U691 ( .A1(n767), .A2(n618), .ZN(n615) );
  XNOR2_X1 U692 ( .A(n615), .B(KEYINPUT42), .ZN(n799) );
  XOR2_X1 U693 ( .A(KEYINPUT46), .B(KEYINPUT89), .Z(n616) );
  XNOR2_X1 U694 ( .A(n617), .B(n616), .ZN(n640) );
  INV_X1 U695 ( .A(KEYINPUT78), .ZN(n624) );
  NOR2_X1 U696 ( .A1(n624), .A2(KEYINPUT47), .ZN(n623) );
  INV_X1 U697 ( .A(n618), .ZN(n620) );
  NOR2_X1 U698 ( .A1(n620), .A2(n619), .ZN(n782) );
  NAND2_X1 U699 ( .A1(n782), .A2(n621), .ZN(n622) );
  XNOR2_X1 U700 ( .A(n623), .B(n622), .ZN(n638) );
  NAND2_X1 U701 ( .A1(n624), .A2(KEYINPUT47), .ZN(n636) );
  OR2_X1 U702 ( .A1(n625), .A2(n603), .ZN(n626) );
  NOR2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n780) );
  NAND2_X1 U704 ( .A1(n781), .A2(n729), .ZN(n644) );
  INV_X1 U705 ( .A(n642), .ZN(n628) );
  NOR2_X1 U706 ( .A1(n644), .A2(n628), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n630), .A2(n629), .ZN(n631) );
  OR2_X1 U708 ( .A1(n631), .A2(n645), .ZN(n633) );
  INV_X1 U709 ( .A(KEYINPUT36), .ZN(n632) );
  XNOR2_X1 U710 ( .A(n633), .B(n632), .ZN(n634) );
  AND2_X1 U711 ( .A1(n634), .A2(n736), .ZN(n785) );
  NOR2_X1 U712 ( .A1(n780), .A2(n785), .ZN(n635) );
  AND2_X1 U713 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U715 ( .A1(n641), .A2(n775), .ZN(n787) );
  NAND2_X1 U716 ( .A1(n642), .A2(n749), .ZN(n643) );
  OR2_X1 U717 ( .A1(n644), .A2(n643), .ZN(n646) );
  NOR2_X1 U718 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U719 ( .A1(n647), .A2(n395), .ZN(n648) );
  XNOR2_X1 U720 ( .A(n648), .B(KEYINPUT43), .ZN(n649) );
  NAND2_X1 U721 ( .A1(n649), .A2(n603), .ZN(n674) );
  AND2_X1 U722 ( .A1(n787), .A2(n674), .ZN(n650) );
  NAND2_X1 U723 ( .A1(n651), .A2(KEYINPUT2), .ZN(n652) );
  NAND2_X1 U724 ( .A1(n709), .A2(G472), .ZN(n656) );
  XOR2_X1 U725 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n653) );
  XNOR2_X1 U726 ( .A(n653), .B(KEYINPUT62), .ZN(n654) );
  XNOR2_X1 U727 ( .A(n658), .B(G110), .ZN(G12) );
  NAND2_X1 U728 ( .A1(n662), .A2(n775), .ZN(n661) );
  XOR2_X1 U729 ( .A(G116), .B(KEYINPUT115), .Z(n660) );
  XNOR2_X1 U730 ( .A(n661), .B(n660), .ZN(G18) );
  NAND2_X1 U731 ( .A1(n662), .A2(n781), .ZN(n663) );
  XNOR2_X1 U732 ( .A(n663), .B(G113), .ZN(G15) );
  NAND2_X1 U733 ( .A1(n669), .A2(n775), .ZN(n668) );
  XOR2_X1 U734 ( .A(KEYINPUT27), .B(KEYINPUT111), .Z(n665) );
  XNOR2_X1 U735 ( .A(G107), .B(KEYINPUT110), .ZN(n664) );
  XNOR2_X1 U736 ( .A(n665), .B(n664), .ZN(n666) );
  XOR2_X1 U737 ( .A(KEYINPUT26), .B(n666), .Z(n667) );
  XNOR2_X1 U738 ( .A(n668), .B(n667), .ZN(G9) );
  NAND2_X1 U739 ( .A1(n669), .A2(n781), .ZN(n671) );
  XOR2_X1 U740 ( .A(G104), .B(KEYINPUT109), .Z(n670) );
  XNOR2_X1 U741 ( .A(n671), .B(n670), .ZN(G6) );
  XNOR2_X1 U742 ( .A(n672), .B(G101), .ZN(G3) );
  XNOR2_X1 U743 ( .A(G140), .B(KEYINPUT116), .ZN(n673) );
  XNOR2_X1 U744 ( .A(n674), .B(n673), .ZN(G42) );
  NAND2_X1 U745 ( .A1(n378), .A2(G478), .ZN(n677) );
  INV_X1 U746 ( .A(n675), .ZN(n676) );
  XNOR2_X1 U747 ( .A(n677), .B(n676), .ZN(n678) );
  NOR2_X2 U748 ( .A1(n678), .A2(n715), .ZN(n679) );
  XNOR2_X1 U749 ( .A(n679), .B(KEYINPUT122), .ZN(G63) );
  INV_X1 U750 ( .A(n374), .ZN(n724) );
  NAND2_X1 U751 ( .A1(n724), .A2(n768), .ZN(n683) );
  NAND2_X1 U752 ( .A1(G953), .A2(G224), .ZN(n680) );
  XNOR2_X1 U753 ( .A(KEYINPUT61), .B(n680), .ZN(n681) );
  NAND2_X1 U754 ( .A1(n681), .A2(G898), .ZN(n682) );
  NAND2_X1 U755 ( .A1(n683), .A2(n682), .ZN(n692) );
  BUF_X1 U756 ( .A(n684), .Z(n685) );
  XOR2_X1 U757 ( .A(G101), .B(KEYINPUT124), .Z(n686) );
  XNOR2_X1 U758 ( .A(n685), .B(n686), .ZN(n688) );
  NAND2_X1 U759 ( .A1(n688), .A2(n687), .ZN(n690) );
  XNOR2_X1 U760 ( .A(KEYINPUT125), .B(KEYINPUT126), .ZN(n689) );
  XNOR2_X1 U761 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U762 ( .A(n692), .B(n691), .ZN(G69) );
  NAND2_X1 U763 ( .A1(n709), .A2(G217), .ZN(n695) );
  XNOR2_X1 U764 ( .A(n693), .B(KEYINPUT123), .ZN(n694) );
  XNOR2_X1 U765 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X1 U766 ( .A1(n696), .A2(n715), .ZN(G66) );
  NAND2_X1 U767 ( .A1(n378), .A2(G475), .ZN(n700) );
  XOR2_X1 U768 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n697) );
  XNOR2_X1 U769 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U770 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X2 U771 ( .A1(n701), .A2(n715), .ZN(n702) );
  XNOR2_X1 U772 ( .A(n702), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U773 ( .A1(n709), .A2(G469), .ZN(n707) );
  XOR2_X1 U774 ( .A(KEYINPUT120), .B(KEYINPUT57), .Z(n703) );
  XNOR2_X1 U775 ( .A(n703), .B(KEYINPUT58), .ZN(n704) );
  XNOR2_X1 U776 ( .A(n705), .B(n704), .ZN(n706) );
  XNOR2_X1 U777 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U778 ( .A1(n708), .A2(n715), .ZN(G54) );
  NAND2_X1 U779 ( .A1(n378), .A2(G210), .ZN(n714) );
  BUF_X1 U780 ( .A(n710), .Z(n712) );
  XOR2_X1 U781 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n711) );
  XNOR2_X1 U782 ( .A(n712), .B(n711), .ZN(n713) );
  XNOR2_X1 U783 ( .A(n714), .B(n713), .ZN(n716) );
  NOR2_X2 U784 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U785 ( .A(n717), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X1 U786 ( .A1(n374), .A2(n423), .ZN(n719) );
  NOR2_X1 U787 ( .A1(n719), .A2(KEYINPUT2), .ZN(n720) );
  NOR2_X1 U788 ( .A1(n720), .A2(KEYINPUT87), .ZN(n726) );
  INV_X1 U789 ( .A(KEYINPUT87), .ZN(n721) );
  NOR2_X1 U790 ( .A1(n721), .A2(KEYINPUT2), .ZN(n722) );
  NAND2_X1 U791 ( .A1(n791), .A2(n722), .ZN(n723) );
  NOR2_X1 U792 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U793 ( .A1(n726), .A2(n725), .ZN(n728) );
  OR2_X1 U794 ( .A1(n728), .A2(n727), .ZN(n773) );
  NAND2_X1 U795 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U796 ( .A(n731), .B(KEYINPUT49), .ZN(n733) );
  OR2_X1 U797 ( .A1(n733), .A2(n732), .ZN(n743) );
  INV_X1 U798 ( .A(KEYINPUT50), .ZN(n734) );
  NAND2_X1 U799 ( .A1(n738), .A2(n734), .ZN(n735) );
  NOR2_X1 U800 ( .A1(n736), .A2(n735), .ZN(n741) );
  NAND2_X1 U801 ( .A1(n738), .A2(n395), .ZN(n739) );
  AND2_X1 U802 ( .A1(n739), .A2(KEYINPUT50), .ZN(n740) );
  NOR2_X1 U803 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U804 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U805 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U806 ( .A(KEYINPUT117), .B(n746), .Z(n747) );
  XNOR2_X1 U807 ( .A(KEYINPUT51), .B(n747), .ZN(n748) );
  NAND2_X1 U808 ( .A1(n748), .A2(n767), .ZN(n761) );
  NOR2_X1 U809 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U810 ( .A1(n752), .A2(n751), .ZN(n756) );
  NOR2_X1 U811 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U812 ( .A1(n756), .A2(n755), .ZN(n758) );
  INV_X1 U813 ( .A(n766), .ZN(n757) );
  NOR2_X1 U814 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U815 ( .A(KEYINPUT118), .B(n759), .Z(n760) );
  NAND2_X1 U816 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U817 ( .A(KEYINPUT52), .B(n762), .Z(n763) );
  NOR2_X1 U818 ( .A1(n764), .A2(n763), .ZN(n765) );
  XOR2_X1 U819 ( .A(KEYINPUT119), .B(n765), .Z(n771) );
  NAND2_X1 U820 ( .A1(n767), .A2(n766), .ZN(n769) );
  NAND2_X1 U821 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X1 U822 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U823 ( .A1(n773), .A2(n772), .ZN(n774) );
  XOR2_X1 U824 ( .A(KEYINPUT53), .B(n774), .Z(G75) );
  XOR2_X1 U825 ( .A(KEYINPUT29), .B(KEYINPUT113), .Z(n777) );
  NAND2_X1 U826 ( .A1(n782), .A2(n775), .ZN(n776) );
  XNOR2_X1 U827 ( .A(n777), .B(n776), .ZN(n779) );
  XOR2_X1 U828 ( .A(G128), .B(KEYINPUT112), .Z(n778) );
  XNOR2_X1 U829 ( .A(n779), .B(n778), .ZN(G30) );
  XOR2_X1 U830 ( .A(G143), .B(n780), .Z(G45) );
  NAND2_X1 U831 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U832 ( .A(n783), .B(KEYINPUT114), .ZN(n784) );
  XNOR2_X1 U833 ( .A(G146), .B(n784), .ZN(G48) );
  XNOR2_X1 U834 ( .A(n785), .B(G125), .ZN(n786) );
  XNOR2_X1 U835 ( .A(n786), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U836 ( .A(G134), .B(n787), .ZN(G36) );
  XNOR2_X1 U837 ( .A(n788), .B(KEYINPUT127), .ZN(n789) );
  XNOR2_X1 U838 ( .A(n790), .B(n789), .ZN(n794) );
  XOR2_X1 U839 ( .A(n794), .B(n791), .Z(n793) );
  NAND2_X1 U840 ( .A1(n793), .A2(n396), .ZN(n798) );
  XNOR2_X1 U841 ( .A(G227), .B(n794), .ZN(n795) );
  NAND2_X1 U842 ( .A1(n795), .A2(G900), .ZN(n796) );
  NAND2_X1 U843 ( .A1(n796), .A2(G953), .ZN(n797) );
  NAND2_X1 U844 ( .A1(n798), .A2(n797), .ZN(G72) );
  XNOR2_X1 U845 ( .A(G137), .B(n799), .ZN(G39) );
endmodule

