

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816;

  AND2_X1 U377 ( .A1(n373), .A2(n623), .ZN(n355) );
  AND2_X1 U378 ( .A1(n695), .A2(n410), .ZN(n356) );
  AND2_X1 U379 ( .A1(n485), .A2(n745), .ZN(n739) );
  NAND2_X1 U380 ( .A1(n399), .A2(n397), .ZN(n396) );
  XNOR2_X1 U381 ( .A(n363), .B(n362), .ZN(n693) );
  NOR2_X2 U382 ( .A1(n461), .A2(n460), .ZN(n423) );
  XNOR2_X1 U383 ( .A(n621), .B(KEYINPUT86), .ZN(n624) );
  XNOR2_X2 U384 ( .A(n640), .B(KEYINPUT41), .ZN(n773) );
  INV_X1 U385 ( .A(n665), .ZN(n667) );
  XNOR2_X1 U386 ( .A(n511), .B(n583), .ZN(n802) );
  NOR2_X2 U387 ( .A1(G953), .A2(G237), .ZN(n591) );
  AND2_X1 U388 ( .A1(n381), .A2(KEYINPUT56), .ZN(n380) );
  AND2_X1 U389 ( .A1(n695), .A2(n358), .ZN(n360) );
  XNOR2_X1 U390 ( .A(n617), .B(n616), .ZN(n702) );
  XNOR2_X1 U391 ( .A(n620), .B(KEYINPUT32), .ZN(n456) );
  INV_X1 U392 ( .A(n644), .ZN(n744) );
  NOR2_X1 U393 ( .A1(n667), .A2(n666), .ZN(n669) );
  OR2_X1 U394 ( .A1(n708), .A2(G902), .ZN(n488) );
  XNOR2_X1 U395 ( .A(n490), .B(n489), .ZN(n797) );
  XNOR2_X1 U396 ( .A(n500), .B(n574), .ZN(n490) );
  XNOR2_X1 U397 ( .A(n802), .B(n512), .ZN(n530) );
  XNOR2_X1 U398 ( .A(n531), .B(n501), .ZN(n500) );
  XNOR2_X1 U399 ( .A(n474), .B(G146), .ZN(n544) );
  INV_X1 U400 ( .A(G125), .ZN(n474) );
  INV_X1 U401 ( .A(KEYINPUT74), .ZN(n513) );
  BUF_X1 U402 ( .A(G128), .Z(n471) );
  XNOR2_X1 U403 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n516) );
  XNOR2_X1 U404 ( .A(G119), .B(KEYINPUT3), .ZN(n515) );
  INV_X1 U405 ( .A(KEYINPUT45), .ZN(n362) );
  NAND2_X1 U406 ( .A1(n382), .A2(n380), .ZN(n379) );
  INV_X1 U407 ( .A(n396), .ZN(n395) );
  INV_X1 U408 ( .A(n388), .ZN(n382) );
  INV_X1 U409 ( .A(n412), .ZN(n357) );
  AND2_X1 U410 ( .A1(n438), .A2(KEYINPUT78), .ZN(n435) );
  AND2_X1 U411 ( .A1(n367), .A2(n355), .ZN(n365) );
  NAND2_X1 U412 ( .A1(n420), .A2(n419), .ZN(n438) );
  XNOR2_X1 U413 ( .A(n377), .B(n494), .ZN(n372) );
  OR2_X1 U414 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U415 ( .A(n366), .B(KEYINPUT72), .ZN(n364) );
  NAND2_X1 U416 ( .A1(n726), .A2(n456), .ZN(n621) );
  NOR2_X1 U417 ( .A1(n409), .A2(KEYINPUT56), .ZN(n385) );
  XNOR2_X1 U418 ( .A(n607), .B(KEYINPUT106), .ZN(n761) );
  OR2_X1 U419 ( .A1(n626), .A2(n565), .ZN(n644) );
  XNOR2_X1 U420 ( .A(n561), .B(n560), .ZN(n626) );
  AND2_X1 U421 ( .A1(n390), .A2(n709), .ZN(n389) );
  AND2_X1 U422 ( .A1(n398), .A2(n709), .ZN(n397) );
  AND2_X1 U423 ( .A1(n409), .A2(n498), .ZN(n392) );
  INV_X1 U424 ( .A(n409), .ZN(n387) );
  INV_X1 U425 ( .A(n706), .ZN(n394) );
  OR2_X1 U426 ( .A1(n706), .A2(n496), .ZN(n398) );
  XNOR2_X1 U427 ( .A(n544), .B(KEYINPUT10), .ZN(n547) );
  XNOR2_X1 U428 ( .A(n426), .B(n425), .ZN(n586) );
  INV_X1 U429 ( .A(n515), .ZN(n517) );
  NOR2_X1 U430 ( .A1(n696), .A2(n427), .ZN(n410) );
  NOR2_X1 U431 ( .A1(n696), .A2(n604), .ZN(n415) );
  INV_X2 U432 ( .A(G953), .ZN(n806) );
  XNOR2_X1 U433 ( .A(KEYINPUT7), .B(G122), .ZN(n582) );
  XNOR2_X1 U434 ( .A(KEYINPUT67), .B(KEYINPUT4), .ZN(n511) );
  XNOR2_X1 U435 ( .A(G122), .B(G104), .ZN(n514) );
  XNOR2_X1 U436 ( .A(G107), .B(G104), .ZN(n533) );
  INV_X1 U437 ( .A(n696), .ZN(n358) );
  NAND2_X1 U438 ( .A1(n359), .A2(n466), .ZN(n465) );
  NOR2_X1 U439 ( .A1(n359), .A2(n493), .ZN(n460) );
  NAND2_X1 U440 ( .A1(n774), .A2(n359), .ZN(n477) );
  XNOR2_X2 U441 ( .A(n378), .B(n455), .ZN(n359) );
  AND2_X2 U442 ( .A1(n467), .A2(n695), .ZN(n412) );
  AND2_X1 U443 ( .A1(n467), .A2(n356), .ZN(n470) );
  AND2_X1 U444 ( .A1(n467), .A2(n360), .ZN(n785) );
  AND2_X1 U445 ( .A1(n467), .A2(n361), .ZN(n413) );
  AND2_X1 U446 ( .A1(n695), .A2(n415), .ZN(n361) );
  NOR2_X1 U447 ( .A1(n412), .A2(n778), .ZN(n779) );
  NAND2_X1 U448 ( .A1(n365), .A2(n364), .ZN(n363) );
  NAND2_X1 U449 ( .A1(n368), .A2(n625), .ZN(n366) );
  NAND2_X1 U450 ( .A1(n369), .A2(n371), .ZN(n367) );
  XNOR2_X1 U451 ( .A(n624), .B(KEYINPUT85), .ZN(n368) );
  NAND2_X1 U452 ( .A1(n370), .A2(n618), .ZN(n369) );
  INV_X1 U453 ( .A(n372), .ZN(n370) );
  NAND2_X1 U454 ( .A1(n375), .A2(n372), .ZN(n371) );
  NAND2_X1 U455 ( .A1(n374), .A2(KEYINPUT84), .ZN(n373) );
  INV_X1 U456 ( .A(n376), .ZN(n374) );
  NAND2_X1 U457 ( .A1(n376), .A2(n618), .ZN(n375) );
  NAND2_X1 U458 ( .A1(n702), .A2(KEYINPUT44), .ZN(n376) );
  NAND2_X1 U459 ( .A1(n495), .A2(n718), .ZN(n377) );
  NAND2_X1 U460 ( .A1(n502), .A2(n378), .ZN(n503) );
  AND2_X1 U461 ( .A1(n454), .A2(n378), .ZN(n405) );
  XNOR2_X2 U462 ( .A(n528), .B(n408), .ZN(n378) );
  NAND2_X1 U463 ( .A1(n383), .A2(n379), .ZN(G51) );
  NAND2_X1 U464 ( .A1(n357), .A2(n387), .ZN(n381) );
  AND2_X1 U465 ( .A1(n386), .A2(n384), .ZN(n383) );
  NAND2_X1 U466 ( .A1(n357), .A2(n385), .ZN(n384) );
  NAND2_X1 U467 ( .A1(n388), .A2(n411), .ZN(n386) );
  NAND2_X1 U468 ( .A1(n391), .A2(n389), .ZN(n388) );
  OR2_X1 U469 ( .A1(n409), .A2(n498), .ZN(n390) );
  NAND2_X1 U470 ( .A1(n412), .A2(n392), .ZN(n391) );
  NAND2_X1 U471 ( .A1(n395), .A2(n393), .ZN(n401) );
  NAND2_X1 U472 ( .A1(n357), .A2(n394), .ZN(n393) );
  NAND2_X1 U473 ( .A1(n412), .A2(n400), .ZN(n399) );
  AND2_X1 U474 ( .A1(n706), .A2(n496), .ZN(n400) );
  XNOR2_X1 U475 ( .A(n401), .B(n707), .ZN(G57) );
  NOR2_X1 U476 ( .A1(n699), .A2(n789), .ZN(n701) );
  NOR2_X2 U477 ( .A1(n606), .A2(n614), .ZN(n668) );
  NOR2_X1 U478 ( .A1(n445), .A2(n444), .ZN(n443) );
  INV_X1 U479 ( .A(n547), .ZN(n601) );
  INV_X1 U480 ( .A(KEYINPUT113), .ZN(n434) );
  INV_X1 U481 ( .A(G902), .ZN(n577) );
  INV_X1 U482 ( .A(KEYINPUT93), .ZN(n455) );
  XNOR2_X1 U483 ( .A(KEYINPUT15), .B(G902), .ZN(n696) );
  INV_X1 U484 ( .A(KEYINPUT81), .ZN(n484) );
  INV_X1 U485 ( .A(KEYINPUT108), .ZN(n494) );
  INV_X1 U486 ( .A(n743), .ZN(n481) );
  INV_X1 U487 ( .A(KEYINPUT48), .ZN(n458) );
  AND2_X1 U488 ( .A1(n743), .A2(KEYINPUT79), .ZN(n482) );
  INV_X1 U489 ( .A(KEYINPUT8), .ZN(n425) );
  NAND2_X1 U490 ( .A1(n806), .A2(G234), .ZN(n426) );
  AND2_X1 U491 ( .A1(n433), .A2(n432), .ZN(n640) );
  INV_X1 U492 ( .A(n761), .ZN(n432) );
  INV_X1 U493 ( .A(KEYINPUT42), .ZN(n452) );
  OR2_X1 U494 ( .A1(n714), .A2(G902), .ZN(n540) );
  AND2_X1 U495 ( .A1(n463), .A2(n632), .ZN(n462) );
  NAND2_X1 U496 ( .A1(n464), .A2(KEYINPUT98), .ZN(n463) );
  XOR2_X1 U497 ( .A(G116), .B(G107), .Z(n581) );
  XNOR2_X1 U498 ( .A(n477), .B(n476), .ZN(n475) );
  INV_X1 U499 ( .A(KEYINPUT34), .ZN(n476) );
  XNOR2_X1 U500 ( .A(n603), .B(G475), .ZN(n487) );
  INV_X1 U501 ( .A(G210), .ZN(n499) );
  NAND2_X1 U502 ( .A1(n626), .A2(n468), .ZN(n666) );
  AND2_X1 U503 ( .A1(n749), .A2(n646), .ZN(n468) );
  OR2_X1 U504 ( .A1(G902), .A2(G237), .ZN(n519) );
  XNOR2_X1 U505 ( .A(G116), .B(G131), .ZN(n570) );
  INV_X1 U506 ( .A(KEYINPUT99), .ZN(n569) );
  XOR2_X1 U507 ( .A(G113), .B(KEYINPUT5), .Z(n568) );
  XNOR2_X1 U508 ( .A(G137), .B(G134), .ZN(n803) );
  INV_X1 U509 ( .A(G101), .ZN(n512) );
  AND2_X1 U510 ( .A1(n480), .A2(n741), .ZN(n479) );
  NAND2_X1 U511 ( .A1(n481), .A2(n419), .ZN(n480) );
  NAND2_X1 U512 ( .A1(G237), .A2(G234), .ZN(n522) );
  XNOR2_X1 U513 ( .A(n687), .B(n638), .ZN(n759) );
  INV_X1 U514 ( .A(KEYINPUT22), .ZN(n431) );
  INV_X1 U515 ( .A(KEYINPUT16), .ZN(n501) );
  XOR2_X1 U516 ( .A(KEYINPUT96), .B(G140), .Z(n552) );
  XNOR2_X1 U517 ( .A(G119), .B(G110), .ZN(n551) );
  XNOR2_X1 U518 ( .A(n547), .B(n546), .ZN(n550) );
  XNOR2_X1 U519 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n553) );
  XOR2_X1 U520 ( .A(KEYINPUT77), .B(KEYINPUT94), .Z(n554) );
  XNOR2_X1 U521 ( .A(n589), .B(n590), .ZN(n697) );
  XNOR2_X1 U522 ( .A(n602), .B(n805), .ZN(n708) );
  XNOR2_X1 U523 ( .A(G140), .B(G131), .ZN(n600) );
  INV_X1 U524 ( .A(KEYINPUT78), .ZN(n436) );
  INV_X1 U525 ( .A(KEYINPUT2), .ZN(n691) );
  XNOR2_X1 U526 ( .A(n612), .B(KEYINPUT33), .ZN(n774) );
  NAND2_X1 U527 ( .A1(n448), .A2(n447), .ZN(n418) );
  NOR2_X1 U528 ( .A1(n641), .A2(n452), .ZN(n447) );
  AND2_X1 U529 ( .A1(n451), .A2(n450), .ZN(n449) );
  NAND2_X1 U530 ( .A1(n641), .A2(n452), .ZN(n450) );
  XNOR2_X1 U531 ( .A(n428), .B(n427), .ZN(n606) );
  NOR2_X1 U532 ( .A1(n697), .A2(G902), .ZN(n428) );
  INV_X1 U533 ( .A(KEYINPUT100), .ZN(n422) );
  INV_X1 U534 ( .A(G472), .ZN(n497) );
  INV_X1 U535 ( .A(n697), .ZN(n469) );
  NAND2_X1 U536 ( .A1(n449), .A2(n418), .ZN(n816) );
  XNOR2_X1 U537 ( .A(KEYINPUT36), .B(KEYINPUT115), .ZN(n673) );
  NAND2_X1 U538 ( .A1(n475), .A2(n654), .ZN(n617) );
  INV_X1 U539 ( .A(n754), .ZN(n454) );
  XNOR2_X1 U540 ( .A(n668), .B(KEYINPUT110), .ZN(n719) );
  INV_X1 U541 ( .A(KEYINPUT56), .ZN(n411) );
  INV_X1 U542 ( .A(n745), .ZN(n429) );
  OR2_X1 U543 ( .A1(n763), .A2(n681), .ZN(n402) );
  AND2_X1 U544 ( .A1(n416), .A2(n429), .ZN(n403) );
  AND2_X1 U545 ( .A1(n457), .A2(n479), .ZN(n404) );
  NOR2_X1 U546 ( .A1(n750), .A2(n619), .ZN(n406) );
  AND2_X1 U547 ( .A1(n626), .A2(n632), .ZN(n407) );
  XOR2_X1 U548 ( .A(KEYINPUT66), .B(KEYINPUT0), .Z(n408) );
  INV_X1 U549 ( .A(KEYINPUT98), .ZN(n493) );
  XOR2_X1 U550 ( .A(n784), .B(n783), .Z(n409) );
  INV_X1 U551 ( .A(G478), .ZN(n427) );
  XNOR2_X1 U552 ( .A(n413), .B(n414), .ZN(n710) );
  XOR2_X1 U553 ( .A(n708), .B(KEYINPUT59), .Z(n414) );
  NAND2_X1 U554 ( .A1(n483), .A2(n482), .ZN(n457) );
  NAND2_X1 U555 ( .A1(n465), .A2(n462), .ZN(n461) );
  XNOR2_X1 U556 ( .A(n503), .B(n431), .ZN(n416) );
  XNOR2_X1 U557 ( .A(n503), .B(n431), .ZN(n430) );
  XNOR2_X1 U558 ( .A(n739), .B(n484), .ZN(n674) );
  NOR2_X1 U559 ( .A1(n761), .A2(n565), .ZN(n502) );
  NOR2_X1 U560 ( .A1(n653), .A2(n759), .ZN(n650) );
  BUF_X1 U561 ( .A(n637), .Z(n687) );
  NAND2_X1 U562 ( .A1(n430), .A2(n429), .ZN(n424) );
  BUF_X1 U563 ( .A(n722), .Z(n417) );
  XNOR2_X1 U564 ( .A(n423), .B(n422), .ZN(n722) );
  NAND2_X1 U565 ( .A1(n418), .A2(n652), .ZN(n444) );
  INV_X1 U566 ( .A(KEYINPUT79), .ZN(n419) );
  INV_X1 U567 ( .A(n483), .ZN(n420) );
  NAND2_X1 U568 ( .A1(n421), .A2(n605), .ZN(n495) );
  NAND2_X1 U569 ( .A1(n722), .A2(n736), .ZN(n421) );
  NAND2_X1 U570 ( .A1(n403), .A2(n667), .ZN(n609) );
  XNOR2_X1 U571 ( .A(n424), .B(KEYINPUT109), .ZN(n478) );
  NAND2_X1 U572 ( .A1(n586), .A2(G217), .ZN(n587) );
  NAND2_X1 U573 ( .A1(n416), .A2(n406), .ZN(n620) );
  AND2_X1 U574 ( .A1(n433), .A2(n605), .ZN(n764) );
  XNOR2_X1 U575 ( .A(n639), .B(n434), .ZN(n433) );
  NAND2_X1 U576 ( .A1(n404), .A2(n438), .ZN(n437) );
  NAND2_X1 U577 ( .A1(n404), .A2(n435), .ZN(n690) );
  AND2_X1 U578 ( .A1(n437), .A2(n436), .ZN(n694) );
  XNOR2_X1 U579 ( .A(n437), .B(n809), .ZN(n807) );
  NAND2_X1 U580 ( .A1(n439), .A2(n453), .ZN(n446) );
  NAND2_X1 U581 ( .A1(n441), .A2(n440), .ZN(n439) );
  INV_X1 U582 ( .A(n814), .ZN(n440) );
  INV_X1 U583 ( .A(n816), .ZN(n441) );
  NAND2_X1 U584 ( .A1(n446), .A2(n442), .ZN(n677) );
  NAND2_X1 U585 ( .A1(n440), .A2(n443), .ZN(n442) );
  INV_X1 U586 ( .A(n449), .ZN(n445) );
  INV_X1 U587 ( .A(n773), .ZN(n448) );
  NAND2_X1 U588 ( .A1(n773), .A2(n452), .ZN(n451) );
  INV_X1 U589 ( .A(n652), .ZN(n453) );
  XNOR2_X1 U590 ( .A(n456), .B(G119), .ZN(G21) );
  XNOR2_X2 U591 ( .A(n459), .B(n458), .ZN(n483) );
  NAND2_X1 U592 ( .A1(n677), .A2(n472), .ZN(n459) );
  NAND2_X1 U593 ( .A1(n667), .A2(n745), .ZN(n619) );
  XNOR2_X2 U594 ( .A(n647), .B(n579), .ZN(n745) );
  XNOR2_X2 U595 ( .A(n540), .B(n539), .ZN(n647) );
  INV_X1 U596 ( .A(n566), .ZN(n464) );
  AND2_X1 U597 ( .A1(n566), .A2(n493), .ZN(n466) );
  XNOR2_X2 U598 ( .A(n692), .B(n691), .ZN(n467) );
  NOR2_X1 U599 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U600 ( .A1(n676), .A2(n402), .ZN(n473) );
  XNOR2_X1 U601 ( .A(n550), .B(n549), .ZN(n558) );
  XNOR2_X1 U602 ( .A(n470), .B(n469), .ZN(n699) );
  INV_X1 U603 ( .A(n473), .ZN(n472) );
  NAND2_X1 U604 ( .A1(n478), .A2(n407), .ZN(n726) );
  XNOR2_X1 U605 ( .A(n486), .B(n673), .ZN(n485) );
  NAND2_X1 U606 ( .A1(n672), .A2(n671), .ZN(n486) );
  XNOR2_X2 U607 ( .A(n488), .B(n487), .ZN(n614) );
  XNOR2_X1 U608 ( .A(n598), .B(n581), .ZN(n489) );
  NOR2_X1 U609 ( .A1(n780), .A2(n358), .ZN(n518) );
  XNOR2_X1 U610 ( .A(n797), .B(n491), .ZN(n780) );
  XNOR2_X1 U611 ( .A(n530), .B(n492), .ZN(n491) );
  XNOR2_X1 U612 ( .A(n507), .B(n510), .ZN(n492) );
  NOR2_X1 U613 ( .A1(n696), .A2(n497), .ZN(n496) );
  NOR2_X1 U614 ( .A1(n696), .A2(n499), .ZN(n498) );
  XNOR2_X2 U615 ( .A(n517), .B(n516), .ZN(n574) );
  XNOR2_X1 U616 ( .A(n518), .B(n504), .ZN(n637) );
  AND2_X1 U617 ( .A1(G210), .A2(n519), .ZN(n504) );
  XOR2_X1 U618 ( .A(KEYINPUT82), .B(KEYINPUT39), .Z(n505) );
  XNOR2_X1 U619 ( .A(n570), .B(n569), .ZN(n571) );
  INV_X1 U620 ( .A(KEYINPUT30), .ZN(n642) );
  XNOR2_X1 U621 ( .A(n572), .B(n571), .ZN(n573) );
  INV_X1 U622 ( .A(KEYINPUT19), .ZN(n521) );
  XNOR2_X1 U623 ( .A(n545), .B(G137), .ZN(n546) );
  AND2_X1 U624 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U625 ( .A(n548), .B(n471), .ZN(n549) );
  BUF_X1 U626 ( .A(n780), .Z(n784) );
  XNOR2_X1 U627 ( .A(n650), .B(n505), .ZN(n689) );
  INV_X1 U628 ( .A(KEYINPUT123), .ZN(n700) );
  NAND2_X1 U629 ( .A1(G224), .A2(n806), .ZN(n506) );
  XNOR2_X1 U630 ( .A(n544), .B(n506), .ZN(n507) );
  XOR2_X1 U631 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n509) );
  XNOR2_X1 U632 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n508) );
  XNOR2_X1 U633 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X2 U634 ( .A(G143), .B(G128), .ZN(n583) );
  XNOR2_X2 U635 ( .A(n513), .B(G110), .ZN(n531) );
  XNOR2_X1 U636 ( .A(n514), .B(G113), .ZN(n598) );
  NAND2_X1 U637 ( .A1(n519), .A2(G214), .ZN(n520) );
  XNOR2_X1 U638 ( .A(KEYINPUT91), .B(n520), .ZN(n758) );
  NOR2_X2 U639 ( .A1(n637), .A2(n758), .ZN(n671) );
  XNOR2_X1 U640 ( .A(n671), .B(n521), .ZN(n658) );
  NOR2_X1 U641 ( .A1(G898), .A2(n806), .ZN(n799) );
  XNOR2_X1 U642 ( .A(n522), .B(KEYINPUT14), .ZN(n524) );
  NAND2_X1 U643 ( .A1(G902), .A2(n524), .ZN(n627) );
  INV_X1 U644 ( .A(n627), .ZN(n523) );
  NAND2_X1 U645 ( .A1(n799), .A2(n523), .ZN(n526) );
  NAND2_X1 U646 ( .A1(G952), .A2(n524), .ZN(n772) );
  NOR2_X1 U647 ( .A1(G953), .A2(n772), .ZN(n525) );
  XOR2_X1 U648 ( .A(KEYINPUT92), .B(n525), .Z(n631) );
  NAND2_X1 U649 ( .A1(n526), .A2(n631), .ZN(n527) );
  NAND2_X1 U650 ( .A1(n527), .A2(n658), .ZN(n528) );
  XNOR2_X1 U651 ( .A(n803), .B(G146), .ZN(n529) );
  XNOR2_X1 U652 ( .A(n530), .B(n529), .ZN(n576) );
  XNOR2_X1 U653 ( .A(n531), .B(n600), .ZN(n535) );
  NAND2_X1 U654 ( .A1(n806), .A2(G227), .ZN(n532) );
  XNOR2_X1 U655 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U656 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U657 ( .A(n576), .B(n536), .ZN(n714) );
  XNOR2_X1 U658 ( .A(KEYINPUT69), .B(G469), .ZN(n538) );
  INV_X1 U659 ( .A(KEYINPUT68), .ZN(n537) );
  XNOR2_X1 U660 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U661 ( .A(KEYINPUT97), .B(KEYINPUT25), .Z(n543) );
  NAND2_X1 U662 ( .A1(G234), .A2(n696), .ZN(n541) );
  XNOR2_X1 U663 ( .A(KEYINPUT20), .B(n541), .ZN(n562) );
  NAND2_X1 U664 ( .A1(n562), .A2(G217), .ZN(n542) );
  XNOR2_X1 U665 ( .A(n543), .B(n542), .ZN(n561) );
  INV_X1 U666 ( .A(KEYINPUT95), .ZN(n545) );
  AND2_X1 U667 ( .A1(G221), .A2(n586), .ZN(n548) );
  XNOR2_X1 U668 ( .A(n552), .B(n551), .ZN(n556) );
  XNOR2_X1 U669 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U670 ( .A(n556), .B(n555), .Z(n557) );
  XNOR2_X1 U671 ( .A(n558), .B(n557), .ZN(n787) );
  NOR2_X1 U672 ( .A1(n787), .A2(G902), .ZN(n559) );
  INV_X1 U673 ( .A(n559), .ZN(n560) );
  NAND2_X1 U674 ( .A1(n562), .A2(G221), .ZN(n564) );
  INV_X1 U675 ( .A(KEYINPUT21), .ZN(n563) );
  XNOR2_X1 U676 ( .A(n564), .B(n563), .ZN(n749) );
  INV_X1 U677 ( .A(n749), .ZN(n565) );
  AND2_X1 U678 ( .A1(n647), .A2(n744), .ZN(n566) );
  NAND2_X1 U679 ( .A1(n591), .A2(G210), .ZN(n567) );
  XNOR2_X1 U680 ( .A(n568), .B(n567), .ZN(n572) );
  XNOR2_X1 U681 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U682 ( .A(n576), .B(n575), .ZN(n705) );
  NAND2_X1 U683 ( .A1(n705), .A2(n577), .ZN(n578) );
  XNOR2_X2 U684 ( .A(n578), .B(G472), .ZN(n748) );
  INV_X1 U685 ( .A(n748), .ZN(n632) );
  NOR2_X1 U686 ( .A1(n632), .A2(n644), .ZN(n580) );
  XNOR2_X1 U687 ( .A(KEYINPUT64), .B(KEYINPUT1), .ZN(n579) );
  NAND2_X1 U688 ( .A1(n580), .A2(n745), .ZN(n754) );
  XNOR2_X1 U689 ( .A(n405), .B(KEYINPUT31), .ZN(n736) );
  XNOR2_X1 U690 ( .A(G134), .B(n581), .ZN(n585) );
  XOR2_X1 U691 ( .A(n583), .B(n582), .Z(n584) );
  XNOR2_X1 U692 ( .A(n585), .B(n584), .ZN(n590) );
  XOR2_X1 U693 ( .A(KEYINPUT9), .B(KEYINPUT105), .Z(n588) );
  XNOR2_X1 U694 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U695 ( .A(KEYINPUT104), .B(KEYINPUT13), .ZN(n603) );
  XOR2_X1 U696 ( .A(KEYINPUT101), .B(KEYINPUT12), .Z(n593) );
  NAND2_X1 U697 ( .A1(n591), .A2(G214), .ZN(n592) );
  XNOR2_X1 U698 ( .A(n593), .B(n592), .ZN(n597) );
  XOR2_X1 U699 ( .A(KEYINPUT11), .B(KEYINPUT102), .Z(n595) );
  XNOR2_X1 U700 ( .A(G143), .B(KEYINPUT103), .ZN(n594) );
  XNOR2_X1 U701 ( .A(n595), .B(n594), .ZN(n596) );
  XOR2_X1 U702 ( .A(n597), .B(n596), .Z(n599) );
  XNOR2_X1 U703 ( .A(n599), .B(n598), .ZN(n602) );
  XNOR2_X1 U704 ( .A(n601), .B(n600), .ZN(n805) );
  INV_X1 U705 ( .A(G475), .ZN(n604) );
  NAND2_X1 U706 ( .A1(n606), .A2(n614), .ZN(n737) );
  INV_X1 U707 ( .A(n737), .ZN(n727) );
  NOR2_X1 U708 ( .A1(n727), .A2(n668), .ZN(n763) );
  INV_X1 U709 ( .A(n763), .ZN(n605) );
  INV_X1 U710 ( .A(n606), .ZN(n613) );
  NAND2_X1 U711 ( .A1(n613), .A2(n614), .ZN(n607) );
  INV_X1 U712 ( .A(KEYINPUT6), .ZN(n608) );
  XNOR2_X1 U713 ( .A(n748), .B(n608), .ZN(n665) );
  XNOR2_X1 U714 ( .A(n609), .B(KEYINPUT83), .ZN(n610) );
  XNOR2_X1 U715 ( .A(n626), .B(KEYINPUT107), .ZN(n750) );
  NAND2_X1 U716 ( .A1(n610), .A2(n750), .ZN(n718) );
  AND2_X1 U717 ( .A1(n745), .A2(n744), .ZN(n611) );
  NAND2_X1 U718 ( .A1(n665), .A2(n611), .ZN(n612) );
  NOR2_X1 U719 ( .A1(n614), .A2(n613), .ZN(n654) );
  INV_X1 U720 ( .A(KEYINPUT75), .ZN(n615) );
  XNOR2_X1 U721 ( .A(n615), .B(KEYINPUT35), .ZN(n616) );
  INV_X1 U722 ( .A(KEYINPUT84), .ZN(n618) );
  BUF_X1 U723 ( .A(n624), .Z(n622) );
  NAND2_X1 U724 ( .A1(n622), .A2(KEYINPUT44), .ZN(n623) );
  NOR2_X1 U725 ( .A1(n702), .A2(KEYINPUT44), .ZN(n625) );
  NOR2_X1 U726 ( .A1(G900), .A2(n627), .ZN(n628) );
  NAND2_X1 U727 ( .A1(G953), .A2(n628), .ZN(n629) );
  XOR2_X1 U728 ( .A(KEYINPUT111), .B(n629), .Z(n630) );
  NAND2_X1 U729 ( .A1(n631), .A2(n630), .ZN(n646) );
  NOR2_X1 U730 ( .A1(n666), .A2(n632), .ZN(n633) );
  XOR2_X1 U731 ( .A(KEYINPUT28), .B(n633), .Z(n636) );
  INV_X1 U732 ( .A(KEYINPUT112), .ZN(n634) );
  XNOR2_X1 U733 ( .A(n647), .B(n634), .ZN(n635) );
  NOR2_X1 U734 ( .A1(n636), .A2(n635), .ZN(n660) );
  INV_X1 U735 ( .A(n660), .ZN(n641) );
  XNOR2_X1 U736 ( .A(KEYINPUT73), .B(KEYINPUT38), .ZN(n638) );
  NOR2_X1 U737 ( .A1(n759), .A2(n758), .ZN(n639) );
  AND2_X1 U738 ( .A1(n748), .A2(n683), .ZN(n643) );
  XNOR2_X1 U739 ( .A(n643), .B(n642), .ZN(n645) );
  NOR2_X1 U740 ( .A1(n645), .A2(n644), .ZN(n649) );
  NAND2_X1 U741 ( .A1(n649), .A2(n648), .ZN(n653) );
  AND2_X1 U742 ( .A1(n668), .A2(n689), .ZN(n651) );
  XNOR2_X1 U743 ( .A(n651), .B(KEYINPUT40), .ZN(n814) );
  XNOR2_X1 U744 ( .A(KEYINPUT46), .B(KEYINPUT80), .ZN(n652) );
  INV_X1 U745 ( .A(n653), .ZN(n655) );
  NAND2_X1 U746 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U747 ( .A1(n687), .A2(n656), .ZN(n731) );
  NOR2_X1 U748 ( .A1(KEYINPUT47), .A2(KEYINPUT76), .ZN(n657) );
  NOR2_X1 U749 ( .A1(n731), .A2(n657), .ZN(n664) );
  NAND2_X1 U750 ( .A1(n763), .A2(KEYINPUT76), .ZN(n661) );
  BUF_X1 U751 ( .A(n658), .Z(n659) );
  NAND2_X1 U752 ( .A1(n660), .A2(n659), .ZN(n678) );
  INV_X1 U753 ( .A(n678), .ZN(n732) );
  NAND2_X1 U754 ( .A1(n661), .A2(n732), .ZN(n662) );
  NAND2_X1 U755 ( .A1(n662), .A2(KEYINPUT47), .ZN(n663) );
  NAND2_X1 U756 ( .A1(n664), .A2(n663), .ZN(n675) );
  NAND2_X1 U757 ( .A1(n669), .A2(n719), .ZN(n682) );
  INV_X1 U758 ( .A(KEYINPUT114), .ZN(n670) );
  XNOR2_X1 U759 ( .A(n682), .B(n670), .ZN(n672) );
  INV_X1 U760 ( .A(KEYINPUT76), .ZN(n680) );
  NOR2_X1 U761 ( .A1(n678), .A2(KEYINPUT47), .ZN(n679) );
  NOR2_X1 U762 ( .A1(n680), .A2(n679), .ZN(n681) );
  INV_X1 U763 ( .A(n682), .ZN(n684) );
  INV_X1 U764 ( .A(n758), .ZN(n683) );
  AND2_X1 U765 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U766 ( .A1(n685), .A2(n429), .ZN(n686) );
  XNOR2_X1 U767 ( .A(n686), .B(KEYINPUT43), .ZN(n688) );
  NAND2_X1 U768 ( .A1(n688), .A2(n687), .ZN(n743) );
  NAND2_X1 U769 ( .A1(n727), .A2(n689), .ZN(n741) );
  NOR2_X2 U770 ( .A1(n693), .A2(n690), .ZN(n692) );
  INV_X1 U771 ( .A(n693), .ZN(n790) );
  NAND2_X1 U772 ( .A1(n790), .A2(n694), .ZN(n695) );
  INV_X1 U773 ( .A(G952), .ZN(n698) );
  AND2_X1 U774 ( .A1(n698), .A2(G953), .ZN(n789) );
  XNOR2_X1 U775 ( .A(n701), .B(n700), .ZN(G63) );
  XOR2_X1 U776 ( .A(G122), .B(n702), .Z(G24) );
  XNOR2_X1 U777 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n703) );
  XOR2_X1 U778 ( .A(n703), .B(KEYINPUT62), .Z(n704) );
  XNOR2_X1 U779 ( .A(n705), .B(n704), .ZN(n706) );
  INV_X1 U780 ( .A(n789), .ZN(n709) );
  XOR2_X1 U781 ( .A(KEYINPUT87), .B(KEYINPUT63), .Z(n707) );
  NAND2_X1 U782 ( .A1(n710), .A2(n709), .ZN(n712) );
  XNOR2_X1 U783 ( .A(KEYINPUT65), .B(KEYINPUT60), .ZN(n711) );
  XNOR2_X1 U784 ( .A(n712), .B(n711), .ZN(G60) );
  NAND2_X1 U785 ( .A1(n785), .A2(G469), .ZN(n716) );
  XOR2_X1 U786 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n713) );
  XNOR2_X1 U787 ( .A(n714), .B(n713), .ZN(n715) );
  XNOR2_X1 U788 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X1 U789 ( .A1(n717), .A2(n789), .ZN(G54) );
  XNOR2_X1 U790 ( .A(G101), .B(n718), .ZN(G3) );
  INV_X1 U791 ( .A(n719), .ZN(n734) );
  NOR2_X1 U792 ( .A1(n734), .A2(n417), .ZN(n720) );
  XOR2_X1 U793 ( .A(KEYINPUT118), .B(n720), .Z(n721) );
  XNOR2_X1 U794 ( .A(G104), .B(n721), .ZN(G6) );
  NOR2_X1 U795 ( .A1(n417), .A2(n737), .ZN(n724) );
  XNOR2_X1 U796 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n723) );
  XNOR2_X1 U797 ( .A(n724), .B(n723), .ZN(n725) );
  XNOR2_X1 U798 ( .A(G107), .B(n725), .ZN(G9) );
  XNOR2_X1 U799 ( .A(n726), .B(G110), .ZN(G12) );
  XOR2_X1 U800 ( .A(KEYINPUT119), .B(KEYINPUT29), .Z(n729) );
  NAND2_X1 U801 ( .A1(n732), .A2(n727), .ZN(n728) );
  XNOR2_X1 U802 ( .A(n729), .B(n728), .ZN(n730) );
  XOR2_X1 U803 ( .A(n471), .B(n730), .Z(G30) );
  XOR2_X1 U804 ( .A(G143), .B(n731), .Z(G45) );
  NAND2_X1 U805 ( .A1(n719), .A2(n732), .ZN(n733) );
  XNOR2_X1 U806 ( .A(n733), .B(G146), .ZN(G48) );
  NOR2_X1 U807 ( .A1(n734), .A2(n736), .ZN(n735) );
  XOR2_X1 U808 ( .A(G113), .B(n735), .Z(G15) );
  NOR2_X1 U809 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U810 ( .A(G116), .B(n738), .Z(G18) );
  XNOR2_X1 U811 ( .A(n739), .B(G125), .ZN(n740) );
  XNOR2_X1 U812 ( .A(n740), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U813 ( .A(G134), .B(KEYINPUT120), .ZN(n742) );
  XNOR2_X1 U814 ( .A(n742), .B(n741), .ZN(G36) );
  XNOR2_X1 U815 ( .A(G140), .B(n743), .ZN(G42) );
  NOR2_X1 U816 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U817 ( .A(n746), .B(KEYINPUT50), .ZN(n747) );
  NOR2_X1 U818 ( .A1(n748), .A2(n747), .ZN(n753) );
  NOR2_X1 U819 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U820 ( .A(n751), .B(KEYINPUT49), .ZN(n752) );
  NAND2_X1 U821 ( .A1(n753), .A2(n752), .ZN(n755) );
  NAND2_X1 U822 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U823 ( .A(KEYINPUT51), .B(n756), .ZN(n757) );
  NOR2_X1 U824 ( .A1(n757), .A2(n773), .ZN(n769) );
  AND2_X1 U825 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U826 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U827 ( .A(KEYINPUT121), .B(n762), .Z(n765) );
  NOR2_X1 U828 ( .A1(n765), .A2(n764), .ZN(n767) );
  INV_X1 U829 ( .A(n774), .ZN(n766) );
  NOR2_X1 U830 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U831 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U832 ( .A(n770), .B(KEYINPUT52), .ZN(n771) );
  NOR2_X1 U833 ( .A1(n772), .A2(n771), .ZN(n777) );
  NAND2_X1 U834 ( .A1(n448), .A2(n774), .ZN(n775) );
  NAND2_X1 U835 ( .A1(n775), .A2(n806), .ZN(n776) );
  XNOR2_X1 U836 ( .A(n779), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U837 ( .A(KEYINPUT88), .B(KEYINPUT55), .Z(n782) );
  XNOR2_X1 U838 ( .A(KEYINPUT122), .B(KEYINPUT54), .ZN(n781) );
  XNOR2_X1 U839 ( .A(n782), .B(n781), .ZN(n783) );
  NAND2_X1 U840 ( .A1(n785), .A2(G217), .ZN(n786) );
  XNOR2_X1 U841 ( .A(n787), .B(n786), .ZN(n788) );
  NOR2_X1 U842 ( .A1(n789), .A2(n788), .ZN(G66) );
  NAND2_X1 U843 ( .A1(n790), .A2(n806), .ZN(n794) );
  NAND2_X1 U844 ( .A1(G953), .A2(G224), .ZN(n791) );
  XNOR2_X1 U845 ( .A(KEYINPUT61), .B(n791), .ZN(n792) );
  NAND2_X1 U846 ( .A1(n792), .A2(G898), .ZN(n793) );
  NAND2_X1 U847 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U848 ( .A(n795), .B(KEYINPUT125), .ZN(n801) );
  XOR2_X1 U849 ( .A(G101), .B(KEYINPUT124), .Z(n796) );
  XNOR2_X1 U850 ( .A(n797), .B(n796), .ZN(n798) );
  NOR2_X1 U851 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U852 ( .A(n801), .B(n800), .Z(G69) );
  XNOR2_X1 U853 ( .A(n802), .B(n803), .ZN(n804) );
  XNOR2_X1 U854 ( .A(n805), .B(n804), .ZN(n809) );
  NAND2_X1 U855 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U856 ( .A(n808), .B(KEYINPUT126), .ZN(n813) );
  XNOR2_X1 U857 ( .A(G227), .B(n809), .ZN(n810) );
  NAND2_X1 U858 ( .A1(n810), .A2(G900), .ZN(n811) );
  NAND2_X1 U859 ( .A1(n811), .A2(G953), .ZN(n812) );
  NAND2_X1 U860 ( .A1(n813), .A2(n812), .ZN(G72) );
  XNOR2_X1 U861 ( .A(G131), .B(KEYINPUT127), .ZN(n815) );
  XNOR2_X1 U862 ( .A(n815), .B(n814), .ZN(G33) );
  XOR2_X1 U863 ( .A(n816), .B(G137), .Z(G39) );
endmodule

