//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n559,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(KEYINPUT68), .B(KEYINPUT2), .Z(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  OR4_X1    g030(.A1(G237), .A2(G238), .A3(G235), .A4(G236), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n455), .A2(new_n456), .ZN(G325));
  XOR2_X1   g032(.A(G325), .B(KEYINPUT69), .Z(G261));
  NAND2_X1  g033(.A1(new_n455), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI211_X1 g040(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT70), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT70), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n466), .A2(new_n470), .A3(new_n467), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  OR2_X1    g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  OAI21_X1  g052(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  XOR2_X1   g054(.A(new_n479), .B(KEYINPUT71), .Z(G160));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT73), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n464), .A2(new_n465), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(new_n463), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n483), .B1(G124), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n484), .A2(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT72), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(G2105), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n485), .B2(G126), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n464), .B2(new_n465), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT74), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n497), .B(KEYINPUT74), .C1(new_n465), .C2(new_n464), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n500), .A2(KEYINPUT75), .A3(KEYINPUT4), .A4(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT76), .B1(new_n498), .B2(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n463), .A2(G138), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n504), .B1(new_n474), .B2(new_n475), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT76), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n502), .A2(new_n503), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n507), .B1(new_n498), .B2(new_n499), .ZN(new_n510));
  AOI21_X1  g085(.A(KEYINPUT75), .B1(new_n510), .B2(new_n501), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n495), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT5), .B(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G62), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n515), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n519));
  XOR2_X1   g094(.A(KEYINPUT6), .B(G651), .Z(new_n520));
  OAI22_X1  g095(.A1(new_n518), .A2(KEYINPUT77), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n518), .A2(KEYINPUT77), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n521), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  INV_X1    g099(.A(KEYINPUT78), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT6), .B(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT78), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n526), .A2(G543), .A3(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G51), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n515), .A2(new_n527), .ZN(new_n535));
  INV_X1    g110(.A(G89), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n533), .B(new_n534), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n531), .A2(new_n537), .ZN(G168));
  AND3_X1   g113(.A1(new_n526), .A2(G543), .A3(new_n528), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G52), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n515), .A2(G64), .ZN(new_n541));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n514), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n535), .ZN(new_n544));
  XOR2_X1   g119(.A(KEYINPUT79), .B(G90), .Z(new_n545));
  AOI21_X1  g120(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n540), .A2(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  AOI22_X1  g123(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n514), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(KEYINPUT80), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n552), .B2(new_n535), .ZN(new_n553));
  INV_X1    g128(.A(G43), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n550), .A2(KEYINPUT80), .B1(new_n529), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g133(.A(KEYINPUT81), .B(KEYINPUT8), .Z(new_n559));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  AOI22_X1  g137(.A1(new_n515), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n563), .A2(new_n514), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT83), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g141(.A(KEYINPUT83), .B1(new_n563), .B2(new_n514), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n566), .A2(new_n567), .B1(G91), .B2(new_n544), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n539), .A2(new_n569), .A3(G53), .ZN(new_n570));
  INV_X1    g145(.A(G53), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT9), .B1(new_n529), .B2(new_n571), .ZN(new_n572));
  AND3_X1   g147(.A1(new_n570), .A2(KEYINPUT82), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g148(.A(KEYINPUT82), .B1(new_n570), .B2(new_n572), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n568), .B1(new_n573), .B2(new_n574), .ZN(G299));
  INV_X1    g150(.A(G168), .ZN(G286));
  NAND2_X1  g151(.A1(new_n544), .A2(G87), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n578));
  INV_X1    g153(.A(G49), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n577), .B(new_n578), .C1(new_n529), .C2(new_n579), .ZN(G288));
  NAND3_X1  g155(.A1(new_n515), .A2(new_n527), .A3(G86), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(KEYINPUT85), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n527), .A2(G48), .A3(G543), .ZN(new_n583));
  AND2_X1   g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n515), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n585));
  OR3_X1    g160(.A1(new_n585), .A2(KEYINPUT84), .A3(new_n514), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n581), .A2(KEYINPUT85), .ZN(new_n587));
  OAI21_X1  g162(.A(KEYINPUT84), .B1(new_n585), .B2(new_n514), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n584), .A2(new_n586), .A3(new_n587), .A4(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n514), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(KEYINPUT86), .B1(G85), .B2(new_n544), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n539), .A2(G47), .ZN(new_n593));
  OAI211_X1 g168(.A(new_n592), .B(new_n593), .C1(KEYINPUT86), .C2(new_n591), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n544), .A2(G92), .ZN(new_n596));
  XOR2_X1   g171(.A(KEYINPUT87), .B(KEYINPUT10), .Z(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n539), .A2(G54), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n515), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n600), .A2(new_n514), .ZN(new_n601));
  AND3_X1   g176(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n595), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n595), .B1(new_n602), .B2(G868), .ZN(G321));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(new_n568), .ZN(new_n606));
  INV_X1    g181(.A(new_n574), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n570), .A2(KEYINPUT82), .A3(new_n572), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n605), .B1(new_n609), .B2(G868), .ZN(G297));
  OAI21_X1  g185(.A(new_n605), .B1(new_n609), .B2(G868), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n602), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n602), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n487), .A2(G135), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n485), .A2(G123), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n463), .A2(G111), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n618), .B(new_n619), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(G2096), .Z(new_n623));
  NAND3_X1  g198(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  INV_X1    g201(.A(G2100), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n623), .A2(new_n628), .A3(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT88), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2427), .B(G2430), .Z(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(G14), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n642), .A2(new_n643), .ZN(new_n647));
  AND2_X1   g222(.A1(new_n647), .A2(KEYINPUT89), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n647), .A2(KEYINPUT89), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(G401));
  XOR2_X1   g226(.A(G2072), .B(G2078), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT17), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n655), .B2(new_n652), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n656), .B1(KEYINPUT90), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(KEYINPUT90), .B2(new_n658), .ZN(new_n660));
  INV_X1    g235(.A(new_n652), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n661), .A2(new_n657), .A3(new_n654), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT18), .Z(new_n663));
  NAND3_X1  g238(.A1(new_n653), .A2(new_n657), .A3(new_n655), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n660), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2096), .B(G2100), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1981), .B(G1986), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1956), .B(G2474), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1961), .B(G1966), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT20), .Z(new_n678));
  NAND2_X1  g253(.A1(new_n673), .A2(KEYINPUT92), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n674), .A2(new_n675), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(new_n672), .B2(new_n676), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n679), .B(new_n681), .Z(new_n682));
  NAND2_X1  g257(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1991), .B(G1996), .Z(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n685), .A2(new_n687), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n669), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n685), .A2(new_n687), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n692), .A2(new_n668), .A3(new_n688), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(G229));
  NOR2_X1   g270(.A1(G29), .A2(G35), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G162), .B2(G29), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT29), .B(G2090), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G21), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G168), .B2(new_n700), .ZN(new_n702));
  INV_X1    g277(.A(G1966), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n700), .A2(G19), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(new_n556), .B2(new_n700), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n706), .A2(G1341), .ZN(new_n707));
  INV_X1    g282(.A(G28), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n708), .A2(KEYINPUT30), .ZN(new_n709));
  AOI21_X1  g284(.A(G29), .B1(new_n708), .B2(KEYINPUT30), .ZN(new_n710));
  OR2_X1    g285(.A1(KEYINPUT31), .A2(G11), .ZN(new_n711));
  NAND2_X1  g286(.A1(KEYINPUT31), .A2(G11), .ZN(new_n712));
  AOI22_X1  g287(.A1(new_n709), .A2(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G32), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n487), .A2(G141), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n485), .A2(G129), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n463), .A2(G105), .A3(G2104), .ZN(new_n718));
  NAND3_X1  g293(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT26), .Z(new_n720));
  NAND4_X1  g295(.A1(new_n716), .A2(new_n717), .A3(new_n718), .A4(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n715), .B1(new_n722), .B2(new_n714), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT27), .B(G1996), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  OAI221_X1 g300(.A(new_n713), .B1(new_n714), .B2(new_n622), .C1(new_n723), .C2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n700), .A2(G5), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G171), .B2(new_n700), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n726), .B1(G1961), .B2(new_n728), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n699), .A2(new_n704), .A3(new_n707), .A4(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(G115), .A2(G2104), .ZN(new_n731));
  INV_X1    g306(.A(G127), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n484), .B2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT98), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n463), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n734), .B2(new_n733), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT25), .ZN(new_n737));
  NAND2_X1  g312(.A1(G103), .A2(G2104), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(G2105), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n463), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n487), .A2(G139), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  MUX2_X1   g317(.A(G33), .B(new_n742), .S(G29), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2072), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n714), .A2(G26), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT28), .Z(new_n746));
  NAND2_X1  g321(.A1(new_n487), .A2(G140), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n485), .A2(G128), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n463), .A2(G116), .ZN(new_n749));
  OAI21_X1  g324(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n747), .B(new_n748), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT97), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n746), .B1(new_n753), .B2(G29), .ZN(new_n754));
  INV_X1    g329(.A(G2067), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NOR3_X1   g331(.A1(new_n730), .A2(new_n744), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n700), .A2(G20), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT23), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n609), .B2(new_n700), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1956), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n723), .A2(new_n725), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n728), .B2(G1961), .ZN(new_n763));
  NAND2_X1  g338(.A1(G160), .A2(G29), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT99), .B(KEYINPUT24), .Z(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G34), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n764), .B1(G29), .B2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(G2084), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n763), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n761), .B1(KEYINPUT100), .B2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(G2078), .ZN(new_n771));
  NOR2_X1   g346(.A1(G164), .A2(new_n714), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G27), .B2(new_n714), .ZN(new_n773));
  OAI22_X1  g348(.A1(new_n767), .A2(new_n768), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G4), .A2(G16), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n602), .B2(G16), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT96), .B(G1348), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n773), .A2(new_n771), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n706), .A2(G1341), .ZN(new_n780));
  NOR4_X1   g355(.A1(new_n774), .A2(new_n778), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n769), .A2(KEYINPUT100), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n757), .A2(new_n770), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  OR2_X1    g358(.A1(G6), .A2(G16), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G305), .B2(new_n700), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT93), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT32), .B(G1981), .Z(new_n787));
  OR2_X1    g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(G23), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n789), .A2(G16), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G288), .B2(G16), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT94), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT33), .B(G1976), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n788), .A2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT34), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n700), .A2(G22), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G303), .B2(G16), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT95), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n802), .A2(G1971), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  INV_X1    g380(.A(G1971), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n805), .A2(new_n806), .B1(new_n787), .B2(new_n786), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n797), .A2(new_n798), .A3(new_n804), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n804), .ZN(new_n809));
  OAI21_X1  g384(.A(KEYINPUT34), .B1(new_n809), .B2(new_n796), .ZN(new_n810));
  MUX2_X1   g385(.A(G24), .B(G290), .S(G16), .Z(new_n811));
  AND2_X1   g386(.A1(new_n811), .A2(G1986), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n811), .A2(G1986), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n714), .A2(G25), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n487), .A2(G131), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n485), .A2(G119), .ZN(new_n816));
  OR2_X1    g391(.A1(G95), .A2(G2105), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n817), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n815), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n814), .B1(new_n820), .B2(new_n714), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT35), .B(G1991), .Z(new_n822));
  XOR2_X1   g397(.A(new_n821), .B(new_n822), .Z(new_n823));
  NOR3_X1   g398(.A1(new_n812), .A2(new_n813), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n808), .A2(new_n810), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(KEYINPUT36), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT36), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n808), .A2(new_n810), .A3(new_n827), .A4(new_n824), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n783), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT101), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(G311));
  INV_X1    g406(.A(new_n829), .ZN(G150));
  NAND2_X1  g407(.A1(new_n539), .A2(G55), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n834), .A2(new_n514), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n544), .A2(G93), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n833), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(G860), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT37), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n602), .A2(G559), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n837), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n556), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n837), .B1(new_n553), .B2(new_n555), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n842), .B(new_n846), .Z(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n849));
  INV_X1    g424(.A(G860), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(new_n848), .B2(KEYINPUT39), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n839), .B1(new_n849), .B2(new_n851), .ZN(G145));
  XNOR2_X1  g427(.A(new_n753), .B(new_n512), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n820), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n485), .A2(G130), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n463), .A2(G118), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n858), .B1(G142), .B2(new_n487), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(new_n625), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n742), .B(new_n722), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n854), .B(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(G160), .B(G162), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n622), .ZN(new_n865));
  AOI21_X1  g440(.A(G37), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n863), .A2(new_n865), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT103), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR3_X1   g444(.A1(new_n863), .A2(KEYINPUT103), .A3(new_n865), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n866), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(KEYINPUT104), .B(KEYINPUT40), .Z(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(G395));
  NAND2_X1  g448(.A1(new_n609), .A2(new_n602), .ZN(new_n874));
  INV_X1    g449(.A(new_n602), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(G299), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(KEYINPUT41), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT41), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n874), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n846), .B(new_n614), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  OR3_X1    g460(.A1(new_n883), .A2(KEYINPUT105), .A3(new_n877), .ZN(new_n886));
  OAI21_X1  g461(.A(KEYINPUT105), .B1(new_n883), .B2(new_n877), .ZN(new_n887));
  AOI22_X1  g462(.A1(KEYINPUT106), .A2(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n885), .A2(KEYINPUT106), .ZN(new_n889));
  XOR2_X1   g464(.A(G303), .B(G305), .Z(new_n890));
  INV_X1    g465(.A(G288), .ZN(new_n891));
  XNOR2_X1  g466(.A(G290), .B(new_n891), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n890), .B(new_n892), .Z(new_n893));
  XOR2_X1   g468(.A(new_n893), .B(KEYINPUT42), .Z(new_n894));
  AND3_X1   g469(.A1(new_n888), .A2(new_n889), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n894), .B1(new_n888), .B2(new_n889), .ZN(new_n896));
  OAI21_X1  g471(.A(G868), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(G868), .B2(new_n843), .ZN(G295));
  OAI21_X1  g473(.A(new_n897), .B1(G868), .B2(new_n843), .ZN(G331));
  INV_X1    g474(.A(G37), .ZN(new_n900));
  AOI21_X1  g475(.A(G171), .B1(G286), .B2(KEYINPUT107), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  OR3_X1    g477(.A1(new_n531), .A2(KEYINPUT107), .A3(new_n537), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n844), .A2(new_n845), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n903), .B1(new_n844), .B2(new_n845), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n903), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n846), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n909), .A2(new_n901), .A3(new_n904), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n881), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n893), .ZN(new_n913));
  INV_X1    g488(.A(new_n877), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n914), .A2(new_n907), .A3(new_n910), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n912), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n879), .B1(new_n874), .B2(new_n876), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n910), .A2(new_n907), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n878), .A2(KEYINPUT108), .A3(new_n880), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n907), .A2(new_n910), .ZN(new_n921));
  AOI22_X1  g496(.A1(new_n919), .A2(new_n920), .B1(new_n921), .B2(new_n914), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n900), .B(new_n916), .C1(new_n922), .C2(new_n913), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT109), .B1(new_n923), .B2(KEYINPUT43), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n916), .A2(new_n900), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n919), .A2(new_n920), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n915), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n893), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n925), .A2(new_n926), .A3(new_n929), .A4(new_n930), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n912), .A2(new_n915), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n932), .A2(new_n913), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n916), .A2(new_n900), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT43), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n924), .A2(new_n931), .A3(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n933), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT43), .B1(new_n939), .B2(new_n925), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n923), .A2(new_n930), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT44), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n938), .A2(new_n942), .ZN(G397));
  INV_X1    g518(.A(G1384), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n512), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT45), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n466), .A2(new_n470), .A3(new_n467), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n470), .B1(new_n466), .B2(new_n467), .ZN(new_n949));
  OAI211_X1 g524(.A(G40), .B(new_n478), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT110), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n472), .A2(KEYINPUT110), .A3(G40), .A4(new_n478), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n947), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n753), .B(G2067), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT112), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n753), .B(new_n755), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT112), .ZN(new_n960));
  INV_X1    g535(.A(G1996), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n721), .B(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n819), .B(new_n822), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n958), .A2(new_n960), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT111), .B1(G290), .B2(G1986), .ZN(new_n965));
  NAND2_X1  g540(.A1(G290), .A2(G1986), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n965), .B(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n955), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT113), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT51), .ZN(new_n970));
  NAND2_X1  g545(.A1(G286), .A2(G8), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n971), .B(KEYINPUT120), .Z(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n952), .A2(new_n953), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT75), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT4), .B1(new_n505), .B2(KEYINPUT74), .ZN(new_n976));
  INV_X1    g551(.A(new_n501), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n503), .A2(new_n508), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(new_n979), .A3(new_n502), .ZN(new_n980));
  AOI21_X1  g555(.A(G1384), .B1(new_n980), .B2(new_n495), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT50), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n974), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AOI211_X1 g558(.A(KEYINPUT50), .B(G1384), .C1(new_n980), .C2(new_n495), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n981), .A2(KEYINPUT45), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n947), .A2(new_n974), .A3(new_n986), .ZN(new_n987));
  AOI22_X1  g562(.A1(new_n985), .A2(new_n768), .B1(new_n987), .B2(new_n703), .ZN(new_n988));
  INV_X1    g563(.A(G8), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n970), .B(new_n973), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT51), .B1(new_n988), .B2(new_n973), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n945), .A2(KEYINPUT50), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n981), .A2(new_n982), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n992), .A2(new_n993), .A3(new_n768), .A4(new_n974), .ZN(new_n994));
  AOI211_X1 g569(.A(new_n946), .B(G1384), .C1(new_n980), .C2(new_n495), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT45), .B1(new_n512), .B2(new_n944), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n995), .A2(new_n996), .A3(new_n954), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n994), .B1(new_n997), .B2(G1966), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n972), .B1(new_n998), .B2(G8), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n990), .B1(new_n991), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT62), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n995), .A2(new_n996), .ZN(new_n1004));
  AOI21_X1  g579(.A(G1971), .B1(new_n1004), .B2(new_n974), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n983), .A2(G2090), .A3(new_n984), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1003), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(G303), .A2(G8), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n1008), .B(KEYINPUT55), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n954), .B1(new_n945), .B2(KEYINPUT50), .ZN(new_n1011));
  INV_X1    g586(.A(G2090), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(new_n1012), .A3(new_n993), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1013), .B(KEYINPUT114), .C1(new_n997), .C2(G1971), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1007), .A2(G8), .A3(new_n1010), .A4(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n974), .A2(new_n981), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n891), .A2(G1976), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(G8), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT115), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n989), .B1(new_n974), .B2(new_n981), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1021), .A2(KEYINPUT115), .A3(new_n1017), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1020), .A2(KEYINPUT52), .A3(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n585), .A2(new_n514), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n581), .A2(new_n583), .ZN(new_n1025));
  OAI21_X1  g600(.A(G1981), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g601(.A(KEYINPUT116), .B(G1981), .ZN(new_n1027));
  OAI211_X1 g602(.A(KEYINPUT49), .B(new_n1026), .C1(G305), .C2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1026), .B1(G305), .B2(new_n1027), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT49), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1021), .A2(new_n1028), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G1976), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT52), .B1(G288), .B2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1021), .A2(new_n1017), .A3(new_n1034), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1023), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(G8), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n1009), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n1015), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G1961), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1011), .A2(new_n993), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n947), .A2(new_n986), .A3(new_n771), .A4(new_n974), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n1041), .A2(new_n1042), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n997), .A2(KEYINPUT53), .A3(new_n771), .ZN(new_n1046));
  AOI21_X1  g621(.A(G301), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1002), .A2(new_n1040), .A3(KEYINPUT122), .A4(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT122), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n973), .B1(new_n988), .B2(new_n989), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n970), .B1(new_n998), .B2(new_n972), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT62), .B1(new_n1052), .B2(new_n990), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1015), .A2(new_n1037), .A3(new_n1039), .A4(new_n1047), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1049), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1000), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT62), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1048), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1032), .A2(new_n1033), .A3(new_n891), .ZN(new_n1059));
  NOR2_X1   g634(.A1(G305), .A2(new_n1027), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n1060), .B(KEYINPUT117), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1021), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1023), .A2(new_n1036), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1062), .B1(new_n1015), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT118), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1066), .B(new_n1062), .C1(new_n1015), .C2(new_n1063), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n988), .A2(new_n989), .A3(G286), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1015), .A2(new_n1037), .A3(new_n1039), .A4(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT63), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1007), .A2(G8), .A3(new_n1014), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n1009), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1063), .A2(new_n1071), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1074), .A2(new_n1015), .A3(new_n1069), .A4(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1072), .A2(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT121), .B(KEYINPUT54), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n950), .A2(new_n1044), .A3(G2078), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1042), .A2(new_n1041), .B1(new_n1004), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1082), .A2(G171), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1078), .B1(new_n1083), .B2(new_n1047), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(G171), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1045), .A2(G301), .A3(new_n1046), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1085), .A2(KEYINPUT54), .A3(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1040), .A2(new_n1056), .A3(new_n1084), .A4(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G1956), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(new_n983), .B2(new_n984), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n570), .A2(new_n572), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n568), .ZN(new_n1092));
  XOR2_X1   g667(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1094), .B1(G299), .B2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT56), .B(G2072), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n947), .A2(new_n986), .A3(new_n974), .A4(new_n1097), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1090), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1090), .A2(new_n1098), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1096), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(G1348), .B1(new_n1011), .B2(new_n993), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n974), .A2(new_n755), .A3(new_n981), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n602), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1099), .B1(new_n1102), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT61), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1096), .B1(new_n1090), .B2(new_n1098), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1108), .B1(new_n1099), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1090), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1102), .A2(new_n1111), .A3(KEYINPUT61), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT60), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1114));
  OAI211_X1 g689(.A(KEYINPUT60), .B(new_n1104), .C1(new_n985), .C2(G1348), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1114), .A2(new_n1115), .A3(new_n602), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1110), .A2(new_n1112), .A3(new_n1116), .ZN(new_n1117));
  XOR2_X1   g692(.A(KEYINPUT58), .B(G1341), .Z(new_n1118));
  NAND2_X1  g693(.A1(new_n1016), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(new_n987), .B2(G1996), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1120), .A2(KEYINPUT59), .A3(new_n556), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1115), .A2(new_n602), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT59), .B1(new_n1120), .B2(new_n556), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1107), .B1(new_n1117), .B2(new_n1124), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1068), .B(new_n1077), .C1(new_n1088), .C2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n969), .B1(new_n1058), .B2(new_n1126), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n958), .A2(new_n960), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n962), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n820), .A2(new_n822), .ZN(new_n1130));
  OAI22_X1  g705(.A1(new_n1129), .A2(new_n1130), .B1(G2067), .B2(new_n753), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n955), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n964), .A2(new_n955), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT125), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1133), .B(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(G290), .A2(G1986), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n955), .A2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1137), .B(KEYINPUT126), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT48), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1135), .A2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1132), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n955), .A2(new_n961), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  OR2_X1    g720(.A1(new_n1145), .A2(KEYINPUT46), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1128), .A2(new_n722), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1147), .A2(new_n1148), .A3(new_n955), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1148), .B1(new_n1147), .B2(new_n955), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1146), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1145), .A2(KEYINPUT46), .ZN(new_n1152));
  XOR2_X1   g727(.A(new_n1152), .B(KEYINPUT123), .Z(new_n1153));
  OR3_X1    g728(.A1(new_n1151), .A2(KEYINPUT47), .A3(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT47), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1143), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1127), .A2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g732(.A1(G227), .A2(new_n461), .ZN(new_n1159));
  NAND2_X1  g733(.A1(new_n650), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g734(.A(KEYINPUT127), .B1(G229), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g735(.A(KEYINPUT127), .ZN(new_n1162));
  NAND4_X1  g736(.A1(new_n694), .A2(new_n650), .A3(new_n1162), .A4(new_n1159), .ZN(new_n1163));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  AND3_X1   g738(.A1(new_n936), .A2(new_n1164), .A3(new_n871), .ZN(G308));
  NAND3_X1  g739(.A1(new_n936), .A2(new_n1164), .A3(new_n871), .ZN(G225));
endmodule


