//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 1 1 0 1 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n555, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n598, new_n601, new_n603, new_n604, new_n605,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT64), .ZN(G319));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  OR2_X1    g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g038(.A(KEYINPUT65), .B1(new_n463), .B2(G125), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI211_X1 g041(.A(KEYINPUT65), .B(G125), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n460), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n463), .A2(G137), .A3(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G112), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n465), .A2(new_n466), .ZN(new_n482));
  OR3_X1    g057(.A1(new_n482), .A2(KEYINPUT66), .A3(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(KEYINPUT66), .B1(new_n482), .B2(G2105), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n482), .A2(new_n471), .ZN(new_n487));
  AOI211_X1 g062(.A(new_n481), .B(new_n486), .C1(G124), .C2(new_n487), .ZN(G162));
  OAI211_X1 g063(.A(G126), .B(G2105), .C1(new_n465), .C2(new_n466), .ZN(new_n489));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n490), .A2(new_n492), .A3(G2104), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n465), .B2(new_n466), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n463), .A2(new_n499), .A3(new_n496), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n494), .B1(new_n498), .B2(new_n500), .ZN(G164));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(KEYINPUT67), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT5), .A3(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT68), .B(G88), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G50), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT69), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n515), .B(new_n516), .ZN(new_n517));
  AOI21_X1  g092(.A(KEYINPUT70), .B1(new_n507), .B2(G62), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n518), .B1(G75), .B2(G543), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n507), .A2(KEYINPUT70), .A3(G62), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n517), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NOR2_X1   g099(.A1(new_n507), .A2(KEYINPUT71), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n526), .B1(new_n504), .B2(new_n506), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n528), .A2(G63), .A3(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n509), .A2(G89), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n513), .A2(G51), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n529), .A2(new_n534), .ZN(G168));
  INV_X1    g110(.A(G651), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n528), .A2(G64), .ZN(new_n537));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n509), .A2(G90), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n541), .B2(new_n512), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(G171));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  NOR3_X1   g119(.A1(new_n525), .A2(new_n544), .A3(new_n527), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT72), .ZN(new_n546));
  AND2_X1   g121(.A1(G68), .A2(G543), .ZN(new_n547));
  OR3_X1    g122(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n545), .B2(new_n547), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n548), .A2(G651), .A3(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n509), .A2(G81), .B1(new_n513), .B2(G43), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n555));
  XOR2_X1   g130(.A(new_n555), .B(KEYINPUT73), .Z(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  XOR2_X1   g134(.A(KEYINPUT75), .B(G65), .Z(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(new_n507), .ZN(new_n561));
  INV_X1    g136(.A(G78), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n562), .B2(new_n503), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n563), .A2(G651), .B1(G91), .B2(new_n509), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n513), .A2(KEYINPUT74), .A3(G53), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT74), .ZN(new_n566));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n512), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n565), .A2(KEYINPUT9), .A3(new_n568), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n568), .A2(KEYINPUT9), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n564), .A2(new_n569), .A3(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(G168), .ZN(G286));
  OAI21_X1  g148(.A(G651), .B1(new_n528), .B2(G74), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n509), .A2(G87), .B1(new_n513), .B2(G49), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(G288));
  AOI22_X1  g151(.A1(new_n507), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(new_n536), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n509), .A2(G86), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n513), .A2(G48), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G305));
  XNOR2_X1  g156(.A(KEYINPUT76), .B(G47), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n509), .A2(G85), .B1(new_n513), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n584), .B2(new_n536), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n507), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n536), .B1(new_n587), .B2(KEYINPUT77), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n588), .B1(KEYINPUT77), .B2(new_n587), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n507), .A2(G92), .A3(new_n508), .ZN(new_n590));
  XOR2_X1   g165(.A(new_n590), .B(KEYINPUT10), .Z(new_n591));
  NAND2_X1  g166(.A1(new_n513), .A2(G54), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n589), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n586), .B1(G868), .B2(new_n594), .ZN(G284));
  OAI21_X1  g170(.A(new_n586), .B1(G868), .B2(new_n594), .ZN(G321));
  NAND2_X1  g171(.A1(G286), .A2(G868), .ZN(new_n597));
  INV_X1    g172(.A(G299), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(G868), .B2(new_n598), .ZN(G297));
  XNOR2_X1  g174(.A(G297), .B(KEYINPUT78), .ZN(G280));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n594), .B1(new_n601), .B2(G860), .ZN(G148));
  NAND2_X1  g177(.A1(new_n594), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G868), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G868), .B2(new_n553), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT79), .ZN(G323));
  XOR2_X1   g181(.A(KEYINPUT80), .B(KEYINPUT11), .Z(new_n607));
  XNOR2_X1  g182(.A(G323), .B(new_n607), .ZN(G282));
  NAND2_X1  g183(.A1(new_n463), .A2(new_n474), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT12), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT13), .ZN(new_n611));
  INV_X1    g186(.A(G2100), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT81), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n485), .A2(G135), .ZN(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n616));
  INV_X1    g191(.A(G111), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G2105), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n618), .B1(new_n487), .B2(G123), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(G2096), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n621), .A2(new_n622), .B1(new_n611), .B2(new_n612), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n614), .B(new_n623), .C1(new_n622), .C2(new_n621), .ZN(G156));
  XNOR2_X1  g199(.A(G2451), .B(G2454), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2443), .B(G2446), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n625), .B(new_n626), .Z(new_n627));
  XNOR2_X1  g202(.A(G1341), .B(G1348), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2427), .B(G2430), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(KEYINPUT14), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT83), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n633), .A2(KEYINPUT83), .A3(KEYINPUT14), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n631), .A2(new_n632), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n629), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  AOI211_X1 g216(.A(new_n639), .B(new_n628), .C1(new_n636), .C2(new_n637), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n627), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(new_n637), .ZN(new_n644));
  AOI21_X1  g219(.A(KEYINPUT83), .B1(new_n633), .B2(KEYINPUT14), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n640), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(new_n628), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n638), .A2(new_n640), .A3(new_n629), .ZN(new_n648));
  INV_X1    g223(.A(new_n627), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n643), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n643), .A2(new_n652), .A3(new_n650), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(G14), .A3(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  XNOR2_X1  g232(.A(KEYINPUT85), .B(G2100), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT84), .ZN(new_n661));
  NOR2_X1   g236(.A1(G2072), .A2(G2078), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n442), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  NAND3_X1  g240(.A1(new_n661), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT18), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n663), .B(KEYINPUT17), .Z(new_n669));
  AOI21_X1  g244(.A(new_n665), .B1(new_n669), .B2(new_n661), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n670), .B1(new_n661), .B2(new_n664), .ZN(new_n671));
  INV_X1    g246(.A(new_n665), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n669), .A2(new_n661), .A3(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n668), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n675), .A2(G2096), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n666), .A2(new_n667), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n666), .A2(new_n667), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n673), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n622), .B1(new_n679), .B2(new_n671), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n659), .B1(new_n676), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n675), .A2(G2096), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n679), .A2(new_n622), .A3(new_n671), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n682), .A2(new_n683), .A3(new_n658), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n681), .A2(new_n684), .ZN(G227));
  XNOR2_X1  g260(.A(G1971), .B(G1976), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G1956), .B(G2474), .Z(new_n689));
  XOR2_X1   g264(.A(G1961), .B(G1966), .Z(new_n690));
  AND2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT20), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n689), .A2(new_n690), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  MUX2_X1   g271(.A(new_n696), .B(new_n695), .S(new_n688), .Z(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  OR3_X1    g274(.A1(new_n694), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(G1991), .B(G1996), .Z(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n699), .B1(new_n694), .B2(new_n697), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n700), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1981), .B(G1986), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n702), .B1(new_n700), .B2(new_n703), .ZN(new_n708));
  OR3_X1    g283(.A1(new_n705), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n707), .B1(new_n705), .B2(new_n708), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(G229));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G22), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G166), .B2(new_n713), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G1971), .ZN(new_n716));
  NOR2_X1   g291(.A1(G6), .A2(G16), .ZN(new_n717));
  AND3_X1   g292(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n717), .B1(new_n718), .B2(G16), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT32), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(G1981), .ZN(new_n721));
  NOR2_X1   g296(.A1(G16), .A2(G23), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT86), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G288), .B2(new_n713), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT33), .B(G1976), .Z(new_n725));
  XOR2_X1   g300(.A(new_n724), .B(new_n725), .Z(new_n726));
  NOR3_X1   g301(.A1(new_n716), .A2(new_n721), .A3(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT34), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G25), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n485), .A2(G131), .ZN(new_n733));
  OAI21_X1  g308(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n734));
  INV_X1    g309(.A(G107), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(G2105), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n487), .B2(G119), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n732), .B1(new_n739), .B2(new_n731), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT35), .B(G1991), .Z(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n740), .B(new_n742), .ZN(new_n743));
  MUX2_X1   g318(.A(G24), .B(G290), .S(G16), .Z(new_n744));
  NOR2_X1   g319(.A1(new_n744), .A2(G1986), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n744), .A2(G1986), .ZN(new_n746));
  NOR3_X1   g321(.A1(new_n743), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n729), .A2(new_n730), .A3(new_n747), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT36), .Z(new_n749));
  NAND2_X1  g324(.A1(new_n731), .A2(G35), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G162), .B2(new_n731), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT29), .B(G2090), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n485), .A2(G141), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n474), .A2(G105), .ZN(new_n755));
  NAND3_X1  g330(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT26), .ZN(new_n757));
  AOI211_X1 g332(.A(new_n755), .B(new_n757), .C1(G129), .C2(new_n487), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(G29), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT91), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n761), .B(new_n762), .C1(G29), .C2(G32), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n762), .B2(new_n761), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT27), .B(G1996), .Z(new_n765));
  OR2_X1    g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n731), .A2(G26), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT28), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n485), .A2(G140), .ZN(new_n770));
  NOR2_X1   g345(.A1(G104), .A2(G2105), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT88), .ZN(new_n772));
  INV_X1    g347(.A(G116), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n473), .B1(new_n773), .B2(G2105), .ZN(new_n774));
  AOI22_X1  g349(.A1(G128), .A2(new_n487), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n769), .B1(new_n776), .B2(G29), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G2067), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n753), .A2(new_n766), .A3(new_n767), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n621), .A2(G29), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT92), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n713), .A2(G21), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G168), .B2(new_n713), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n783), .A2(G1966), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(G1966), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n781), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(G29), .A2(G33), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT89), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT90), .B(KEYINPUT25), .Z(new_n789));
  NAND3_X1  g364(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n483), .A2(new_n484), .ZN(new_n793));
  INV_X1    g368(.A(G139), .ZN(new_n794));
  OAI221_X1 g369(.A(new_n791), .B1(new_n471), .B2(new_n792), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n788), .B1(new_n795), .B2(new_n731), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G2072), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT30), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n798), .A2(G28), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n731), .B1(new_n798), .B2(G28), .ZN(new_n800));
  AND2_X1   g375(.A1(KEYINPUT31), .A2(G11), .ZN(new_n801));
  NOR2_X1   g376(.A1(KEYINPUT31), .A2(G11), .ZN(new_n802));
  OAI22_X1  g377(.A1(new_n799), .A2(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(G164), .A2(G29), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G27), .B2(G29), .ZN(new_n805));
  INV_X1    g380(.A(G2078), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n803), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n797), .B(new_n807), .C1(new_n806), .C2(new_n805), .ZN(new_n808));
  NOR3_X1   g383(.A1(new_n779), .A2(new_n786), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n713), .A2(G20), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT23), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n598), .B2(new_n713), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(G1956), .Z(new_n813));
  NOR2_X1   g388(.A1(new_n594), .A2(new_n713), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G4), .B2(new_n713), .ZN(new_n815));
  INV_X1    g390(.A(G1348), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n713), .A2(G5), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G171), .B2(new_n713), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n817), .B1(G1961), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n553), .A2(G16), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G16), .B2(G19), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT87), .B(G1341), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT24), .ZN(new_n826));
  INV_X1    g401(.A(G34), .ZN(new_n827));
  AOI21_X1  g402(.A(G29), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n826), .B2(new_n827), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(G160), .B2(new_n731), .ZN(new_n830));
  INV_X1    g405(.A(G2084), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n815), .B2(new_n816), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n820), .A2(new_n825), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n819), .A2(G1961), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT93), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(new_n822), .B2(new_n824), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n809), .A2(new_n813), .A3(new_n834), .A4(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n749), .A2(new_n838), .ZN(G311));
  INV_X1    g414(.A(G311), .ZN(G150));
  NAND2_X1  g415(.A1(new_n594), .A2(G559), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT38), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n509), .A2(G93), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n513), .A2(G55), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(KEYINPUT94), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT94), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n843), .A2(new_n847), .A3(new_n844), .ZN(new_n848));
  NAND2_X1  g423(.A1(G80), .A2(G543), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n507), .B(KEYINPUT71), .ZN(new_n850));
  INV_X1    g425(.A(G67), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n846), .A2(new_n848), .B1(new_n852), .B2(G651), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n552), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n550), .A2(new_n853), .A3(new_n551), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n842), .B(new_n857), .Z(new_n858));
  OR2_X1    g433(.A1(new_n858), .A2(KEYINPUT39), .ZN(new_n859));
  INV_X1    g434(.A(G860), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(KEYINPUT39), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n853), .A2(new_n860), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT37), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(G145));
  XOR2_X1   g440(.A(KEYINPUT95), .B(G37), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n759), .B(new_n776), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n739), .ZN(new_n868));
  INV_X1    g443(.A(G164), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n795), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n487), .A2(G130), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n471), .A2(G118), .ZN(new_n872));
  OAI21_X1  g447(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n873));
  INV_X1    g448(.A(G142), .ZN(new_n874));
  OAI221_X1 g449(.A(new_n871), .B1(new_n872), .B2(new_n873), .C1(new_n793), .C2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n610), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n870), .B(new_n876), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n868), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n868), .A2(new_n877), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n620), .B(new_n477), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n881), .B(G162), .Z(new_n882));
  NOR2_X1   g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n882), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(new_n878), .B2(new_n879), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n866), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT40), .ZN(G395));
  OR2_X1    g462(.A1(G290), .A2(G288), .ZN(new_n888));
  NAND2_X1  g463(.A1(G290), .A2(G288), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT98), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n890), .A2(new_n891), .ZN(new_n894));
  AOI21_X1  g469(.A(KEYINPUT97), .B1(new_n517), .B2(new_n522), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n517), .A2(KEYINPUT97), .A3(new_n522), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(G305), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(G305), .B1(new_n896), .B2(new_n897), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n893), .B(new_n894), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n900), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n902), .A2(new_n892), .A3(new_n898), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  XOR2_X1   g479(.A(new_n904), .B(KEYINPUT42), .Z(new_n905));
  XNOR2_X1  g480(.A(new_n857), .B(new_n603), .ZN(new_n906));
  NAND2_X1  g481(.A1(G299), .A2(KEYINPUT96), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT96), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n564), .A2(new_n569), .A3(new_n570), .A4(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n594), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n593), .A2(G299), .A3(KEYINPUT96), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n906), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT41), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n910), .A2(new_n915), .A3(new_n911), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n915), .B1(new_n910), .B2(new_n911), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n914), .B1(new_n906), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT99), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n920), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n905), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n905), .A2(new_n922), .ZN(new_n924));
  OAI21_X1  g499(.A(G868), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n925), .B1(G868), .B2(new_n853), .ZN(G295));
  OAI21_X1  g501(.A(new_n925), .B1(G868), .B2(new_n853), .ZN(G331));
  INV_X1    g502(.A(new_n918), .ZN(new_n928));
  NOR2_X1   g503(.A1(G171), .A2(KEYINPUT100), .ZN(new_n929));
  INV_X1    g504(.A(new_n856), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n853), .B1(new_n550), .B2(new_n551), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n929), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n855), .A2(new_n933), .A3(new_n856), .ZN(new_n934));
  AOI21_X1  g509(.A(G286), .B1(G171), .B2(KEYINPUT100), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n932), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n935), .B1(new_n932), .B2(new_n934), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n928), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(KEYINPUT101), .ZN(new_n939));
  INV_X1    g514(.A(new_n935), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n930), .A2(new_n931), .A3(new_n929), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n933), .B1(new_n855), .B2(new_n856), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n932), .A2(new_n934), .A3(new_n935), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(new_n913), .A3(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT101), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n946), .B(new_n928), .C1(new_n936), .C2(new_n937), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n939), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n904), .A2(KEYINPUT102), .ZN(new_n949));
  AOI21_X1  g524(.A(G37), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n904), .A2(KEYINPUT102), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n939), .A2(new_n951), .A3(new_n945), .A4(new_n947), .ZN(new_n952));
  AOI21_X1  g527(.A(KEYINPUT43), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n904), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n939), .A2(new_n954), .A3(new_n945), .A4(new_n947), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n866), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT104), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n943), .A2(new_n944), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT103), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n912), .A2(new_n959), .A3(KEYINPUT41), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n960), .B1(new_n918), .B2(new_n959), .ZN(new_n961));
  AOI22_X1  g536(.A1(new_n945), .A2(new_n957), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n943), .A2(KEYINPUT104), .A3(new_n913), .A4(new_n944), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n954), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n956), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT44), .B1(new_n953), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n947), .A2(new_n945), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n946), .B1(new_n958), .B2(new_n928), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n949), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G37), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n970), .A2(new_n971), .A3(new_n952), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n945), .A2(new_n957), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n958), .A2(new_n961), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n974), .A2(new_n963), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n904), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n977), .A2(new_n965), .A3(new_n866), .A4(new_n955), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n973), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n967), .B1(new_n980), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g556(.A(KEYINPUT121), .ZN(new_n982));
  XOR2_X1   g557(.A(KEYINPUT119), .B(KEYINPUT51), .Z(new_n983));
  INV_X1    g558(.A(G1966), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n472), .A2(G40), .A3(new_n475), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n985), .B1(new_n469), .B2(G2105), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n987), .B1(G164), .B2(G1384), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n498), .A2(new_n500), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n489), .A2(new_n493), .ZN(new_n990));
  AOI211_X1 g565(.A(new_n987), .B(G1384), .C1(new_n989), .C2(new_n990), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n986), .B(new_n988), .C1(new_n991), .C2(KEYINPUT113), .ZN(new_n992));
  AOI21_X1  g567(.A(G1384), .B1(new_n989), .B2(new_n990), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n993), .A2(KEYINPUT113), .A3(KEYINPUT45), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n984), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT118), .ZN(new_n996));
  INV_X1    g571(.A(new_n985), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT65), .ZN(new_n998));
  INV_X1    g573(.A(G125), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n998), .B1(new_n482), .B2(new_n999), .ZN(new_n1000));
  AOI22_X1  g575(.A1(new_n1000), .A2(new_n467), .B1(G113), .B2(G2104), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n997), .B(new_n831), .C1(new_n1001), .C2(new_n471), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT108), .B1(new_n993), .B2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g580(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n993), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1008), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1003), .A2(new_n1005), .A3(new_n1007), .A4(new_n1009), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n995), .A2(new_n996), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n996), .B1(new_n995), .B2(new_n1010), .ZN(new_n1012));
  OAI211_X1 g587(.A(KEYINPUT120), .B(G8), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G8), .ZN(new_n1014));
  NOR2_X1   g589(.A1(G168), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n470), .B(new_n997), .C1(new_n993), .C2(KEYINPUT45), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT113), .B1(new_n993), .B2(KEYINPUT45), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n994), .ZN(new_n1021));
  AOI21_X1  g596(.A(G1966), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1010), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT118), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n995), .A2(new_n996), .A3(new_n1010), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT120), .B1(new_n1026), .B2(G8), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n983), .B1(new_n1017), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1014), .B1(new_n995), .B2(new_n1010), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n1029), .A2(KEYINPUT51), .A3(new_n1015), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1016), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n982), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  AOI211_X1 g610(.A(KEYINPUT121), .B(new_n1033), .C1(new_n1028), .C2(new_n1031), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT62), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(G8), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT120), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1040), .A2(new_n1016), .A3(new_n1013), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1030), .B1(new_n1041), .B2(new_n983), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT121), .B1(new_n1042), .B2(new_n1033), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1032), .A2(new_n982), .A3(new_n1034), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT62), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(G303), .A2(G8), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1047), .B(KEYINPUT55), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n470), .A2(new_n997), .ZN(new_n1049));
  INV_X1    g624(.A(new_n993), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1006), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n993), .A2(new_n1004), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(G2090), .ZN(new_n1055));
  INV_X1    g630(.A(G1971), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n993), .A2(KEYINPUT45), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1057), .A2(new_n988), .A3(new_n986), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1055), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1048), .B1(new_n1059), .B2(new_n1014), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n1047), .B(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1058), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1005), .A2(new_n986), .A3(new_n1007), .A4(new_n1009), .ZN(new_n1064));
  OAI22_X1  g639(.A1(new_n1063), .A2(G1971), .B1(new_n1064), .B2(G2090), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1062), .A2(G8), .A3(new_n1065), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n1060), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(G1981), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1068), .B1(new_n578), .B2(KEYINPUT109), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n718), .B(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT49), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1072), .A2(new_n1014), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1070), .A2(KEYINPUT110), .A3(KEYINPUT49), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT110), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n1069), .B(G305), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT49), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1075), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1071), .B(new_n1073), .C1(new_n1074), .C2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G288), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(G1976), .ZN(new_n1081));
  INV_X1    g656(.A(G1976), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT52), .B1(G288), .B2(new_n1082), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1073), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1073), .A2(new_n1081), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1084), .B1(KEYINPUT52), .B2(new_n1085), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n1079), .A2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1087), .A2(KEYINPUT112), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1079), .A2(new_n1086), .A3(KEYINPUT112), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1067), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT53), .B1(new_n1063), .B2(new_n806), .ZN(new_n1091));
  INV_X1    g666(.A(G1961), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1091), .B1(new_n1092), .B2(new_n1064), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n806), .A2(KEYINPUT53), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(G171), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1090), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1037), .A2(new_n1046), .A3(new_n1098), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1029), .A2(G168), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT63), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1067), .B(new_n1102), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1079), .A2(new_n1082), .A3(new_n1080), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n718), .A2(new_n1068), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT111), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1104), .A2(KEYINPUT111), .A3(new_n1105), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(new_n1109), .A3(new_n1073), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1065), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1048), .B1(new_n1014), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1087), .A2(new_n1100), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1066), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1113), .A2(KEYINPUT63), .B1(new_n1087), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1103), .A2(new_n1110), .A3(new_n1115), .ZN(new_n1116));
  XOR2_X1   g691(.A(G171), .B(KEYINPUT54), .Z(new_n1117));
  OR2_X1    g692(.A1(new_n1001), .A2(KEYINPUT122), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n471), .B1(new_n1001), .B2(KEYINPUT122), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n985), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n1121));
  OR2_X1    g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1057), .A2(new_n988), .ZN(new_n1123));
  AOI211_X1 g698(.A(new_n1095), .B(new_n1123), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1117), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1096), .A2(new_n1117), .B1(new_n1125), .B2(new_n1093), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1067), .B(new_n1126), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1127));
  AOI21_X1  g702(.A(G1956), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1128));
  XOR2_X1   g703(.A(KEYINPUT56), .B(G2072), .Z(new_n1129));
  NOR2_X1   g704(.A1(new_n1058), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT115), .ZN(new_n1132));
  NAND2_X1  g707(.A1(G299), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(KEYINPUT57), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT114), .ZN(new_n1135));
  NAND2_X1  g710(.A1(G299), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(KEYINPUT115), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT57), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1138), .B1(new_n1139), .B2(new_n1137), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1131), .A2(new_n1140), .ZN(new_n1141));
  OAI221_X1 g716(.A(new_n1138), .B1(new_n1139), .B2(new_n1137), .C1(new_n1128), .C2(new_n1130), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1141), .A2(KEYINPUT61), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(G2067), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1072), .A2(new_n1144), .ZN(new_n1145));
  XOR2_X1   g720(.A(new_n1145), .B(KEYINPUT116), .Z(new_n1146));
  NAND2_X1  g721(.A1(new_n1064), .A2(new_n816), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n593), .A2(KEYINPUT60), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g724(.A(KEYINPUT58), .B(G1341), .ZN(new_n1150));
  OAI22_X1  g725(.A1(new_n1072), .A2(new_n1150), .B1(new_n1058), .B2(G1996), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n553), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(KEYINPUT59), .ZN(new_n1153));
  OR2_X1    g728(.A1(new_n1152), .A2(KEYINPUT59), .ZN(new_n1154));
  AND4_X1   g729(.A1(new_n1143), .A2(new_n1149), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1146), .A2(new_n593), .A3(new_n1147), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n593), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1157));
  OAI21_X1  g732(.A(KEYINPUT60), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1159), .A2(KEYINPUT117), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(KEYINPUT117), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1155), .B(new_n1158), .C1(new_n1161), .C2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1142), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1164), .B1(new_n1157), .B2(new_n1141), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1127), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1116), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1099), .A2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1049), .A2(new_n988), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1171), .A2(G1996), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(new_n760), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT105), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n776), .B(new_n1144), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1175), .A2(new_n1171), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1170), .A2(G1996), .A3(new_n759), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT106), .ZN(new_n1178));
  NOR3_X1   g753(.A1(new_n1174), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n739), .A2(new_n741), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n738), .A2(new_n742), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1170), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g758(.A(G290), .B(G1986), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1183), .B1(new_n1170), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1169), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n770), .A2(new_n1144), .A3(new_n775), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1171), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1172), .A2(KEYINPUT46), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1190), .B(KEYINPUT124), .ZN(new_n1191));
  AND2_X1   g766(.A1(new_n1175), .A2(new_n760), .ZN(new_n1192));
  OAI221_X1 g767(.A(new_n1191), .B1(KEYINPUT46), .B2(new_n1172), .C1(new_n1171), .C2(new_n1192), .ZN(new_n1193));
  XOR2_X1   g768(.A(new_n1193), .B(KEYINPUT47), .Z(new_n1194));
  INV_X1    g769(.A(new_n1183), .ZN(new_n1195));
  NOR3_X1   g770(.A1(new_n1171), .A2(G1986), .A3(G290), .ZN(new_n1196));
  XOR2_X1   g771(.A(new_n1196), .B(KEYINPUT48), .Z(new_n1197));
  AOI211_X1 g772(.A(new_n1189), .B(new_n1194), .C1(new_n1195), .C2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1186), .A2(new_n1198), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n1201));
  AOI21_X1  g775(.A(new_n458), .B1(new_n681), .B2(new_n684), .ZN(new_n1202));
  NAND2_X1  g776(.A1(new_n655), .A2(G14), .ZN(new_n1203));
  AOI21_X1  g777(.A(new_n652), .B1(new_n643), .B2(new_n650), .ZN(new_n1204));
  OAI211_X1 g778(.A(KEYINPUT125), .B(new_n1202), .C1(new_n1203), .C2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g779(.A1(new_n1205), .A2(new_n711), .ZN(new_n1206));
  AOI21_X1  g780(.A(KEYINPUT125), .B1(new_n656), .B2(new_n1202), .ZN(new_n1207));
  OAI21_X1  g781(.A(KEYINPUT126), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g782(.A(new_n1202), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1209));
  INV_X1    g783(.A(KEYINPUT125), .ZN(new_n1210));
  NAND2_X1  g784(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n1212));
  NAND4_X1  g786(.A1(new_n1211), .A2(new_n1212), .A3(new_n711), .A4(new_n1205), .ZN(new_n1213));
  NAND2_X1  g787(.A1(new_n1208), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g788(.A1(new_n1214), .A2(new_n886), .ZN(new_n1215));
  INV_X1    g789(.A(new_n1215), .ZN(new_n1216));
  AOI21_X1  g790(.A(new_n1201), .B1(new_n979), .B2(new_n1216), .ZN(new_n1217));
  AOI211_X1 g791(.A(KEYINPUT127), .B(new_n1215), .C1(new_n973), .C2(new_n978), .ZN(new_n1218));
  NOR2_X1   g792(.A1(new_n1217), .A2(new_n1218), .ZN(G308));
  AOI21_X1  g793(.A(new_n965), .B1(new_n950), .B2(new_n952), .ZN(new_n1220));
  NOR3_X1   g794(.A1(new_n956), .A2(new_n964), .A3(KEYINPUT43), .ZN(new_n1221));
  OAI21_X1  g795(.A(new_n1216), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g796(.A1(new_n1222), .A2(KEYINPUT127), .ZN(new_n1223));
  NAND3_X1  g797(.A1(new_n979), .A2(new_n1201), .A3(new_n1216), .ZN(new_n1224));
  NAND2_X1  g798(.A1(new_n1223), .A2(new_n1224), .ZN(G225));
endmodule


