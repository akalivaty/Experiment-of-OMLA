

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U554 ( .A1(n697), .A2(n803), .ZN(n726) );
  NAND2_X1 U555 ( .A1(n730), .A2(n729), .ZN(n751) );
  XNOR2_X1 U556 ( .A(n724), .B(n723), .ZN(n730) );
  INV_X1 U557 ( .A(KEYINPUT29), .ZN(n723) );
  NOR2_X2 U558 ( .A1(G2104), .A2(n534), .ZN(n551) );
  NOR2_X1 U559 ( .A1(n744), .A2(n743), .ZN(n519) );
  INV_X1 U560 ( .A(KEYINPUT98), .ZN(n737) );
  XNOR2_X1 U561 ( .A(n737), .B(KEYINPUT31), .ZN(n738) );
  XNOR2_X1 U562 ( .A(n739), .B(n738), .ZN(n753) );
  INV_X1 U563 ( .A(KEYINPUT102), .ZN(n781) );
  XNOR2_X1 U564 ( .A(KEYINPUT65), .B(G651), .ZN(n524) );
  XNOR2_X1 U565 ( .A(KEYINPUT15), .B(n601), .ZN(n978) );
  NOR2_X1 U566 ( .A1(G651), .A2(n635), .ZN(n657) );
  NOR2_X1 U567 ( .A1(G543), .A2(G651), .ZN(n648) );
  NAND2_X1 U568 ( .A1(n648), .A2(G90), .ZN(n521) );
  XOR2_X1 U569 ( .A(G543), .B(KEYINPUT0), .Z(n635) );
  NOR2_X1 U570 ( .A1(n635), .A2(n524), .ZN(n652) );
  NAND2_X1 U571 ( .A1(G77), .A2(n652), .ZN(n520) );
  NAND2_X1 U572 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U573 ( .A(KEYINPUT9), .B(n522), .ZN(n531) );
  NAND2_X1 U574 ( .A1(G52), .A2(n657), .ZN(n523) );
  XNOR2_X1 U575 ( .A(n523), .B(KEYINPUT69), .ZN(n529) );
  XNOR2_X1 U576 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n526) );
  NOR2_X1 U577 ( .A1(G543), .A2(n524), .ZN(n525) );
  XNOR2_X2 U578 ( .A(n526), .B(n525), .ZN(n649) );
  NAND2_X1 U579 ( .A1(G64), .A2(n649), .ZN(n527) );
  XOR2_X1 U580 ( .A(KEYINPUT68), .B(n527), .Z(n528) );
  NOR2_X1 U581 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U582 ( .A1(n531), .A2(n530), .ZN(G301) );
  INV_X1 U583 ( .A(G301), .ZN(G171) );
  INV_X1 U584 ( .A(G2105), .ZN(n534) );
  AND2_X1 U585 ( .A1(G126), .A2(n551), .ZN(n533) );
  AND2_X1 U586 ( .A1(G2104), .A2(G2105), .ZN(n881) );
  AND2_X1 U587 ( .A1(G114), .A2(n881), .ZN(n532) );
  NOR2_X1 U588 ( .A1(n533), .A2(n532), .ZN(n536) );
  AND2_X1 U589 ( .A1(n534), .A2(G2104), .ZN(n884) );
  NAND2_X1 U590 ( .A1(G102), .A2(n884), .ZN(n535) );
  AND2_X1 U591 ( .A1(n536), .A2(n535), .ZN(n691) );
  NOR2_X1 U592 ( .A1(G2104), .A2(G2105), .ZN(n537) );
  XOR2_X2 U593 ( .A(KEYINPUT17), .B(n537), .Z(n885) );
  NAND2_X1 U594 ( .A1(n885), .A2(G138), .ZN(n538) );
  AND2_X1 U595 ( .A1(n691), .A2(n538), .ZN(G164) );
  XOR2_X1 U596 ( .A(G2443), .B(KEYINPUT106), .Z(n540) );
  XNOR2_X1 U597 ( .A(G2451), .B(G2427), .ZN(n539) );
  XNOR2_X1 U598 ( .A(n540), .B(n539), .ZN(n544) );
  XOR2_X1 U599 ( .A(G2435), .B(G2438), .Z(n542) );
  XNOR2_X1 U600 ( .A(G2454), .B(G2430), .ZN(n541) );
  XNOR2_X1 U601 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U602 ( .A(n544), .B(n543), .Z(n546) );
  XNOR2_X1 U603 ( .A(G2446), .B(KEYINPUT104), .ZN(n545) );
  XNOR2_X1 U604 ( .A(n546), .B(n545), .ZN(n549) );
  XOR2_X1 U605 ( .A(G1348), .B(G1341), .Z(n547) );
  XNOR2_X1 U606 ( .A(KEYINPUT105), .B(n547), .ZN(n548) );
  XOR2_X1 U607 ( .A(n549), .B(n548), .Z(n550) );
  AND2_X1 U608 ( .A1(G14), .A2(n550), .ZN(G401) );
  AND2_X1 U609 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U610 ( .A1(n551), .A2(G123), .ZN(n553) );
  XNOR2_X1 U611 ( .A(KEYINPUT18), .B(KEYINPUT80), .ZN(n552) );
  XNOR2_X1 U612 ( .A(n553), .B(n552), .ZN(n560) );
  NAND2_X1 U613 ( .A1(G99), .A2(n884), .ZN(n555) );
  NAND2_X1 U614 ( .A1(G111), .A2(n881), .ZN(n554) );
  NAND2_X1 U615 ( .A1(n555), .A2(n554), .ZN(n558) );
  NAND2_X1 U616 ( .A1(G135), .A2(n885), .ZN(n556) );
  XNOR2_X1 U617 ( .A(KEYINPUT81), .B(n556), .ZN(n557) );
  NOR2_X1 U618 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U619 ( .A1(n560), .A2(n559), .ZN(n929) );
  XNOR2_X1 U620 ( .A(G2096), .B(n929), .ZN(n561) );
  OR2_X1 U621 ( .A1(G2100), .A2(n561), .ZN(G156) );
  INV_X1 U622 ( .A(G57), .ZN(G237) );
  INV_X1 U623 ( .A(G132), .ZN(G219) );
  INV_X1 U624 ( .A(G82), .ZN(G220) );
  NAND2_X1 U625 ( .A1(G50), .A2(n657), .ZN(n563) );
  NAND2_X1 U626 ( .A1(G62), .A2(n649), .ZN(n562) );
  NAND2_X1 U627 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U628 ( .A(KEYINPUT86), .B(n564), .Z(n568) );
  NAND2_X1 U629 ( .A1(n652), .A2(G75), .ZN(n566) );
  NAND2_X1 U630 ( .A1(n648), .A2(G88), .ZN(n565) );
  AND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n568), .A2(n567), .ZN(G303) );
  NAND2_X1 U633 ( .A1(G51), .A2(n657), .ZN(n570) );
  NAND2_X1 U634 ( .A1(G63), .A2(n649), .ZN(n569) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(KEYINPUT6), .B(n571), .ZN(n577) );
  NAND2_X1 U637 ( .A1(n648), .A2(G89), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(KEYINPUT4), .ZN(n574) );
  NAND2_X1 U639 ( .A1(G76), .A2(n652), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U641 ( .A(n575), .B(KEYINPUT5), .Z(n576) );
  NOR2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U643 ( .A(KEYINPUT76), .B(n578), .Z(n579) );
  XNOR2_X1 U644 ( .A(KEYINPUT7), .B(n579), .ZN(G168) );
  XOR2_X1 U645 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U646 ( .A1(G7), .A2(G661), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n580), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U648 ( .A(G223), .ZN(n835) );
  NAND2_X1 U649 ( .A1(n835), .A2(G567), .ZN(n581) );
  XNOR2_X1 U650 ( .A(n581), .B(KEYINPUT71), .ZN(n582) );
  XNOR2_X1 U651 ( .A(KEYINPUT11), .B(n582), .ZN(G234) );
  NAND2_X1 U652 ( .A1(n648), .A2(G81), .ZN(n583) );
  XNOR2_X1 U653 ( .A(n583), .B(KEYINPUT12), .ZN(n585) );
  NAND2_X1 U654 ( .A1(G68), .A2(n652), .ZN(n584) );
  NAND2_X1 U655 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U656 ( .A(n586), .B(KEYINPUT13), .ZN(n588) );
  NAND2_X1 U657 ( .A1(G43), .A2(n657), .ZN(n587) );
  NAND2_X1 U658 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U659 ( .A1(n649), .A2(G56), .ZN(n589) );
  XOR2_X1 U660 ( .A(KEYINPUT14), .B(n589), .Z(n590) );
  NOR2_X1 U661 ( .A1(n591), .A2(n590), .ZN(n990) );
  XOR2_X1 U662 ( .A(G860), .B(KEYINPUT72), .Z(n613) );
  INV_X1 U663 ( .A(n613), .ZN(n592) );
  NAND2_X1 U664 ( .A1(n990), .A2(n592), .ZN(G153) );
  NAND2_X1 U665 ( .A1(G54), .A2(n657), .ZN(n593) );
  XNOR2_X1 U666 ( .A(n593), .B(KEYINPUT74), .ZN(n600) );
  NAND2_X1 U667 ( .A1(n648), .A2(G92), .ZN(n595) );
  NAND2_X1 U668 ( .A1(G79), .A2(n652), .ZN(n594) );
  NAND2_X1 U669 ( .A1(n595), .A2(n594), .ZN(n598) );
  NAND2_X1 U670 ( .A1(G66), .A2(n649), .ZN(n596) );
  XNOR2_X1 U671 ( .A(KEYINPUT73), .B(n596), .ZN(n597) );
  NOR2_X1 U672 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U673 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U674 ( .A1(n978), .A2(G868), .ZN(n602) );
  XNOR2_X1 U675 ( .A(n602), .B(KEYINPUT75), .ZN(n604) );
  NAND2_X1 U676 ( .A1(G868), .A2(G301), .ZN(n603) );
  NAND2_X1 U677 ( .A1(n604), .A2(n603), .ZN(G284) );
  NAND2_X1 U678 ( .A1(G53), .A2(n657), .ZN(n606) );
  NAND2_X1 U679 ( .A1(G65), .A2(n649), .ZN(n605) );
  NAND2_X1 U680 ( .A1(n606), .A2(n605), .ZN(n610) );
  NAND2_X1 U681 ( .A1(n648), .A2(G91), .ZN(n608) );
  NAND2_X1 U682 ( .A1(G78), .A2(n652), .ZN(n607) );
  NAND2_X1 U683 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U684 ( .A1(n610), .A2(n609), .ZN(n969) );
  XOR2_X1 U685 ( .A(KEYINPUT70), .B(n969), .Z(G299) );
  NAND2_X1 U686 ( .A1(G868), .A2(G286), .ZN(n612) );
  INV_X1 U687 ( .A(G868), .ZN(n620) );
  NAND2_X1 U688 ( .A1(G299), .A2(n620), .ZN(n611) );
  NAND2_X1 U689 ( .A1(n612), .A2(n611), .ZN(G297) );
  NAND2_X1 U690 ( .A1(n613), .A2(G559), .ZN(n614) );
  NAND2_X1 U691 ( .A1(n614), .A2(n978), .ZN(n615) );
  XNOR2_X1 U692 ( .A(n615), .B(KEYINPUT16), .ZN(n616) );
  XOR2_X1 U693 ( .A(KEYINPUT77), .B(n616), .Z(G148) );
  INV_X1 U694 ( .A(n978), .ZN(n617) );
  NOR2_X1 U695 ( .A1(G559), .A2(n617), .ZN(n618) );
  NAND2_X1 U696 ( .A1(G868), .A2(n618), .ZN(n619) );
  XNOR2_X1 U697 ( .A(n619), .B(KEYINPUT78), .ZN(n622) );
  NAND2_X1 U698 ( .A1(n990), .A2(n620), .ZN(n621) );
  NAND2_X1 U699 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U700 ( .A(KEYINPUT79), .B(n623), .ZN(G282) );
  NAND2_X1 U701 ( .A1(G559), .A2(n978), .ZN(n624) );
  XOR2_X1 U702 ( .A(n990), .B(n624), .Z(n667) );
  NOR2_X1 U703 ( .A1(G860), .A2(n667), .ZN(n634) );
  NAND2_X1 U704 ( .A1(n648), .A2(G93), .ZN(n626) );
  NAND2_X1 U705 ( .A1(G80), .A2(n652), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U707 ( .A(n627), .B(KEYINPUT83), .ZN(n629) );
  NAND2_X1 U708 ( .A1(G55), .A2(n657), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n649), .A2(G67), .ZN(n630) );
  XOR2_X1 U711 ( .A(KEYINPUT84), .B(n630), .Z(n631) );
  NOR2_X1 U712 ( .A1(n632), .A2(n631), .ZN(n661) );
  XNOR2_X1 U713 ( .A(n661), .B(KEYINPUT82), .ZN(n633) );
  XNOR2_X1 U714 ( .A(n634), .B(n633), .ZN(G145) );
  NAND2_X1 U715 ( .A1(G87), .A2(n635), .ZN(n637) );
  NAND2_X1 U716 ( .A1(G74), .A2(G651), .ZN(n636) );
  NAND2_X1 U717 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U718 ( .A1(n649), .A2(n638), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n657), .A2(G49), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n640), .A2(n639), .ZN(G288) );
  NAND2_X1 U721 ( .A1(n648), .A2(G85), .ZN(n642) );
  NAND2_X1 U722 ( .A1(G72), .A2(n652), .ZN(n641) );
  NAND2_X1 U723 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U724 ( .A(KEYINPUT66), .B(n643), .Z(n647) );
  NAND2_X1 U725 ( .A1(n649), .A2(G60), .ZN(n645) );
  NAND2_X1 U726 ( .A1(G47), .A2(n657), .ZN(n644) );
  AND2_X1 U727 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U728 ( .A1(n647), .A2(n646), .ZN(G290) );
  NAND2_X1 U729 ( .A1(n648), .A2(G86), .ZN(n651) );
  NAND2_X1 U730 ( .A1(G61), .A2(n649), .ZN(n650) );
  NAND2_X1 U731 ( .A1(n651), .A2(n650), .ZN(n655) );
  NAND2_X1 U732 ( .A1(G73), .A2(n652), .ZN(n653) );
  XOR2_X1 U733 ( .A(KEYINPUT2), .B(n653), .Z(n654) );
  NOR2_X1 U734 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U735 ( .A(KEYINPUT85), .B(n656), .Z(n659) );
  NAND2_X1 U736 ( .A1(n657), .A2(G48), .ZN(n658) );
  NAND2_X1 U737 ( .A1(n659), .A2(n658), .ZN(G305) );
  NOR2_X1 U738 ( .A1(G868), .A2(n661), .ZN(n660) );
  XNOR2_X1 U739 ( .A(n660), .B(KEYINPUT87), .ZN(n670) );
  XNOR2_X1 U740 ( .A(KEYINPUT19), .B(G299), .ZN(n663) );
  XNOR2_X1 U741 ( .A(G288), .B(n661), .ZN(n662) );
  XNOR2_X1 U742 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U743 ( .A(n664), .B(G290), .ZN(n665) );
  XNOR2_X1 U744 ( .A(n665), .B(G303), .ZN(n666) );
  XNOR2_X1 U745 ( .A(n666), .B(G305), .ZN(n905) );
  XNOR2_X1 U746 ( .A(n905), .B(n667), .ZN(n668) );
  NAND2_X1 U747 ( .A1(G868), .A2(n668), .ZN(n669) );
  NAND2_X1 U748 ( .A1(n670), .A2(n669), .ZN(G295) );
  NAND2_X1 U749 ( .A1(G2084), .A2(G2078), .ZN(n671) );
  XOR2_X1 U750 ( .A(KEYINPUT20), .B(n671), .Z(n672) );
  NAND2_X1 U751 ( .A1(G2090), .A2(n672), .ZN(n674) );
  XNOR2_X1 U752 ( .A(KEYINPUT88), .B(KEYINPUT21), .ZN(n673) );
  XNOR2_X1 U753 ( .A(n674), .B(n673), .ZN(n675) );
  NAND2_X1 U754 ( .A1(G2072), .A2(n675), .ZN(G158) );
  XNOR2_X1 U755 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U756 ( .A1(G220), .A2(G219), .ZN(n676) );
  XOR2_X1 U757 ( .A(KEYINPUT22), .B(n676), .Z(n677) );
  NOR2_X1 U758 ( .A1(G218), .A2(n677), .ZN(n678) );
  NAND2_X1 U759 ( .A1(G96), .A2(n678), .ZN(n842) );
  NAND2_X1 U760 ( .A1(G2106), .A2(n842), .ZN(n682) );
  NAND2_X1 U761 ( .A1(G69), .A2(G120), .ZN(n679) );
  NOR2_X1 U762 ( .A1(G237), .A2(n679), .ZN(n680) );
  NAND2_X1 U763 ( .A1(G108), .A2(n680), .ZN(n843) );
  NAND2_X1 U764 ( .A1(G567), .A2(n843), .ZN(n681) );
  NAND2_X1 U765 ( .A1(n682), .A2(n681), .ZN(n844) );
  NAND2_X1 U766 ( .A1(G483), .A2(G661), .ZN(n683) );
  NOR2_X1 U767 ( .A1(n844), .A2(n683), .ZN(n839) );
  NAND2_X1 U768 ( .A1(n839), .A2(G36), .ZN(G176) );
  NAND2_X1 U769 ( .A1(n881), .A2(G113), .ZN(n686) );
  NAND2_X1 U770 ( .A1(G101), .A2(n884), .ZN(n684) );
  XOR2_X1 U771 ( .A(KEYINPUT23), .B(n684), .Z(n685) );
  NAND2_X1 U772 ( .A1(n686), .A2(n685), .ZN(n690) );
  NAND2_X1 U773 ( .A1(G137), .A2(n885), .ZN(n688) );
  NAND2_X1 U774 ( .A1(G125), .A2(n551), .ZN(n687) );
  NAND2_X1 U775 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U776 ( .A1(n690), .A2(n689), .ZN(G160) );
  INV_X1 U777 ( .A(G303), .ZN(G166) );
  OR2_X1 U778 ( .A1(n691), .A2(G1384), .ZN(n695) );
  INV_X1 U779 ( .A(G1384), .ZN(n692) );
  AND2_X1 U780 ( .A1(G138), .A2(n692), .ZN(n693) );
  NAND2_X1 U781 ( .A1(n885), .A2(n693), .ZN(n694) );
  NAND2_X1 U782 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U783 ( .A(n696), .B(KEYINPUT64), .ZN(n802) );
  INV_X1 U784 ( .A(n802), .ZN(n697) );
  NAND2_X1 U785 ( .A1(G160), .A2(G40), .ZN(n803) );
  INV_X1 U786 ( .A(n726), .ZN(n746) );
  NAND2_X1 U787 ( .A1(G8), .A2(n746), .ZN(n775) );
  NOR2_X1 U788 ( .A1(G1981), .A2(G305), .ZN(n698) );
  XOR2_X1 U789 ( .A(n698), .B(KEYINPUT24), .Z(n699) );
  NOR2_X1 U790 ( .A1(n775), .A2(n699), .ZN(n780) );
  NAND2_X1 U791 ( .A1(G1996), .A2(n726), .ZN(n700) );
  XNOR2_X1 U792 ( .A(KEYINPUT26), .B(n700), .ZN(n701) );
  NAND2_X1 U793 ( .A1(n701), .A2(n990), .ZN(n704) );
  NAND2_X1 U794 ( .A1(G1341), .A2(n746), .ZN(n702) );
  XNOR2_X1 U795 ( .A(KEYINPUT95), .B(n702), .ZN(n703) );
  NOR2_X1 U796 ( .A1(n704), .A2(n703), .ZN(n710) );
  NAND2_X1 U797 ( .A1(n978), .A2(n710), .ZN(n709) );
  NAND2_X1 U798 ( .A1(n746), .A2(G1348), .ZN(n705) );
  XNOR2_X1 U799 ( .A(n705), .B(KEYINPUT96), .ZN(n707) );
  NAND2_X1 U800 ( .A1(n726), .A2(G2067), .ZN(n706) );
  NAND2_X1 U801 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U802 ( .A1(n709), .A2(n708), .ZN(n712) );
  OR2_X1 U803 ( .A1(n978), .A2(n710), .ZN(n711) );
  NAND2_X1 U804 ( .A1(n712), .A2(n711), .ZN(n718) );
  NAND2_X1 U805 ( .A1(n726), .A2(G2072), .ZN(n713) );
  XNOR2_X1 U806 ( .A(n713), .B(KEYINPUT27), .ZN(n715) );
  INV_X1 U807 ( .A(G1956), .ZN(n998) );
  NOR2_X1 U808 ( .A1(n998), .A2(n726), .ZN(n714) );
  NOR2_X1 U809 ( .A1(n715), .A2(n714), .ZN(n719) );
  AND2_X1 U810 ( .A1(n969), .A2(n719), .ZN(n716) );
  XNOR2_X1 U811 ( .A(KEYINPUT97), .B(n716), .ZN(n717) );
  NAND2_X1 U812 ( .A1(n718), .A2(n717), .ZN(n722) );
  NOR2_X1 U813 ( .A1(n969), .A2(n719), .ZN(n720) );
  XOR2_X1 U814 ( .A(KEYINPUT28), .B(n720), .Z(n721) );
  NAND2_X1 U815 ( .A1(n722), .A2(n721), .ZN(n724) );
  XNOR2_X1 U816 ( .A(G2078), .B(KEYINPUT25), .ZN(n945) );
  NAND2_X1 U817 ( .A1(n726), .A2(n945), .ZN(n725) );
  XNOR2_X1 U818 ( .A(n725), .B(KEYINPUT94), .ZN(n728) );
  OR2_X1 U819 ( .A1(G1961), .A2(n726), .ZN(n727) );
  NAND2_X1 U820 ( .A1(n728), .A2(n727), .ZN(n731) );
  NAND2_X1 U821 ( .A1(n731), .A2(G171), .ZN(n729) );
  NOR2_X1 U822 ( .A1(G171), .A2(n731), .ZN(n736) );
  NOR2_X1 U823 ( .A1(G1966), .A2(n775), .ZN(n744) );
  NOR2_X1 U824 ( .A1(n746), .A2(G2084), .ZN(n742) );
  NOR2_X1 U825 ( .A1(n744), .A2(n742), .ZN(n732) );
  NAND2_X1 U826 ( .A1(G8), .A2(n732), .ZN(n733) );
  XNOR2_X1 U827 ( .A(n733), .B(KEYINPUT30), .ZN(n734) );
  NOR2_X1 U828 ( .A1(n734), .A2(G168), .ZN(n735) );
  NOR2_X1 U829 ( .A1(n736), .A2(n735), .ZN(n739) );
  NAND2_X1 U830 ( .A1(n751), .A2(n753), .ZN(n741) );
  INV_X1 U831 ( .A(KEYINPUT99), .ZN(n740) );
  XNOR2_X1 U832 ( .A(n741), .B(n740), .ZN(n745) );
  AND2_X1 U833 ( .A1(n742), .A2(G8), .ZN(n743) );
  AND2_X1 U834 ( .A1(n745), .A2(n519), .ZN(n761) );
  NOR2_X1 U835 ( .A1(G1971), .A2(n775), .ZN(n748) );
  NOR2_X1 U836 ( .A1(G2090), .A2(n746), .ZN(n747) );
  NOR2_X1 U837 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U838 ( .A1(n749), .A2(G303), .ZN(n750) );
  XNOR2_X1 U839 ( .A(n750), .B(KEYINPUT100), .ZN(n754) );
  AND2_X1 U840 ( .A1(n751), .A2(n754), .ZN(n752) );
  NAND2_X1 U841 ( .A1(n753), .A2(n752), .ZN(n758) );
  INV_X1 U842 ( .A(n754), .ZN(n755) );
  OR2_X1 U843 ( .A1(n755), .A2(G286), .ZN(n756) );
  AND2_X1 U844 ( .A1(G8), .A2(n756), .ZN(n757) );
  NAND2_X1 U845 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U846 ( .A(KEYINPUT32), .B(n759), .Z(n760) );
  OR2_X2 U847 ( .A1(n761), .A2(n760), .ZN(n770) );
  NOR2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n970) );
  NOR2_X1 U849 ( .A1(G1971), .A2(G303), .ZN(n975) );
  NOR2_X1 U850 ( .A1(n970), .A2(n975), .ZN(n762) );
  NAND2_X1 U851 ( .A1(n770), .A2(n762), .ZN(n763) );
  NAND2_X1 U852 ( .A1(G1976), .A2(G288), .ZN(n972) );
  NAND2_X1 U853 ( .A1(n763), .A2(n972), .ZN(n764) );
  NOR2_X1 U854 ( .A1(n775), .A2(n764), .ZN(n765) );
  NOR2_X1 U855 ( .A1(KEYINPUT33), .A2(n765), .ZN(n768) );
  NAND2_X1 U856 ( .A1(n970), .A2(KEYINPUT33), .ZN(n766) );
  NOR2_X1 U857 ( .A1(n766), .A2(n775), .ZN(n767) );
  NOR2_X1 U858 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U859 ( .A(G1981), .B(G305), .Z(n986) );
  NAND2_X1 U860 ( .A1(n769), .A2(n986), .ZN(n778) );
  INV_X1 U861 ( .A(n770), .ZN(n773) );
  NAND2_X1 U862 ( .A1(G166), .A2(G8), .ZN(n771) );
  NOR2_X1 U863 ( .A1(G2090), .A2(n771), .ZN(n772) );
  NOR2_X1 U864 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U865 ( .A(n774), .B(KEYINPUT101), .ZN(n776) );
  NAND2_X1 U866 ( .A1(n776), .A2(n775), .ZN(n777) );
  NAND2_X1 U867 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n782) );
  XNOR2_X1 U869 ( .A(n782), .B(n781), .ZN(n818) );
  NAND2_X1 U870 ( .A1(G95), .A2(n884), .ZN(n784) );
  NAND2_X1 U871 ( .A1(G107), .A2(n881), .ZN(n783) );
  NAND2_X1 U872 ( .A1(n784), .A2(n783), .ZN(n787) );
  NAND2_X1 U873 ( .A1(n885), .A2(G131), .ZN(n785) );
  XOR2_X1 U874 ( .A(KEYINPUT92), .B(n785), .Z(n786) );
  NOR2_X1 U875 ( .A1(n787), .A2(n786), .ZN(n789) );
  NAND2_X1 U876 ( .A1(n551), .A2(G119), .ZN(n788) );
  NAND2_X1 U877 ( .A1(n789), .A2(n788), .ZN(n878) );
  NAND2_X1 U878 ( .A1(n878), .A2(G1991), .ZN(n799) );
  NAND2_X1 U879 ( .A1(G129), .A2(n551), .ZN(n791) );
  NAND2_X1 U880 ( .A1(G117), .A2(n881), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n791), .A2(n790), .ZN(n794) );
  NAND2_X1 U882 ( .A1(n884), .A2(G105), .ZN(n792) );
  XOR2_X1 U883 ( .A(KEYINPUT38), .B(n792), .Z(n793) );
  NOR2_X1 U884 ( .A1(n794), .A2(n793), .ZN(n795) );
  XOR2_X1 U885 ( .A(KEYINPUT93), .B(n795), .Z(n797) );
  NAND2_X1 U886 ( .A1(n885), .A2(G141), .ZN(n796) );
  NAND2_X1 U887 ( .A1(n797), .A2(n796), .ZN(n879) );
  NAND2_X1 U888 ( .A1(n879), .A2(G1996), .ZN(n798) );
  NAND2_X1 U889 ( .A1(n799), .A2(n798), .ZN(n916) );
  INV_X1 U890 ( .A(n916), .ZN(n801) );
  XNOR2_X1 U891 ( .A(KEYINPUT89), .B(G1986), .ZN(n800) );
  XNOR2_X1 U892 ( .A(n800), .B(G290), .ZN(n982) );
  NAND2_X1 U893 ( .A1(n801), .A2(n982), .ZN(n804) );
  NOR2_X1 U894 ( .A1(n803), .A2(n802), .ZN(n829) );
  NAND2_X1 U895 ( .A1(n804), .A2(n829), .ZN(n816) );
  NAND2_X1 U896 ( .A1(n884), .A2(G104), .ZN(n805) );
  XNOR2_X1 U897 ( .A(n805), .B(KEYINPUT90), .ZN(n807) );
  NAND2_X1 U898 ( .A1(G140), .A2(n885), .ZN(n806) );
  NAND2_X1 U899 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U900 ( .A(KEYINPUT34), .B(n808), .ZN(n814) );
  NAND2_X1 U901 ( .A1(G128), .A2(n551), .ZN(n810) );
  NAND2_X1 U902 ( .A1(G116), .A2(n881), .ZN(n809) );
  NAND2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U904 ( .A(KEYINPUT35), .B(n811), .ZN(n812) );
  XNOR2_X1 U905 ( .A(KEYINPUT91), .B(n812), .ZN(n813) );
  NOR2_X1 U906 ( .A1(n814), .A2(n813), .ZN(n815) );
  XOR2_X1 U907 ( .A(KEYINPUT36), .B(n815), .Z(n901) );
  XOR2_X1 U908 ( .A(G2067), .B(KEYINPUT37), .Z(n828) );
  AND2_X1 U909 ( .A1(n901), .A2(n828), .ZN(n923) );
  NAND2_X1 U910 ( .A1(n923), .A2(n829), .ZN(n819) );
  AND2_X1 U911 ( .A1(n816), .A2(n819), .ZN(n817) );
  NAND2_X1 U912 ( .A1(n818), .A2(n817), .ZN(n833) );
  INV_X1 U913 ( .A(n819), .ZN(n827) );
  NOR2_X1 U914 ( .A1(G1996), .A2(n879), .ZN(n927) );
  NOR2_X1 U915 ( .A1(G1986), .A2(G290), .ZN(n821) );
  NOR2_X1 U916 ( .A1(G1991), .A2(n878), .ZN(n820) );
  XOR2_X1 U917 ( .A(KEYINPUT103), .B(n820), .Z(n932) );
  NOR2_X1 U918 ( .A1(n821), .A2(n932), .ZN(n822) );
  NOR2_X1 U919 ( .A1(n916), .A2(n822), .ZN(n823) );
  NOR2_X1 U920 ( .A1(n927), .A2(n823), .ZN(n824) );
  XNOR2_X1 U921 ( .A(KEYINPUT39), .B(n824), .ZN(n825) );
  NAND2_X1 U922 ( .A1(n825), .A2(n829), .ZN(n826) );
  OR2_X1 U923 ( .A1(n827), .A2(n826), .ZN(n831) );
  NOR2_X1 U924 ( .A1(n901), .A2(n828), .ZN(n917) );
  NAND2_X1 U925 ( .A1(n917), .A2(n829), .ZN(n830) );
  AND2_X1 U926 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U927 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U928 ( .A(n834), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n835), .ZN(G217) );
  NAND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n837) );
  INV_X1 U931 ( .A(G661), .ZN(n836) );
  NOR2_X1 U932 ( .A1(n837), .A2(n836), .ZN(n838) );
  XNOR2_X1 U933 ( .A(n838), .B(KEYINPUT107), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G1), .A2(G3), .ZN(n840) );
  NAND2_X1 U935 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U936 ( .A(n841), .B(KEYINPUT108), .ZN(G188) );
  INV_X1 U938 ( .A(G120), .ZN(G236) );
  INV_X1 U939 ( .A(G96), .ZN(G221) );
  INV_X1 U940 ( .A(G69), .ZN(G235) );
  NOR2_X1 U941 ( .A1(n843), .A2(n842), .ZN(G325) );
  INV_X1 U942 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U943 ( .A(KEYINPUT109), .B(n844), .ZN(G319) );
  XOR2_X1 U944 ( .A(G2100), .B(G2096), .Z(n846) );
  XNOR2_X1 U945 ( .A(KEYINPUT42), .B(G2678), .ZN(n845) );
  XNOR2_X1 U946 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U947 ( .A(KEYINPUT43), .B(G2090), .Z(n848) );
  XNOR2_X1 U948 ( .A(G2067), .B(G2072), .ZN(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U950 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U951 ( .A(G2084), .B(G2078), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n852), .B(n851), .ZN(G227) );
  XOR2_X1 U953 ( .A(KEYINPUT41), .B(G1981), .Z(n854) );
  XNOR2_X1 U954 ( .A(G1966), .B(G1971), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U956 ( .A(n855), .B(KEYINPUT110), .Z(n857) );
  XNOR2_X1 U957 ( .A(G1991), .B(G1996), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U959 ( .A(G1976), .B(G1956), .Z(n859) );
  XNOR2_X1 U960 ( .A(G1986), .B(G1961), .ZN(n858) );
  XNOR2_X1 U961 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U962 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U963 ( .A(KEYINPUT111), .B(G2474), .ZN(n862) );
  XNOR2_X1 U964 ( .A(n863), .B(n862), .ZN(G229) );
  NAND2_X1 U965 ( .A1(n551), .A2(G124), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n864), .B(KEYINPUT44), .ZN(n866) );
  NAND2_X1 U967 ( .A1(G112), .A2(n881), .ZN(n865) );
  NAND2_X1 U968 ( .A1(n866), .A2(n865), .ZN(n870) );
  NAND2_X1 U969 ( .A1(G100), .A2(n884), .ZN(n868) );
  NAND2_X1 U970 ( .A1(G136), .A2(n885), .ZN(n867) );
  NAND2_X1 U971 ( .A1(n868), .A2(n867), .ZN(n869) );
  NOR2_X1 U972 ( .A1(n870), .A2(n869), .ZN(G162) );
  NAND2_X1 U973 ( .A1(G103), .A2(n884), .ZN(n872) );
  NAND2_X1 U974 ( .A1(G139), .A2(n885), .ZN(n871) );
  NAND2_X1 U975 ( .A1(n872), .A2(n871), .ZN(n877) );
  NAND2_X1 U976 ( .A1(G127), .A2(n551), .ZN(n874) );
  NAND2_X1 U977 ( .A1(G115), .A2(n881), .ZN(n873) );
  NAND2_X1 U978 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U979 ( .A(KEYINPUT47), .B(n875), .Z(n876) );
  NOR2_X1 U980 ( .A1(n877), .A2(n876), .ZN(n918) );
  XNOR2_X1 U981 ( .A(n918), .B(n878), .ZN(n880) );
  XNOR2_X1 U982 ( .A(n880), .B(n879), .ZN(n892) );
  NAND2_X1 U983 ( .A1(G130), .A2(n551), .ZN(n883) );
  NAND2_X1 U984 ( .A1(G118), .A2(n881), .ZN(n882) );
  NAND2_X1 U985 ( .A1(n883), .A2(n882), .ZN(n890) );
  NAND2_X1 U986 ( .A1(G106), .A2(n884), .ZN(n887) );
  NAND2_X1 U987 ( .A1(G142), .A2(n885), .ZN(n886) );
  NAND2_X1 U988 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U989 ( .A(KEYINPUT45), .B(n888), .Z(n889) );
  NOR2_X1 U990 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U991 ( .A(n892), .B(n891), .Z(n894) );
  XNOR2_X1 U992 ( .A(G160), .B(G162), .ZN(n893) );
  XNOR2_X1 U993 ( .A(n894), .B(n893), .ZN(n903) );
  XNOR2_X1 U994 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n929), .B(KEYINPUT46), .ZN(n895) );
  XNOR2_X1 U996 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U997 ( .A(n897), .B(KEYINPUT112), .Z(n899) );
  XNOR2_X1 U998 ( .A(G164), .B(KEYINPUT48), .ZN(n898) );
  XNOR2_X1 U999 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U1000 ( .A(n901), .B(n900), .Z(n902) );
  XNOR2_X1 U1001 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n904), .ZN(G395) );
  XNOR2_X1 U1003 ( .A(G286), .B(n905), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(G171), .B(n990), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n908), .B(n978), .ZN(n909) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n909), .ZN(G397) );
  NOR2_X1 U1008 ( .A1(G227), .A2(G229), .ZN(n910) );
  XOR2_X1 U1009 ( .A(KEYINPUT49), .B(n910), .Z(n911) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n911), .ZN(n912) );
  NOR2_X1 U1011 ( .A1(G401), .A2(n912), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n913) );
  XOR2_X1 U1013 ( .A(KEYINPUT115), .B(n913), .Z(n914) );
  NAND2_X1 U1014 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(G108), .ZN(G238) );
  NOR2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n925) );
  XOR2_X1 U1018 ( .A(G2072), .B(n918), .Z(n920) );
  XOR2_X1 U1019 ( .A(G164), .B(G2078), .Z(n919) );
  NOR2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1021 ( .A(KEYINPUT50), .B(n921), .Z(n922) );
  NOR2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n937) );
  XOR2_X1 U1024 ( .A(G2090), .B(G162), .Z(n926) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1026 ( .A(KEYINPUT51), .B(n928), .Z(n935) );
  XNOR2_X1 U1027 ( .A(G160), .B(G2084), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1030 ( .A(n933), .B(KEYINPUT116), .ZN(n934) );
  NAND2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1033 ( .A(KEYINPUT52), .B(n938), .ZN(n939) );
  INV_X1 U1034 ( .A(KEYINPUT55), .ZN(n962) );
  NAND2_X1 U1035 ( .A1(n939), .A2(n962), .ZN(n940) );
  NAND2_X1 U1036 ( .A1(n940), .A2(G29), .ZN(n1027) );
  XNOR2_X1 U1037 ( .A(KEYINPUT117), .B(G2090), .ZN(n941) );
  XNOR2_X1 U1038 ( .A(n941), .B(G35), .ZN(n960) );
  XNOR2_X1 U1039 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n955) );
  XNOR2_X1 U1040 ( .A(G2067), .B(G26), .ZN(n943) );
  XNOR2_X1 U1041 ( .A(G33), .B(G2072), .ZN(n942) );
  NOR2_X1 U1042 ( .A1(n943), .A2(n942), .ZN(n952) );
  XOR2_X1 U1043 ( .A(G1991), .B(G25), .Z(n944) );
  NAND2_X1 U1044 ( .A1(n944), .A2(G28), .ZN(n950) );
  XOR2_X1 U1045 ( .A(G1996), .B(G32), .Z(n947) );
  XNOR2_X1 U1046 ( .A(n945), .B(G27), .ZN(n946) );
  NAND2_X1 U1047 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1048 ( .A(KEYINPUT118), .B(n948), .ZN(n949) );
  NOR2_X1 U1049 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1050 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1051 ( .A(KEYINPUT53), .B(n953), .ZN(n954) );
  XNOR2_X1 U1052 ( .A(n955), .B(n954), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(G2084), .B(G34), .ZN(n956) );
  XNOR2_X1 U1054 ( .A(KEYINPUT54), .B(n956), .ZN(n957) );
  NOR2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(n962), .B(n961), .ZN(n964) );
  INV_X1 U1058 ( .A(G29), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1060 ( .A1(G11), .A2(n965), .ZN(n1025) );
  INV_X1 U1061 ( .A(G16), .ZN(n1021) );
  XNOR2_X1 U1062 ( .A(KEYINPUT56), .B(KEYINPUT121), .ZN(n966) );
  XNOR2_X1 U1063 ( .A(n1021), .B(n966), .ZN(n997) );
  XNOR2_X1 U1064 ( .A(G171), .B(G1961), .ZN(n968) );
  NAND2_X1 U1065 ( .A1(G1971), .A2(G303), .ZN(n967) );
  NAND2_X1 U1066 ( .A1(n968), .A2(n967), .ZN(n984) );
  XNOR2_X1 U1067 ( .A(n969), .B(G1956), .ZN(n977) );
  INV_X1 U1068 ( .A(n970), .ZN(n971) );
  NAND2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1070 ( .A(KEYINPUT123), .B(n973), .Z(n974) );
  NOR2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n980) );
  XOR2_X1 U1073 ( .A(G1348), .B(n978), .Z(n979) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(KEYINPUT124), .B(n985), .ZN(n995) );
  XNOR2_X1 U1078 ( .A(G1966), .B(G168), .ZN(n987) );
  NAND2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n989) );
  XOR2_X1 U1080 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n988) );
  XNOR2_X1 U1081 ( .A(n989), .B(n988), .ZN(n993) );
  XNOR2_X1 U1082 ( .A(n990), .B(G1341), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(KEYINPUT125), .B(n991), .ZN(n992) );
  NOR2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n1023) );
  XNOR2_X1 U1087 ( .A(G20), .B(n998), .ZN(n1002) );
  XNOR2_X1 U1088 ( .A(G1341), .B(G19), .ZN(n1000) );
  XNOR2_X1 U1089 ( .A(G6), .B(G1981), .ZN(n999) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XOR2_X1 U1092 ( .A(KEYINPUT59), .B(G1348), .Z(n1003) );
  XNOR2_X1 U1093 ( .A(G4), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(KEYINPUT60), .B(n1006), .ZN(n1016) );
  XNOR2_X1 U1096 ( .A(G1961), .B(KEYINPUT126), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(n1007), .B(G5), .ZN(n1014) );
  XNOR2_X1 U1098 ( .A(G1971), .B(G22), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(G23), .B(G1976), .ZN(n1008) );
  NOR2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  XOR2_X1 U1101 ( .A(G1986), .B(G24), .Z(n1010) );
  NAND2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1103 ( .A(KEYINPUT58), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(G21), .B(G1966), .ZN(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1108 ( .A(KEYINPUT61), .B(n1019), .ZN(n1020) );
  NAND2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1113 ( .A(n1028), .B(KEYINPUT127), .ZN(n1029) );
  XNOR2_X1 U1114 ( .A(KEYINPUT62), .B(n1029), .ZN(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

