

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U554 ( .A(n731), .ZN(n705) );
  NAND2_X2 U555 ( .A1(n780), .A2(n782), .ZN(n731) );
  XOR2_X1 U556 ( .A(KEYINPUT17), .B(n531), .Z(n870) );
  XNOR2_X1 U557 ( .A(n681), .B(KEYINPUT83), .ZN(n780) );
  OR2_X1 U558 ( .A1(n968), .A2(n753), .ZN(n522) );
  NAND2_X1 U559 ( .A1(n750), .A2(n749), .ZN(n523) );
  AND2_X1 U560 ( .A1(n685), .A2(n684), .ZN(n524) );
  OR2_X1 U561 ( .A1(n761), .A2(n760), .ZN(n525) );
  XOR2_X1 U562 ( .A(n747), .B(KEYINPUT96), .Z(n526) );
  NOR2_X1 U563 ( .A1(n752), .A2(n751), .ZN(n527) );
  INV_X1 U564 ( .A(n982), .ZN(n684) );
  AND2_X1 U565 ( .A1(n686), .A2(n524), .ZN(n696) );
  NOR2_X1 U566 ( .A1(n721), .A2(n713), .ZN(n715) );
  NOR2_X1 U567 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U568 ( .A1(G2084), .A2(n731), .ZN(n712) );
  AND2_X1 U569 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U570 ( .A1(n526), .A2(n523), .ZN(n751) );
  NAND2_X1 U571 ( .A1(G160), .A2(G40), .ZN(n681) );
  AND2_X1 U572 ( .A1(n762), .A2(n525), .ZN(n763) );
  AND2_X1 U573 ( .A1(n532), .A2(G2104), .ZN(n869) );
  NOR2_X1 U574 ( .A1(G2104), .A2(n532), .ZN(n866) );
  NOR2_X1 U575 ( .A1(G651), .A2(n631), .ZN(n643) );
  NOR2_X1 U576 ( .A1(n536), .A2(n535), .ZN(G160) );
  AND2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n865) );
  NAND2_X1 U578 ( .A1(n865), .A2(G113), .ZN(n530) );
  INV_X1 U579 ( .A(G2105), .ZN(n532) );
  NAND2_X1 U580 ( .A1(G101), .A2(n869), .ZN(n528) );
  XOR2_X1 U581 ( .A(KEYINPUT23), .B(n528), .Z(n529) );
  NAND2_X1 U582 ( .A1(n530), .A2(n529), .ZN(n536) );
  NOR2_X1 U583 ( .A1(G2105), .A2(G2104), .ZN(n531) );
  NAND2_X1 U584 ( .A1(G137), .A2(n870), .ZN(n534) );
  NAND2_X1 U585 ( .A1(G125), .A2(n866), .ZN(n533) );
  NAND2_X1 U586 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U587 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U588 ( .A(G57), .ZN(G237) );
  INV_X1 U589 ( .A(G132), .ZN(G219) );
  INV_X1 U590 ( .A(G82), .ZN(G220) );
  NOR2_X1 U591 ( .A1(G651), .A2(G543), .ZN(n638) );
  NAND2_X1 U592 ( .A1(G88), .A2(n638), .ZN(n538) );
  XOR2_X1 U593 ( .A(KEYINPUT0), .B(G543), .Z(n631) );
  INV_X1 U594 ( .A(G651), .ZN(n539) );
  NOR2_X1 U595 ( .A1(n631), .A2(n539), .ZN(n639) );
  NAND2_X1 U596 ( .A1(G75), .A2(n639), .ZN(n537) );
  NAND2_X1 U597 ( .A1(n538), .A2(n537), .ZN(n544) );
  NOR2_X1 U598 ( .A1(G543), .A2(n539), .ZN(n540) );
  XOR2_X1 U599 ( .A(KEYINPUT1), .B(n540), .Z(n642) );
  NAND2_X1 U600 ( .A1(G62), .A2(n642), .ZN(n542) );
  NAND2_X1 U601 ( .A1(G50), .A2(n643), .ZN(n541) );
  NAND2_X1 U602 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U603 ( .A1(n544), .A2(n543), .ZN(G166) );
  NAND2_X1 U604 ( .A1(G90), .A2(n638), .ZN(n546) );
  NAND2_X1 U605 ( .A1(G77), .A2(n639), .ZN(n545) );
  NAND2_X1 U606 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U607 ( .A(n547), .B(KEYINPUT9), .ZN(n549) );
  NAND2_X1 U608 ( .A1(G52), .A2(n643), .ZN(n548) );
  NAND2_X1 U609 ( .A1(n549), .A2(n548), .ZN(n552) );
  NAND2_X1 U610 ( .A1(G64), .A2(n642), .ZN(n550) );
  XNOR2_X1 U611 ( .A(KEYINPUT65), .B(n550), .ZN(n551) );
  NOR2_X1 U612 ( .A1(n552), .A2(n551), .ZN(G171) );
  NAND2_X1 U613 ( .A1(G63), .A2(n642), .ZN(n554) );
  NAND2_X1 U614 ( .A1(G51), .A2(n643), .ZN(n553) );
  NAND2_X1 U615 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U616 ( .A(n555), .B(KEYINPUT71), .ZN(n556) );
  XNOR2_X1 U617 ( .A(n556), .B(KEYINPUT6), .ZN(n563) );
  XNOR2_X1 U618 ( .A(KEYINPUT5), .B(KEYINPUT70), .ZN(n561) );
  NAND2_X1 U619 ( .A1(n638), .A2(G89), .ZN(n557) );
  XNOR2_X1 U620 ( .A(n557), .B(KEYINPUT4), .ZN(n559) );
  NAND2_X1 U621 ( .A1(G76), .A2(n639), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U623 ( .A(n561), .B(n560), .ZN(n562) );
  NAND2_X1 U624 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U625 ( .A(KEYINPUT7), .B(n564), .ZN(G168) );
  XOR2_X1 U626 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U627 ( .A1(G7), .A2(G661), .ZN(n565) );
  XNOR2_X1 U628 ( .A(n565), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U629 ( .A(G223), .ZN(n818) );
  NAND2_X1 U630 ( .A1(n818), .A2(G567), .ZN(n566) );
  XOR2_X1 U631 ( .A(KEYINPUT11), .B(n566), .Z(G234) );
  NAND2_X1 U632 ( .A1(G56), .A2(n642), .ZN(n567) );
  XOR2_X1 U633 ( .A(KEYINPUT14), .B(n567), .Z(n573) );
  NAND2_X1 U634 ( .A1(n638), .A2(G81), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n568), .B(KEYINPUT12), .ZN(n570) );
  NAND2_X1 U636 ( .A1(G68), .A2(n639), .ZN(n569) );
  NAND2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U638 ( .A(KEYINPUT13), .B(n571), .Z(n572) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U640 ( .A1(n643), .A2(G43), .ZN(n574) );
  NAND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n982) );
  INV_X1 U642 ( .A(G860), .ZN(n597) );
  OR2_X1 U643 ( .A1(n982), .A2(n597), .ZN(G153) );
  INV_X1 U644 ( .A(G868), .ZN(n657) );
  NOR2_X1 U645 ( .A1(n657), .A2(G171), .ZN(n576) );
  XNOR2_X1 U646 ( .A(n576), .B(KEYINPUT67), .ZN(n587) );
  NAND2_X1 U647 ( .A1(G79), .A2(n639), .ZN(n577) );
  XNOR2_X1 U648 ( .A(n577), .B(KEYINPUT68), .ZN(n584) );
  NAND2_X1 U649 ( .A1(G92), .A2(n638), .ZN(n579) );
  NAND2_X1 U650 ( .A1(G66), .A2(n642), .ZN(n578) );
  NAND2_X1 U651 ( .A1(n579), .A2(n578), .ZN(n582) );
  NAND2_X1 U652 ( .A1(G54), .A2(n643), .ZN(n580) );
  XNOR2_X1 U653 ( .A(KEYINPUT69), .B(n580), .ZN(n581) );
  NOR2_X1 U654 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U655 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U656 ( .A(KEYINPUT15), .B(n585), .ZN(n981) );
  OR2_X1 U657 ( .A1(G868), .A2(n981), .ZN(n586) );
  NAND2_X1 U658 ( .A1(n587), .A2(n586), .ZN(G284) );
  NAND2_X1 U659 ( .A1(G91), .A2(n638), .ZN(n589) );
  NAND2_X1 U660 ( .A1(G78), .A2(n639), .ZN(n588) );
  NAND2_X1 U661 ( .A1(n589), .A2(n588), .ZN(n592) );
  NAND2_X1 U662 ( .A1(n642), .A2(G65), .ZN(n590) );
  XOR2_X1 U663 ( .A(KEYINPUT66), .B(n590), .Z(n591) );
  NOR2_X1 U664 ( .A1(n592), .A2(n591), .ZN(n594) );
  NAND2_X1 U665 ( .A1(n643), .A2(G53), .ZN(n593) );
  NAND2_X1 U666 ( .A1(n594), .A2(n593), .ZN(G299) );
  NOR2_X1 U667 ( .A1(G286), .A2(n657), .ZN(n596) );
  NOR2_X1 U668 ( .A1(G868), .A2(G299), .ZN(n595) );
  NOR2_X1 U669 ( .A1(n596), .A2(n595), .ZN(G297) );
  NAND2_X1 U670 ( .A1(n597), .A2(G559), .ZN(n598) );
  NAND2_X1 U671 ( .A1(n598), .A2(n981), .ZN(n599) );
  XNOR2_X1 U672 ( .A(n599), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U673 ( .A1(G868), .A2(n982), .ZN(n602) );
  NAND2_X1 U674 ( .A1(G868), .A2(n981), .ZN(n600) );
  NOR2_X1 U675 ( .A1(G559), .A2(n600), .ZN(n601) );
  NOR2_X1 U676 ( .A1(n602), .A2(n601), .ZN(G282) );
  NAND2_X1 U677 ( .A1(n865), .A2(G111), .ZN(n603) );
  XNOR2_X1 U678 ( .A(n603), .B(KEYINPUT72), .ZN(n605) );
  NAND2_X1 U679 ( .A1(G99), .A2(n869), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U681 ( .A(n606), .B(KEYINPUT73), .ZN(n608) );
  NAND2_X1 U682 ( .A1(G135), .A2(n870), .ZN(n607) );
  NAND2_X1 U683 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n866), .A2(G123), .ZN(n609) );
  XOR2_X1 U685 ( .A(KEYINPUT18), .B(n609), .Z(n610) );
  NOR2_X1 U686 ( .A1(n611), .A2(n610), .ZN(n947) );
  XNOR2_X1 U687 ( .A(G2096), .B(n947), .ZN(n613) );
  INV_X1 U688 ( .A(G2100), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n613), .A2(n612), .ZN(G156) );
  NAND2_X1 U690 ( .A1(G86), .A2(n638), .ZN(n615) );
  NAND2_X1 U691 ( .A1(G61), .A2(n642), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U693 ( .A1(n639), .A2(G73), .ZN(n616) );
  XOR2_X1 U694 ( .A(KEYINPUT2), .B(n616), .Z(n617) );
  NOR2_X1 U695 ( .A1(n618), .A2(n617), .ZN(n619) );
  XOR2_X1 U696 ( .A(KEYINPUT77), .B(n619), .Z(n621) );
  NAND2_X1 U697 ( .A1(n643), .A2(G48), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U699 ( .A(KEYINPUT78), .B(n622), .ZN(G305) );
  NAND2_X1 U700 ( .A1(G72), .A2(n639), .ZN(n624) );
  NAND2_X1 U701 ( .A1(G60), .A2(n642), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n638), .A2(G85), .ZN(n625) );
  XOR2_X1 U704 ( .A(KEYINPUT64), .B(n625), .Z(n626) );
  NOR2_X1 U705 ( .A1(n627), .A2(n626), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n643), .A2(G47), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n629), .A2(n628), .ZN(G290) );
  NAND2_X1 U708 ( .A1(G74), .A2(G651), .ZN(n630) );
  XNOR2_X1 U709 ( .A(n630), .B(KEYINPUT76), .ZN(n636) );
  NAND2_X1 U710 ( .A1(G49), .A2(n643), .ZN(n633) );
  NAND2_X1 U711 ( .A1(G87), .A2(n631), .ZN(n632) );
  NAND2_X1 U712 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U713 ( .A1(n642), .A2(n634), .ZN(n635) );
  NAND2_X1 U714 ( .A1(n636), .A2(n635), .ZN(G288) );
  NAND2_X1 U715 ( .A1(G559), .A2(n981), .ZN(n637) );
  XNOR2_X1 U716 ( .A(n637), .B(n982), .ZN(n826) );
  NAND2_X1 U717 ( .A1(G93), .A2(n638), .ZN(n641) );
  NAND2_X1 U718 ( .A1(G80), .A2(n639), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n641), .A2(n640), .ZN(n648) );
  NAND2_X1 U720 ( .A1(G67), .A2(n642), .ZN(n645) );
  NAND2_X1 U721 ( .A1(G55), .A2(n643), .ZN(n644) );
  NAND2_X1 U722 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U723 ( .A(KEYINPUT74), .B(n646), .ZN(n647) );
  NOR2_X1 U724 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U725 ( .A(n649), .B(KEYINPUT75), .ZN(n828) );
  XNOR2_X1 U726 ( .A(G305), .B(n828), .ZN(n655) );
  XNOR2_X1 U727 ( .A(KEYINPUT19), .B(KEYINPUT79), .ZN(n651) );
  XNOR2_X1 U728 ( .A(G299), .B(G166), .ZN(n650) );
  XNOR2_X1 U729 ( .A(n651), .B(n650), .ZN(n652) );
  XOR2_X1 U730 ( .A(n652), .B(G288), .Z(n653) );
  XNOR2_X1 U731 ( .A(G290), .B(n653), .ZN(n654) );
  XNOR2_X1 U732 ( .A(n655), .B(n654), .ZN(n892) );
  XNOR2_X1 U733 ( .A(n826), .B(n892), .ZN(n656) );
  NAND2_X1 U734 ( .A1(n656), .A2(G868), .ZN(n659) );
  NAND2_X1 U735 ( .A1(n657), .A2(n828), .ZN(n658) );
  NAND2_X1 U736 ( .A1(n659), .A2(n658), .ZN(G295) );
  NAND2_X1 U737 ( .A1(G2084), .A2(G2078), .ZN(n660) );
  XOR2_X1 U738 ( .A(KEYINPUT20), .B(n660), .Z(n661) );
  NAND2_X1 U739 ( .A1(G2090), .A2(n661), .ZN(n662) );
  XNOR2_X1 U740 ( .A(KEYINPUT21), .B(n662), .ZN(n663) );
  NAND2_X1 U741 ( .A1(n663), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U742 ( .A(KEYINPUT80), .B(G44), .ZN(n664) );
  XNOR2_X1 U743 ( .A(n664), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U744 ( .A1(G220), .A2(G219), .ZN(n665) );
  XNOR2_X1 U745 ( .A(KEYINPUT22), .B(n665), .ZN(n666) );
  NAND2_X1 U746 ( .A1(n666), .A2(G96), .ZN(n667) );
  NOR2_X1 U747 ( .A1(n667), .A2(G218), .ZN(n668) );
  XNOR2_X1 U748 ( .A(n668), .B(KEYINPUT81), .ZN(n824) );
  NAND2_X1 U749 ( .A1(n824), .A2(G2106), .ZN(n672) );
  NAND2_X1 U750 ( .A1(G69), .A2(G120), .ZN(n669) );
  NOR2_X1 U751 ( .A1(G237), .A2(n669), .ZN(n670) );
  NAND2_X1 U752 ( .A1(G108), .A2(n670), .ZN(n825) );
  NAND2_X1 U753 ( .A1(n825), .A2(G567), .ZN(n671) );
  NAND2_X1 U754 ( .A1(n672), .A2(n671), .ZN(n829) );
  NAND2_X1 U755 ( .A1(G483), .A2(G661), .ZN(n673) );
  NOR2_X1 U756 ( .A1(n829), .A2(n673), .ZN(n823) );
  NAND2_X1 U757 ( .A1(n823), .A2(G36), .ZN(G176) );
  NAND2_X1 U758 ( .A1(G126), .A2(n866), .ZN(n675) );
  NAND2_X1 U759 ( .A1(G114), .A2(n865), .ZN(n674) );
  NAND2_X1 U760 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U761 ( .A(n676), .B(KEYINPUT82), .ZN(n680) );
  NAND2_X1 U762 ( .A1(G102), .A2(n869), .ZN(n678) );
  NAND2_X1 U763 ( .A1(G138), .A2(n870), .ZN(n677) );
  NAND2_X1 U764 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U765 ( .A1(n680), .A2(n679), .ZN(G164) );
  INV_X1 U766 ( .A(G166), .ZN(G303) );
  INV_X1 U767 ( .A(G171), .ZN(G301) );
  XNOR2_X1 U768 ( .A(G305), .B(G1981), .ZN(n968) );
  NOR2_X1 U769 ( .A1(G164), .A2(G1384), .ZN(n782) );
  NAND2_X1 U770 ( .A1(G8), .A2(n731), .ZN(n761) );
  NOR2_X1 U771 ( .A1(G1966), .A2(n761), .ZN(n721) );
  INV_X1 U772 ( .A(G1996), .ZN(n848) );
  NOR2_X1 U773 ( .A1(n731), .A2(n848), .ZN(n683) );
  INV_X1 U774 ( .A(KEYINPUT26), .ZN(n682) );
  XNOR2_X1 U775 ( .A(n683), .B(n682), .ZN(n686) );
  NAND2_X1 U776 ( .A1(n731), .A2(G1341), .ZN(n685) );
  NOR2_X1 U777 ( .A1(n981), .A2(n696), .ZN(n690) );
  NAND2_X1 U778 ( .A1(n705), .A2(G2067), .ZN(n688) );
  NAND2_X1 U779 ( .A1(G1348), .A2(n731), .ZN(n687) );
  NAND2_X1 U780 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U781 ( .A1(n690), .A2(n689), .ZN(n695) );
  NAND2_X1 U782 ( .A1(n705), .A2(G2072), .ZN(n691) );
  XOR2_X1 U783 ( .A(KEYINPUT27), .B(n691), .Z(n693) );
  NAND2_X1 U784 ( .A1(G1956), .A2(n731), .ZN(n692) );
  NAND2_X1 U785 ( .A1(n693), .A2(n692), .ZN(n700) );
  NOR2_X1 U786 ( .A1(G299), .A2(n700), .ZN(n694) );
  NOR2_X1 U787 ( .A1(n695), .A2(n694), .ZN(n698) );
  NAND2_X1 U788 ( .A1(n981), .A2(n696), .ZN(n697) );
  NAND2_X1 U789 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U790 ( .A(n699), .B(KEYINPUT91), .ZN(n703) );
  NAND2_X1 U791 ( .A1(G299), .A2(n700), .ZN(n701) );
  XOR2_X1 U792 ( .A(KEYINPUT28), .B(n701), .Z(n702) );
  NOR2_X1 U793 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U794 ( .A(n704), .B(KEYINPUT29), .ZN(n709) );
  NAND2_X1 U795 ( .A1(G1961), .A2(n731), .ZN(n707) );
  XOR2_X1 U796 ( .A(G2078), .B(KEYINPUT25), .Z(n919) );
  NAND2_X1 U797 ( .A1(n705), .A2(n919), .ZN(n706) );
  NAND2_X1 U798 ( .A1(n707), .A2(n706), .ZN(n710) );
  OR2_X1 U799 ( .A1(n710), .A2(G301), .ZN(n708) );
  NAND2_X1 U800 ( .A1(n709), .A2(n708), .ZN(n727) );
  NAND2_X1 U801 ( .A1(G301), .A2(n710), .ZN(n711) );
  XNOR2_X1 U802 ( .A(n711), .B(KEYINPUT93), .ZN(n718) );
  XOR2_X1 U803 ( .A(KEYINPUT90), .B(n712), .Z(n723) );
  NAND2_X1 U804 ( .A1(G8), .A2(n723), .ZN(n713) );
  XOR2_X1 U805 ( .A(KEYINPUT92), .B(KEYINPUT30), .Z(n714) );
  XNOR2_X1 U806 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U807 ( .A1(n716), .A2(G168), .ZN(n717) );
  XOR2_X1 U808 ( .A(KEYINPUT31), .B(n719), .Z(n728) );
  AND2_X1 U809 ( .A1(n727), .A2(n728), .ZN(n720) );
  NOR2_X1 U810 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U811 ( .A(n722), .B(KEYINPUT94), .ZN(n726) );
  INV_X1 U812 ( .A(n723), .ZN(n724) );
  NAND2_X1 U813 ( .A1(G8), .A2(n724), .ZN(n725) );
  NAND2_X1 U814 ( .A1(n726), .A2(n725), .ZN(n741) );
  NAND2_X1 U815 ( .A1(n728), .A2(n727), .ZN(n730) );
  AND2_X1 U816 ( .A1(G286), .A2(G8), .ZN(n729) );
  NAND2_X1 U817 ( .A1(n730), .A2(n729), .ZN(n738) );
  INV_X1 U818 ( .A(G8), .ZN(n736) );
  NOR2_X1 U819 ( .A1(G1971), .A2(n761), .ZN(n733) );
  NOR2_X1 U820 ( .A1(G2090), .A2(n731), .ZN(n732) );
  NOR2_X1 U821 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U822 ( .A1(n734), .A2(G303), .ZN(n735) );
  OR2_X1 U823 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U824 ( .A(n739), .B(KEYINPUT32), .ZN(n740) );
  NAND2_X1 U825 ( .A1(n741), .A2(n740), .ZN(n754) );
  NOR2_X1 U826 ( .A1(G1971), .A2(G303), .ZN(n742) );
  NOR2_X1 U827 ( .A1(G1976), .A2(G288), .ZN(n976) );
  NOR2_X1 U828 ( .A1(n742), .A2(n976), .ZN(n743) );
  INV_X1 U829 ( .A(KEYINPUT33), .ZN(n750) );
  AND2_X1 U830 ( .A1(n743), .A2(n750), .ZN(n744) );
  AND2_X1 U831 ( .A1(n754), .A2(n744), .ZN(n752) );
  NAND2_X1 U832 ( .A1(KEYINPUT33), .A2(n976), .ZN(n745) );
  XOR2_X1 U833 ( .A(KEYINPUT95), .B(n745), .Z(n746) );
  NOR2_X1 U834 ( .A1(n761), .A2(n746), .ZN(n747) );
  NAND2_X1 U835 ( .A1(G1976), .A2(G288), .ZN(n973) );
  INV_X1 U836 ( .A(n761), .ZN(n748) );
  NAND2_X1 U837 ( .A1(n973), .A2(n748), .ZN(n749) );
  XNOR2_X1 U838 ( .A(n527), .B(KEYINPUT97), .ZN(n753) );
  NOR2_X1 U839 ( .A1(G2090), .A2(G303), .ZN(n755) );
  NAND2_X1 U840 ( .A1(G8), .A2(n755), .ZN(n756) );
  NAND2_X1 U841 ( .A1(n754), .A2(n756), .ZN(n757) );
  NAND2_X1 U842 ( .A1(n757), .A2(n761), .ZN(n762) );
  NOR2_X1 U843 ( .A1(G305), .A2(G1981), .ZN(n758) );
  XNOR2_X1 U844 ( .A(n758), .B(KEYINPUT89), .ZN(n759) );
  XNOR2_X1 U845 ( .A(KEYINPUT24), .B(n759), .ZN(n760) );
  NAND2_X1 U846 ( .A1(n522), .A2(n763), .ZN(n800) );
  NAND2_X1 U847 ( .A1(G95), .A2(n869), .ZN(n765) );
  NAND2_X1 U848 ( .A1(G131), .A2(n870), .ZN(n764) );
  NAND2_X1 U849 ( .A1(n765), .A2(n764), .ZN(n769) );
  NAND2_X1 U850 ( .A1(G107), .A2(n865), .ZN(n767) );
  NAND2_X1 U851 ( .A1(G119), .A2(n866), .ZN(n766) );
  NAND2_X1 U852 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U853 ( .A1(n769), .A2(n768), .ZN(n885) );
  INV_X1 U854 ( .A(G1991), .ZN(n916) );
  NOR2_X1 U855 ( .A1(n885), .A2(n916), .ZN(n779) );
  NAND2_X1 U856 ( .A1(n866), .A2(G129), .ZN(n776) );
  NAND2_X1 U857 ( .A1(G117), .A2(n865), .ZN(n771) );
  NAND2_X1 U858 ( .A1(G141), .A2(n870), .ZN(n770) );
  NAND2_X1 U859 ( .A1(n771), .A2(n770), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n869), .A2(G105), .ZN(n772) );
  XOR2_X1 U861 ( .A(KEYINPUT38), .B(n772), .Z(n773) );
  NOR2_X1 U862 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U863 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U864 ( .A(KEYINPUT87), .B(n777), .ZN(n886) );
  NOR2_X1 U865 ( .A1(n886), .A2(n848), .ZN(n778) );
  NOR2_X1 U866 ( .A1(n779), .A2(n778), .ZN(n952) );
  INV_X1 U867 ( .A(n780), .ZN(n781) );
  NOR2_X1 U868 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U869 ( .A(KEYINPUT84), .B(n783), .ZN(n812) );
  XOR2_X1 U870 ( .A(KEYINPUT88), .B(n812), .Z(n784) );
  NOR2_X1 U871 ( .A1(n952), .A2(n784), .ZN(n803) );
  INV_X1 U872 ( .A(n803), .ZN(n796) );
  NAND2_X1 U873 ( .A1(G104), .A2(n869), .ZN(n786) );
  NAND2_X1 U874 ( .A1(G140), .A2(n870), .ZN(n785) );
  NAND2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U876 ( .A(KEYINPUT34), .B(n787), .ZN(n793) );
  NAND2_X1 U877 ( .A1(n865), .A2(G116), .ZN(n788) );
  XOR2_X1 U878 ( .A(KEYINPUT85), .B(n788), .Z(n790) );
  NAND2_X1 U879 ( .A1(n866), .A2(G128), .ZN(n789) );
  NAND2_X1 U880 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U881 ( .A(n791), .B(KEYINPUT35), .Z(n792) );
  NOR2_X1 U882 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U883 ( .A(KEYINPUT36), .B(n794), .Z(n795) );
  XOR2_X1 U884 ( .A(KEYINPUT86), .B(n795), .Z(n889) );
  XNOR2_X1 U885 ( .A(G2067), .B(KEYINPUT37), .ZN(n810) );
  NOR2_X1 U886 ( .A1(n889), .A2(n810), .ZN(n955) );
  NAND2_X1 U887 ( .A1(n955), .A2(n812), .ZN(n808) );
  NAND2_X1 U888 ( .A1(n796), .A2(n808), .ZN(n798) );
  XNOR2_X1 U889 ( .A(G1986), .B(G290), .ZN(n972) );
  AND2_X1 U890 ( .A1(n972), .A2(n812), .ZN(n797) );
  NOR2_X1 U891 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U892 ( .A1(n800), .A2(n799), .ZN(n815) );
  AND2_X1 U893 ( .A1(n848), .A2(n886), .ZN(n943) );
  NOR2_X1 U894 ( .A1(G1986), .A2(G290), .ZN(n801) );
  AND2_X1 U895 ( .A1(n916), .A2(n885), .ZN(n948) );
  NOR2_X1 U896 ( .A1(n801), .A2(n948), .ZN(n802) );
  NOR2_X1 U897 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U898 ( .A(n804), .B(KEYINPUT98), .ZN(n805) );
  NOR2_X1 U899 ( .A1(n943), .A2(n805), .ZN(n807) );
  XOR2_X1 U900 ( .A(KEYINPUT39), .B(KEYINPUT99), .Z(n806) );
  XNOR2_X1 U901 ( .A(n807), .B(n806), .ZN(n809) );
  NAND2_X1 U902 ( .A1(n809), .A2(n808), .ZN(n811) );
  NAND2_X1 U903 ( .A1(n889), .A2(n810), .ZN(n958) );
  NAND2_X1 U904 ( .A1(n811), .A2(n958), .ZN(n813) );
  NAND2_X1 U905 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U906 ( .A1(n815), .A2(n814), .ZN(n817) );
  XNOR2_X1 U907 ( .A(KEYINPUT100), .B(KEYINPUT40), .ZN(n816) );
  XNOR2_X1 U908 ( .A(n817), .B(n816), .ZN(G329) );
  NAND2_X1 U909 ( .A1(n818), .A2(G2106), .ZN(n819) );
  XNOR2_X1 U910 ( .A(n819), .B(KEYINPUT102), .ZN(G217) );
  AND2_X1 U911 ( .A1(G15), .A2(G2), .ZN(n820) );
  NAND2_X1 U912 ( .A1(G661), .A2(n820), .ZN(G259) );
  NAND2_X1 U913 ( .A1(G3), .A2(G1), .ZN(n821) );
  XOR2_X1 U914 ( .A(KEYINPUT103), .B(n821), .Z(n822) );
  NAND2_X1 U915 ( .A1(n823), .A2(n822), .ZN(G188) );
  INV_X1 U917 ( .A(G120), .ZN(G236) );
  INV_X1 U918 ( .A(G96), .ZN(G221) );
  INV_X1 U919 ( .A(G69), .ZN(G235) );
  NOR2_X1 U920 ( .A1(n825), .A2(n824), .ZN(G325) );
  INV_X1 U921 ( .A(G325), .ZN(G261) );
  NOR2_X1 U922 ( .A1(G860), .A2(n826), .ZN(n827) );
  XOR2_X1 U923 ( .A(n828), .B(n827), .Z(G145) );
  INV_X1 U924 ( .A(n829), .ZN(G319) );
  XOR2_X1 U925 ( .A(G2096), .B(KEYINPUT43), .Z(n831) );
  XNOR2_X1 U926 ( .A(G2090), .B(G2678), .ZN(n830) );
  XNOR2_X1 U927 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U928 ( .A(n832), .B(KEYINPUT104), .Z(n834) );
  XNOR2_X1 U929 ( .A(G2067), .B(G2072), .ZN(n833) );
  XNOR2_X1 U930 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U931 ( .A(KEYINPUT42), .B(G2100), .Z(n836) );
  XNOR2_X1 U932 ( .A(G2084), .B(G2078), .ZN(n835) );
  XNOR2_X1 U933 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U934 ( .A(n838), .B(n837), .ZN(G227) );
  XOR2_X1 U935 ( .A(G1991), .B(G1981), .Z(n840) );
  XNOR2_X1 U936 ( .A(G1966), .B(G1961), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U938 ( .A(G1986), .B(G1976), .Z(n842) );
  XNOR2_X1 U939 ( .A(G1956), .B(G1971), .ZN(n841) );
  XNOR2_X1 U940 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U941 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U942 ( .A(G2474), .B(KEYINPUT41), .ZN(n845) );
  XNOR2_X1 U943 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U944 ( .A(KEYINPUT105), .B(n847), .ZN(n849) );
  XNOR2_X1 U945 ( .A(n849), .B(n848), .ZN(G229) );
  NAND2_X1 U946 ( .A1(G124), .A2(n866), .ZN(n850) );
  XNOR2_X1 U947 ( .A(n850), .B(KEYINPUT44), .ZN(n852) );
  NAND2_X1 U948 ( .A1(n865), .A2(G112), .ZN(n851) );
  NAND2_X1 U949 ( .A1(n852), .A2(n851), .ZN(n856) );
  NAND2_X1 U950 ( .A1(G100), .A2(n869), .ZN(n854) );
  NAND2_X1 U951 ( .A1(G136), .A2(n870), .ZN(n853) );
  NAND2_X1 U952 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U953 ( .A1(n856), .A2(n855), .ZN(G162) );
  XNOR2_X1 U954 ( .A(G164), .B(n947), .ZN(n864) );
  NAND2_X1 U955 ( .A1(G103), .A2(n869), .ZN(n858) );
  NAND2_X1 U956 ( .A1(G139), .A2(n870), .ZN(n857) );
  NAND2_X1 U957 ( .A1(n858), .A2(n857), .ZN(n863) );
  NAND2_X1 U958 ( .A1(G115), .A2(n865), .ZN(n860) );
  NAND2_X1 U959 ( .A1(G127), .A2(n866), .ZN(n859) );
  NAND2_X1 U960 ( .A1(n860), .A2(n859), .ZN(n861) );
  XOR2_X1 U961 ( .A(KEYINPUT47), .B(n861), .Z(n862) );
  NOR2_X1 U962 ( .A1(n863), .A2(n862), .ZN(n938) );
  XNOR2_X1 U963 ( .A(n864), .B(n938), .ZN(n878) );
  NAND2_X1 U964 ( .A1(G118), .A2(n865), .ZN(n868) );
  NAND2_X1 U965 ( .A1(G130), .A2(n866), .ZN(n867) );
  NAND2_X1 U966 ( .A1(n868), .A2(n867), .ZN(n876) );
  NAND2_X1 U967 ( .A1(G106), .A2(n869), .ZN(n872) );
  NAND2_X1 U968 ( .A1(G142), .A2(n870), .ZN(n871) );
  NAND2_X1 U969 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U970 ( .A(KEYINPUT45), .B(n873), .Z(n874) );
  XNOR2_X1 U971 ( .A(KEYINPUT106), .B(n874), .ZN(n875) );
  NOR2_X1 U972 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U973 ( .A(n878), .B(n877), .Z(n880) );
  XNOR2_X1 U974 ( .A(G160), .B(G162), .ZN(n879) );
  XNOR2_X1 U975 ( .A(n880), .B(n879), .ZN(n884) );
  XOR2_X1 U976 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n882) );
  XNOR2_X1 U977 ( .A(KEYINPUT108), .B(KEYINPUT107), .ZN(n881) );
  XNOR2_X1 U978 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U979 ( .A(n884), .B(n883), .Z(n888) );
  XNOR2_X1 U980 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U981 ( .A(n888), .B(n887), .ZN(n890) );
  XNOR2_X1 U982 ( .A(n890), .B(n889), .ZN(n891) );
  NOR2_X1 U983 ( .A1(G37), .A2(n891), .ZN(G395) );
  XNOR2_X1 U984 ( .A(n982), .B(n892), .ZN(n894) );
  XNOR2_X1 U985 ( .A(G171), .B(n981), .ZN(n893) );
  XNOR2_X1 U986 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U987 ( .A(G286), .B(n895), .Z(n896) );
  NOR2_X1 U988 ( .A1(G37), .A2(n896), .ZN(G397) );
  XOR2_X1 U989 ( .A(KEYINPUT101), .B(G2451), .Z(n898) );
  XNOR2_X1 U990 ( .A(G2446), .B(G2427), .ZN(n897) );
  XNOR2_X1 U991 ( .A(n898), .B(n897), .ZN(n905) );
  XOR2_X1 U992 ( .A(G2438), .B(G2435), .Z(n900) );
  XNOR2_X1 U993 ( .A(G2443), .B(G2430), .ZN(n899) );
  XNOR2_X1 U994 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U995 ( .A(n901), .B(G2454), .Z(n903) );
  XNOR2_X1 U996 ( .A(G1348), .B(G1341), .ZN(n902) );
  XNOR2_X1 U997 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U998 ( .A(n905), .B(n904), .ZN(n906) );
  NAND2_X1 U999 ( .A1(n906), .A2(G14), .ZN(n912) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n912), .ZN(n909) );
  NOR2_X1 U1001 ( .A1(G227), .A2(G229), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(KEYINPUT49), .B(n907), .ZN(n908) );
  NOR2_X1 U1003 ( .A1(n909), .A2(n908), .ZN(n911) );
  NOR2_X1 U1004 ( .A1(G395), .A2(G397), .ZN(n910) );
  NAND2_X1 U1005 ( .A1(n911), .A2(n910), .ZN(G225) );
  INV_X1 U1006 ( .A(G225), .ZN(G308) );
  INV_X1 U1007 ( .A(G108), .ZN(G238) );
  INV_X1 U1008 ( .A(n912), .ZN(G401) );
  XNOR2_X1 U1009 ( .A(KEYINPUT54), .B(KEYINPUT116), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(n913), .B(G34), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(G2084), .B(n914), .ZN(n934) );
  XNOR2_X1 U1012 ( .A(KEYINPUT114), .B(KEYINPUT53), .ZN(n928) );
  XNOR2_X1 U1013 ( .A(KEYINPUT113), .B(G1996), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(n915), .B(G32), .ZN(n923) );
  XOR2_X1 U1015 ( .A(G2067), .B(G26), .Z(n918) );
  XNOR2_X1 U1016 ( .A(n916), .B(G25), .ZN(n917) );
  NAND2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n921) );
  XNOR2_X1 U1018 ( .A(G27), .B(n919), .ZN(n920) );
  NOR2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1020 ( .A1(n923), .A2(n922), .ZN(n926) );
  XOR2_X1 U1021 ( .A(G2072), .B(G33), .Z(n924) );
  NAND2_X1 U1022 ( .A1(G28), .A2(n924), .ZN(n925) );
  NOR2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1024 ( .A(n928), .B(n927), .ZN(n931) );
  XNOR2_X1 U1025 ( .A(G2090), .B(G35), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(KEYINPUT112), .B(n929), .ZN(n930) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1028 ( .A(KEYINPUT115), .B(n932), .ZN(n933) );
  NOR2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1030 ( .A(n935), .B(KEYINPUT55), .ZN(n937) );
  XNOR2_X1 U1031 ( .A(G29), .B(KEYINPUT117), .ZN(n936) );
  NAND2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n1025) );
  XOR2_X1 U1033 ( .A(G2072), .B(n938), .Z(n940) );
  XOR2_X1 U1034 ( .A(G164), .B(G2078), .Z(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1036 ( .A(KEYINPUT50), .B(n941), .ZN(n946) );
  XOR2_X1 U1037 ( .A(G2090), .B(G162), .Z(n942) );
  NOR2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1039 ( .A(KEYINPUT51), .B(n944), .Z(n945) );
  NAND2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n960) );
  XNOR2_X1 U1041 ( .A(G160), .B(G2084), .ZN(n950) );
  NOR2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1043 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(KEYINPUT109), .B(n951), .ZN(n953) );
  NAND2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1046 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1047 ( .A(n956), .B(KEYINPUT110), .ZN(n957) );
  NAND2_X1 U1048 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1049 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1050 ( .A(KEYINPUT52), .B(n961), .Z(n962) );
  NOR2_X1 U1051 ( .A1(KEYINPUT55), .A2(n962), .ZN(n963) );
  XNOR2_X1 U1052 ( .A(KEYINPUT111), .B(n963), .ZN(n964) );
  NAND2_X1 U1053 ( .A1(n964), .A2(G29), .ZN(n965) );
  NAND2_X1 U1054 ( .A1(n965), .A2(G11), .ZN(n1023) );
  XNOR2_X1 U1055 ( .A(G16), .B(KEYINPUT56), .ZN(n993) );
  XOR2_X1 U1056 ( .A(G1966), .B(G168), .Z(n966) );
  XNOR2_X1 U1057 ( .A(KEYINPUT118), .B(n966), .ZN(n967) );
  NOR2_X1 U1058 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1059 ( .A(KEYINPUT119), .B(n969), .ZN(n970) );
  XNOR2_X1 U1060 ( .A(n970), .B(KEYINPUT57), .ZN(n991) );
  XNOR2_X1 U1061 ( .A(G1956), .B(G299), .ZN(n971) );
  NOR2_X1 U1062 ( .A1(n972), .A2(n971), .ZN(n974) );
  NAND2_X1 U1063 ( .A1(n974), .A2(n973), .ZN(n988) );
  XNOR2_X1 U1064 ( .A(G1961), .B(KEYINPUT120), .ZN(n975) );
  XNOR2_X1 U1065 ( .A(n975), .B(G301), .ZN(n980) );
  XNOR2_X1 U1066 ( .A(n976), .B(KEYINPUT121), .ZN(n978) );
  XNOR2_X1 U1067 ( .A(G166), .B(G1971), .ZN(n977) );
  NAND2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1069 ( .A1(n980), .A2(n979), .ZN(n986) );
  XOR2_X1 U1070 ( .A(G1348), .B(n981), .Z(n984) );
  XNOR2_X1 U1071 ( .A(n982), .B(G1341), .ZN(n983) );
  NOR2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1073 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1074 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1075 ( .A(KEYINPUT122), .B(n989), .ZN(n990) );
  NAND2_X1 U1076 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1077 ( .A1(n993), .A2(n992), .ZN(n1020) );
  XNOR2_X1 U1078 ( .A(G1971), .B(G22), .ZN(n995) );
  XNOR2_X1 U1079 ( .A(G1976), .B(G23), .ZN(n994) );
  NOR2_X1 U1080 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1081 ( .A(KEYINPUT126), .B(n996), .Z(n998) );
  XNOR2_X1 U1082 ( .A(G1986), .B(G24), .ZN(n997) );
  NOR2_X1 U1083 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1084 ( .A(KEYINPUT58), .B(n999), .ZN(n1003) );
  XNOR2_X1 U1085 ( .A(G1966), .B(G21), .ZN(n1001) );
  XNOR2_X1 U1086 ( .A(G1961), .B(G5), .ZN(n1000) );
  NOR2_X1 U1087 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1088 ( .A1(n1003), .A2(n1002), .ZN(n1015) );
  XOR2_X1 U1089 ( .A(G1341), .B(G19), .Z(n1006) );
  XOR2_X1 U1090 ( .A(G20), .B(KEYINPUT124), .Z(n1004) );
  XNOR2_X1 U1091 ( .A(G1956), .B(n1004), .ZN(n1005) );
  NAND2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1009) );
  XOR2_X1 U1093 ( .A(KEYINPUT59), .B(G1348), .Z(n1007) );
  XNOR2_X1 U1094 ( .A(G4), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1012) );
  XNOR2_X1 U1096 ( .A(G1981), .B(KEYINPUT125), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(n1010), .B(G6), .ZN(n1011) );
  NAND2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(KEYINPUT60), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1101 ( .A(n1016), .B(KEYINPUT61), .ZN(n1018) );
  XNOR2_X1 U1102 ( .A(G16), .B(KEYINPUT123), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1105 ( .A(KEYINPUT127), .B(n1021), .Z(n1022) );
  NOR2_X1 U1106 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1107 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1026), .Z(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

