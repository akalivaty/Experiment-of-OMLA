

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805;

  INV_X1 U373 ( .A(n804), .ZN(n356) );
  XNOR2_X1 U374 ( .A(n635), .B(n634), .ZN(n804) );
  NAND2_X1 U375 ( .A1(n355), .A2(n354), .ZN(n353) );
  XNOR2_X1 U376 ( .A(n613), .B(KEYINPUT30), .ZN(n355) );
  INV_X1 U377 ( .A(n615), .ZN(n354) );
  OR2_X1 U378 ( .A1(n688), .A2(G902), .ZN(n481) );
  INV_X1 U379 ( .A(n622), .ZN(n504) );
  BUF_X1 U380 ( .A(n493), .Z(n494) );
  XNOR2_X1 U381 ( .A(n476), .B(n360), .ZN(n478) );
  XNOR2_X2 U382 ( .A(n352), .B(n641), .ZN(n426) );
  NAND2_X1 U383 ( .A1(n639), .A2(n640), .ZN(n352) );
  XNOR2_X2 U384 ( .A(KEYINPUT5), .B(G137), .ZN(n471) );
  INV_X1 U385 ( .A(n353), .ZN(n617) );
  NAND2_X1 U386 ( .A1(n357), .A2(n356), .ZN(n638) );
  INV_X1 U387 ( .A(n670), .ZN(n357) );
  NAND2_X1 U388 ( .A1(n358), .A2(n361), .ZN(n552) );
  NAND2_X1 U389 ( .A1(n370), .A2(n398), .ZN(n358) );
  NAND2_X1 U390 ( .A1(n437), .A2(n436), .ZN(n374) );
  XNOR2_X2 U391 ( .A(n468), .B(n438), .ZN(n437) );
  XNOR2_X2 U392 ( .A(n500), .B(KEYINPUT90), .ZN(n501) );
  NAND2_X2 U393 ( .A1(n602), .A2(n509), .ZN(n511) );
  XNOR2_X2 U394 ( .A(n365), .B(KEYINPUT19), .ZN(n602) );
  XNOR2_X2 U395 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X2 U396 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X2 U397 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X2 U398 ( .A(n460), .B(n459), .ZN(n693) );
  NAND2_X2 U399 ( .A1(n371), .A2(n504), .ZN(n365) );
  NOR2_X1 U400 ( .A1(G953), .A2(G237), .ZN(n531) );
  NAND2_X2 U401 ( .A1(n552), .A2(n734), .ZN(n468) );
  NAND2_X1 U402 ( .A1(n426), .A2(n651), .ZN(n720) );
  AND2_X1 U403 ( .A1(n408), .A2(n406), .ZN(n410) );
  AND2_X1 U404 ( .A1(n559), .A2(n647), .ZN(n587) );
  OR2_X1 U405 ( .A1(n644), .A2(n633), .ZN(n635) );
  XNOR2_X1 U406 ( .A(n626), .B(KEYINPUT41), .ZN(n750) );
  NOR2_X1 U407 ( .A1(n420), .A2(n418), .ZN(n598) );
  AND2_X1 U408 ( .A1(n368), .A2(n448), .ZN(n369) );
  INV_X1 U409 ( .A(G146), .ZN(n470) );
  XNOR2_X2 U410 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n483) );
  XNOR2_X1 U411 ( .A(G140), .B(G137), .ZN(n452) );
  BUF_X1 U412 ( .A(n477), .Z(n359) );
  BUF_X1 U413 ( .A(n491), .Z(n360) );
  XNOR2_X2 U414 ( .A(n491), .B(n490), .ZN(n794) );
  INV_X1 U415 ( .A(KEYINPUT47), .ZN(n413) );
  NAND2_X1 U416 ( .A1(n391), .A2(n390), .ZN(n389) );
  OR2_X1 U417 ( .A1(n693), .A2(n392), .ZN(n391) );
  OR2_X1 U418 ( .A1(n416), .A2(n413), .ZN(n407) );
  INV_X1 U419 ( .A(n665), .ZN(n411) );
  NAND2_X1 U420 ( .A1(n402), .A2(n525), .ZN(n401) );
  NAND2_X1 U421 ( .A1(n410), .A2(n409), .ZN(n415) );
  OR2_X1 U422 ( .A1(n771), .A2(n413), .ZN(n409) );
  NAND2_X1 U423 ( .A1(n654), .A2(n423), .ZN(n422) );
  INV_X1 U424 ( .A(KEYINPUT8), .ZN(n450) );
  XOR2_X1 U425 ( .A(G107), .B(KEYINPUT7), .Z(n515) );
  XNOR2_X1 U426 ( .A(KEYINPUT101), .B(KEYINPUT9), .ZN(n514) );
  XNOR2_X1 U427 ( .A(G113), .B(G119), .ZN(n428) );
  XNOR2_X1 U428 ( .A(G128), .B(G119), .ZN(n455) );
  XNOR2_X1 U429 ( .A(n454), .B(KEYINPUT23), .ZN(n405) );
  AND2_X1 U430 ( .A1(n518), .A2(G221), .ZN(n404) );
  XNOR2_X1 U431 ( .A(n551), .B(n550), .ZN(n559) );
  INV_X1 U432 ( .A(n389), .ZN(n381) );
  AND2_X1 U433 ( .A1(n407), .A2(n411), .ZN(n406) );
  NAND2_X1 U434 ( .A1(n385), .A2(n363), .ZN(n396) );
  NAND2_X1 U435 ( .A1(n402), .A2(n403), .ZN(n384) );
  NAND2_X1 U436 ( .A1(n395), .A2(KEYINPUT1), .ZN(n394) );
  INV_X1 U437 ( .A(n401), .ZN(n395) );
  XNOR2_X1 U438 ( .A(G104), .B(G140), .ZN(n533) );
  XNOR2_X1 U439 ( .A(G113), .B(G131), .ZN(n534) );
  XNOR2_X1 U440 ( .A(G143), .B(KEYINPUT12), .ZN(n529) );
  XNOR2_X1 U441 ( .A(G122), .B(KEYINPUT99), .ZN(n528) );
  XNOR2_X1 U442 ( .A(KEYINPUT87), .B(KEYINPUT89), .ZN(n486) );
  NAND2_X1 U443 ( .A1(G237), .A2(G234), .ZN(n505) );
  XNOR2_X1 U444 ( .A(n609), .B(KEYINPUT38), .ZN(n728) );
  NAND2_X1 U445 ( .A1(n738), .A2(n383), .ZN(n420) );
  NAND2_X1 U446 ( .A1(n419), .A2(n616), .ZN(n418) );
  NOR2_X2 U447 ( .A1(n389), .A2(n382), .ZN(n734) );
  NAND2_X1 U448 ( .A1(n387), .A2(n383), .ZN(n382) );
  XNOR2_X1 U449 ( .A(KEYINPUT70), .B(G101), .ZN(n474) );
  XNOR2_X1 U450 ( .A(G131), .B(G134), .ZN(n441) );
  NAND2_X1 U451 ( .A1(n654), .A2(KEYINPUT2), .ZN(n427) );
  INV_X1 U452 ( .A(KEYINPUT66), .ZN(n439) );
  XNOR2_X1 U453 ( .A(G122), .B(G134), .ZN(n513) );
  BUF_X1 U454 ( .A(n724), .Z(n760) );
  INV_X1 U455 ( .A(KEYINPUT94), .ZN(n512) );
  XNOR2_X1 U456 ( .A(n405), .B(n404), .ZN(n460) );
  NAND2_X1 U457 ( .A1(n661), .A2(n660), .ZN(n706) );
  AND2_X1 U458 ( .A1(n414), .A2(n553), .ZN(n783) );
  XNOR2_X1 U459 ( .A(n555), .B(n554), .ZN(n556) );
  INV_X1 U460 ( .A(KEYINPUT68), .ZN(n554) );
  XNOR2_X1 U461 ( .A(n374), .B(n364), .ZN(n724) );
  INV_X1 U462 ( .A(n737), .ZN(n383) );
  INV_X1 U463 ( .A(KEYINPUT1), .ZN(n399) );
  NAND2_X1 U464 ( .A1(n381), .A2(n387), .ZN(n738) );
  AND2_X1 U465 ( .A1(n396), .A2(n393), .ZN(n361) );
  AND2_X1 U466 ( .A1(n651), .A2(n654), .ZN(n362) );
  AND2_X1 U467 ( .A1(n384), .A2(KEYINPUT1), .ZN(n363) );
  AND2_X1 U468 ( .A1(n602), .A2(n627), .ZN(n771) );
  XOR2_X1 U469 ( .A(KEYINPUT86), .B(KEYINPUT33), .Z(n364) );
  INV_X1 U470 ( .A(KEYINPUT78), .ZN(n423) );
  XNOR2_X2 U471 ( .A(n372), .B(n501), .ZN(n371) );
  XNOR2_X2 U472 ( .A(n373), .B(n439), .ZN(n366) );
  XNOR2_X1 U473 ( .A(n373), .B(n439), .ZN(n701) );
  NAND2_X2 U474 ( .A1(n376), .A2(n378), .ZN(n373) );
  BUF_X1 U475 ( .A(n655), .Z(n657) );
  BUF_X1 U476 ( .A(n669), .Z(n367) );
  XNOR2_X1 U477 ( .A(n672), .B(n447), .ZN(n368) );
  XNOR2_X1 U478 ( .A(n672), .B(n447), .ZN(n711) );
  OR2_X2 U479 ( .A1(n711), .A2(n401), .ZN(n400) );
  NOR2_X1 U480 ( .A1(n369), .A2(n386), .ZN(n370) );
  NAND2_X1 U481 ( .A1(n424), .A2(n422), .ZN(n425) );
  AND2_X1 U482 ( .A1(n416), .A2(n413), .ZN(n412) );
  AND2_X1 U483 ( .A1(n725), .A2(n417), .ZN(n416) );
  BUF_X1 U484 ( .A(n653), .Z(n790) );
  INV_X1 U485 ( .A(n371), .ZN(n609) );
  XNOR2_X2 U486 ( .A(n633), .B(n603), .ZN(n777) );
  NOR2_X2 U487 ( .A1(n415), .A2(n783), .ZN(n621) );
  OR2_X2 U488 ( .A1(n583), .A2(n582), .ZN(n633) );
  NAND2_X1 U489 ( .A1(n426), .A2(n362), .ZN(n424) );
  INV_X1 U490 ( .A(n742), .ZN(n419) );
  XNOR2_X1 U491 ( .A(n742), .B(n482), .ZN(n604) );
  NOR2_X2 U492 ( .A1(n655), .A2(n654), .ZN(n372) );
  XNOR2_X1 U493 ( .A(n472), .B(n473), .ZN(n475) );
  XNOR2_X1 U494 ( .A(n375), .B(KEYINPUT34), .ZN(n542) );
  NOR2_X2 U495 ( .A1(n577), .A2(n724), .ZN(n375) );
  NAND2_X1 U496 ( .A1(n421), .A2(n425), .ZN(n377) );
  XNOR2_X2 U497 ( .A(n653), .B(n652), .ZN(n421) );
  NAND2_X1 U498 ( .A1(n377), .A2(n427), .ZN(n376) );
  NAND2_X1 U499 ( .A1(n379), .A2(n719), .ZN(n378) );
  NAND2_X1 U500 ( .A1(n421), .A2(n380), .ZN(n379) );
  NAND2_X1 U501 ( .A1(n790), .A2(n423), .ZN(n380) );
  OR2_X1 U502 ( .A1(n711), .A2(n386), .ZN(n385) );
  INV_X1 U503 ( .A(n403), .ZN(n386) );
  NAND2_X1 U504 ( .A1(n693), .A2(n388), .ZN(n387) );
  NOR2_X1 U505 ( .A1(n464), .A2(G902), .ZN(n388) );
  NAND2_X1 U506 ( .A1(n464), .A2(G902), .ZN(n390) );
  INV_X1 U507 ( .A(n464), .ZN(n392) );
  OR2_X1 U508 ( .A1(n368), .A2(n394), .ZN(n393) );
  NAND2_X1 U509 ( .A1(n370), .A2(n400), .ZN(n600) );
  AND2_X2 U510 ( .A1(n400), .A2(n399), .ZN(n398) );
  INV_X1 U511 ( .A(n448), .ZN(n402) );
  NAND2_X1 U512 ( .A1(n448), .A2(G902), .ZN(n403) );
  NAND2_X1 U513 ( .A1(n771), .A2(n412), .ZN(n408) );
  XNOR2_X1 U514 ( .A(n612), .B(n611), .ZN(n414) );
  INV_X1 U515 ( .A(KEYINPUT71), .ZN(n417) );
  INV_X1 U516 ( .A(n738), .ZN(n593) );
  INV_X1 U517 ( .A(n420), .ZN(n606) );
  NAND2_X1 U518 ( .A1(n719), .A2(n421), .ZN(n722) );
  XNOR2_X2 U519 ( .A(n432), .B(KEYINPUT45), .ZN(n653) );
  XNOR2_X2 U520 ( .A(n429), .B(n428), .ZN(n491) );
  XNOR2_X2 U521 ( .A(n469), .B(KEYINPUT3), .ZN(n429) );
  AND2_X2 U522 ( .A1(n431), .A2(n430), .ZN(n433) );
  AND2_X2 U523 ( .A1(n592), .A2(n591), .ZN(n430) );
  NAND2_X1 U524 ( .A1(n569), .A2(n570), .ZN(n431) );
  NAND2_X2 U525 ( .A1(n434), .A2(n433), .ZN(n432) );
  NAND2_X1 U526 ( .A1(n435), .A2(n563), .ZN(n434) );
  NAND2_X1 U527 ( .A1(n562), .A2(n567), .ZN(n435) );
  INV_X1 U528 ( .A(n604), .ZN(n436) );
  AND2_X1 U529 ( .A1(n437), .A2(n419), .ZN(n747) );
  INV_X1 U530 ( .A(KEYINPUT76), .ZN(n438) );
  NAND2_X1 U531 ( .A1(n556), .A2(n738), .ZN(n684) );
  XNOR2_X1 U532 ( .A(n471), .B(n470), .ZN(n472) );
  BUF_X1 U533 ( .A(n368), .Z(n714) );
  INV_X1 U534 ( .A(KEYINPUT56), .ZN(n663) );
  XNOR2_X2 U535 ( .A(G143), .B(KEYINPUT65), .ZN(n440) );
  XNOR2_X2 U536 ( .A(n440), .B(G128), .ZN(n521) );
  XNOR2_X2 U537 ( .A(n521), .B(KEYINPUT4), .ZN(n493) );
  XNOR2_X2 U538 ( .A(n493), .B(n441), .ZN(n477) );
  XNOR2_X2 U539 ( .A(n477), .B(n452), .ZN(n672) );
  XNOR2_X1 U540 ( .A(G104), .B(G110), .ZN(n442) );
  XNOR2_X1 U541 ( .A(n442), .B(G107), .ZN(n797) );
  XNOR2_X1 U542 ( .A(n797), .B(n474), .ZN(n495) );
  XOR2_X1 U543 ( .A(G146), .B(KEYINPUT79), .Z(n445) );
  INV_X2 U544 ( .A(KEYINPUT64), .ZN(n443) );
  XNOR2_X2 U545 ( .A(n443), .B(G953), .ZN(n449) );
  NAND2_X1 U546 ( .A1(n449), .A2(G227), .ZN(n444) );
  XNOR2_X1 U547 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U548 ( .A(n495), .B(n446), .ZN(n447) );
  XOR2_X1 U549 ( .A(KEYINPUT73), .B(G469), .Z(n448) );
  NAND2_X1 U550 ( .A1(n449), .A2(G234), .ZN(n451) );
  XNOR2_X1 U551 ( .A(n451), .B(n450), .ZN(n518) );
  INV_X1 U552 ( .A(n452), .ZN(n453) );
  XOR2_X1 U553 ( .A(n453), .B(KEYINPUT95), .Z(n454) );
  XOR2_X1 U554 ( .A(KEYINPUT24), .B(G110), .Z(n457) );
  XNOR2_X1 U555 ( .A(KEYINPUT96), .B(n455), .ZN(n456) );
  XNOR2_X1 U556 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U557 ( .A(G146), .B(G125), .ZN(n487) );
  XNOR2_X1 U558 ( .A(n487), .B(KEYINPUT10), .ZN(n671) );
  XNOR2_X1 U559 ( .A(n458), .B(n671), .ZN(n459) );
  INV_X1 U560 ( .A(G902), .ZN(n525) );
  XOR2_X1 U561 ( .A(KEYINPUT25), .B(KEYINPUT97), .Z(n463) );
  XNOR2_X1 U562 ( .A(G902), .B(KEYINPUT15), .ZN(n498) );
  NAND2_X1 U563 ( .A1(G234), .A2(n498), .ZN(n461) );
  XNOR2_X1 U564 ( .A(KEYINPUT20), .B(n461), .ZN(n465) );
  NAND2_X1 U565 ( .A1(n465), .A2(G217), .ZN(n462) );
  XNOR2_X1 U566 ( .A(n463), .B(n462), .ZN(n464) );
  AND2_X1 U567 ( .A1(n465), .A2(G221), .ZN(n467) );
  INV_X1 U568 ( .A(KEYINPUT21), .ZN(n466) );
  XNOR2_X1 U569 ( .A(n467), .B(n466), .ZN(n737) );
  XNOR2_X2 U570 ( .A(G116), .B(KEYINPUT88), .ZN(n469) );
  NAND2_X1 U571 ( .A1(n531), .A2(G210), .ZN(n473) );
  XNOR2_X1 U572 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U573 ( .A(n478), .B(n359), .ZN(n688) );
  INV_X1 U574 ( .A(KEYINPUT74), .ZN(n479) );
  XNOR2_X1 U575 ( .A(n479), .B(G472), .ZN(n480) );
  XNOR2_X2 U576 ( .A(n481), .B(n480), .ZN(n742) );
  INV_X1 U577 ( .A(KEYINPUT6), .ZN(n482) );
  NAND2_X1 U578 ( .A1(n449), .A2(G224), .ZN(n485) );
  XNOR2_X1 U579 ( .A(n483), .B(KEYINPUT80), .ZN(n484) );
  XNOR2_X1 U580 ( .A(n485), .B(n484), .ZN(n489) );
  XNOR2_X1 U581 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U582 ( .A(n489), .B(n488), .ZN(n492) );
  XNOR2_X1 U583 ( .A(G122), .B(KEYINPUT16), .ZN(n490) );
  XNOR2_X1 U584 ( .A(n794), .B(n492), .ZN(n497) );
  XOR2_X1 U585 ( .A(n495), .B(n494), .Z(n496) );
  XNOR2_X1 U586 ( .A(n497), .B(n496), .ZN(n655) );
  INV_X1 U587 ( .A(n498), .ZN(n654) );
  NOR2_X1 U588 ( .A1(G237), .A2(G902), .ZN(n499) );
  XNOR2_X1 U589 ( .A(KEYINPUT77), .B(n499), .ZN(n502) );
  NAND2_X1 U590 ( .A1(n502), .A2(G210), .ZN(n500) );
  NAND2_X1 U591 ( .A1(n502), .A2(G214), .ZN(n503) );
  XNOR2_X1 U592 ( .A(n503), .B(KEYINPUT91), .ZN(n622) );
  XNOR2_X1 U593 ( .A(n505), .B(KEYINPUT14), .ZN(n507) );
  NAND2_X1 U594 ( .A1(G952), .A2(n507), .ZN(n756) );
  NOR2_X1 U595 ( .A1(G953), .A2(n756), .ZN(n506) );
  XNOR2_X1 U596 ( .A(n506), .B(KEYINPUT92), .ZN(n597) );
  NAND2_X1 U597 ( .A1(G902), .A2(n507), .ZN(n594) );
  XNOR2_X1 U598 ( .A(G898), .B(KEYINPUT93), .ZN(n788) );
  NAND2_X1 U599 ( .A1(G953), .A2(n788), .ZN(n799) );
  NOR2_X1 U600 ( .A1(n594), .A2(n799), .ZN(n508) );
  OR2_X1 U601 ( .A1(n597), .A2(n508), .ZN(n509) );
  XNOR2_X1 U602 ( .A(KEYINPUT85), .B(KEYINPUT0), .ZN(n510) );
  XNOR2_X2 U603 ( .A(n511), .B(n510), .ZN(n572) );
  XNOR2_X1 U604 ( .A(n572), .B(n512), .ZN(n577) );
  XNOR2_X1 U605 ( .A(n513), .B(G116), .ZN(n517) );
  XNOR2_X1 U606 ( .A(n515), .B(n514), .ZN(n516) );
  XOR2_X1 U607 ( .A(n517), .B(n516), .Z(n520) );
  NAND2_X1 U608 ( .A1(G217), .A2(n518), .ZN(n519) );
  XNOR2_X1 U609 ( .A(n520), .B(n519), .ZN(n524) );
  BUF_X1 U610 ( .A(n521), .Z(n522) );
  INV_X1 U611 ( .A(n522), .ZN(n523) );
  XNOR2_X1 U612 ( .A(n524), .B(n523), .ZN(n697) );
  NAND2_X1 U613 ( .A1(n697), .A2(n525), .ZN(n527) );
  INV_X1 U614 ( .A(G478), .ZN(n526) );
  XNOR2_X1 U615 ( .A(n527), .B(n526), .ZN(n580) );
  INV_X1 U616 ( .A(n580), .ZN(n583) );
  XNOR2_X1 U617 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U618 ( .A(n671), .B(n530), .ZN(n538) );
  NAND2_X1 U619 ( .A1(n531), .A2(G214), .ZN(n532) );
  XNOR2_X1 U620 ( .A(n532), .B(KEYINPUT11), .ZN(n536) );
  XNOR2_X1 U621 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U622 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U623 ( .A(n538), .B(n537), .ZN(n703) );
  OR2_X1 U624 ( .A1(n703), .A2(G902), .ZN(n541) );
  INV_X1 U625 ( .A(KEYINPUT13), .ZN(n539) );
  XNOR2_X1 U626 ( .A(n539), .B(G475), .ZN(n540) );
  XNOR2_X1 U627 ( .A(n541), .B(n540), .ZN(n579) );
  AND2_X1 U628 ( .A1(n583), .A2(n579), .ZN(n618) );
  NAND2_X1 U629 ( .A1(n542), .A2(n618), .ZN(n544) );
  INV_X1 U630 ( .A(KEYINPUT35), .ZN(n543) );
  XNOR2_X2 U631 ( .A(n544), .B(n543), .ZN(n685) );
  INV_X1 U632 ( .A(KEYINPUT84), .ZN(n545) );
  NAND2_X1 U633 ( .A1(n685), .A2(n545), .ZN(n546) );
  INV_X1 U634 ( .A(KEYINPUT44), .ZN(n565) );
  NAND2_X1 U635 ( .A1(n546), .A2(n565), .ZN(n561) );
  OR2_X1 U636 ( .A1(n583), .A2(n579), .ZN(n548) );
  INV_X1 U637 ( .A(KEYINPUT104), .ZN(n547) );
  XNOR2_X1 U638 ( .A(n548), .B(n547), .ZN(n625) );
  AND2_X1 U639 ( .A1(n625), .A2(n383), .ZN(n549) );
  NAND2_X1 U640 ( .A1(n572), .A2(n549), .ZN(n551) );
  XNOR2_X1 U641 ( .A(KEYINPUT75), .B(KEYINPUT22), .ZN(n550) );
  BUF_X1 U642 ( .A(n552), .Z(n553) );
  INV_X1 U643 ( .A(n553), .ZN(n647) );
  NAND2_X1 U644 ( .A1(n587), .A2(n742), .ZN(n555) );
  AND2_X1 U645 ( .A1(n604), .A2(n738), .ZN(n557) );
  AND2_X1 U646 ( .A1(n553), .A2(n557), .ZN(n558) );
  NAND2_X1 U647 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U648 ( .A(n560), .B(KEYINPUT32), .ZN(n668) );
  NAND2_X1 U649 ( .A1(n684), .A2(n668), .ZN(n564) );
  NAND2_X1 U650 ( .A1(n561), .A2(n564), .ZN(n562) );
  INV_X1 U651 ( .A(KEYINPUT67), .ZN(n567) );
  NAND2_X1 U652 ( .A1(KEYINPUT67), .A2(KEYINPUT44), .ZN(n563) );
  INV_X1 U653 ( .A(n564), .ZN(n570) );
  AND2_X1 U654 ( .A1(n565), .A2(KEYINPUT84), .ZN(n566) );
  NAND2_X1 U655 ( .A1(n685), .A2(n566), .ZN(n568) );
  NAND2_X1 U656 ( .A1(n568), .A2(n567), .ZN(n569) );
  INV_X1 U657 ( .A(n685), .ZN(n571) );
  NAND2_X1 U658 ( .A1(n571), .A2(KEYINPUT44), .ZN(n592) );
  BUF_X1 U659 ( .A(n572), .Z(n573) );
  NAND2_X1 U660 ( .A1(n747), .A2(n573), .ZN(n575) );
  INV_X1 U661 ( .A(KEYINPUT31), .ZN(n574) );
  XNOR2_X1 U662 ( .A(n575), .B(n574), .ZN(n780) );
  NAND2_X1 U663 ( .A1(n734), .A2(n600), .ZN(n615) );
  OR2_X1 U664 ( .A1(n615), .A2(n419), .ZN(n576) );
  OR2_X1 U665 ( .A1(n577), .A2(n576), .ZN(n767) );
  NAND2_X1 U666 ( .A1(n780), .A2(n767), .ZN(n578) );
  XNOR2_X1 U667 ( .A(n578), .B(KEYINPUT98), .ZN(n586) );
  XNOR2_X1 U668 ( .A(n579), .B(KEYINPUT100), .ZN(n581) );
  OR2_X1 U669 ( .A1(n580), .A2(n581), .ZN(n781) );
  XNOR2_X1 U670 ( .A(n781), .B(KEYINPUT102), .ZN(n643) );
  INV_X1 U671 ( .A(n581), .ZN(n582) );
  NAND2_X1 U672 ( .A1(n643), .A2(n633), .ZN(n585) );
  INV_X1 U673 ( .A(KEYINPUT103), .ZN(n584) );
  XNOR2_X1 U674 ( .A(n585), .B(n584), .ZN(n725) );
  NAND2_X1 U675 ( .A1(n586), .A2(n725), .ZN(n590) );
  NAND2_X1 U676 ( .A1(n587), .A2(n604), .ZN(n588) );
  XNOR2_X1 U677 ( .A(n588), .B(KEYINPUT83), .ZN(n589) );
  NAND2_X1 U678 ( .A1(n589), .A2(n593), .ZN(n669) );
  AND2_X1 U679 ( .A1(n590), .A2(n669), .ZN(n591) );
  INV_X1 U680 ( .A(KEYINPUT2), .ZN(n652) );
  NOR2_X1 U681 ( .A1(G900), .A2(n594), .ZN(n595) );
  INV_X1 U682 ( .A(n449), .ZN(n661) );
  AND2_X1 U683 ( .A1(n595), .A2(n661), .ZN(n596) );
  OR2_X1 U684 ( .A1(n597), .A2(n596), .ZN(n616) );
  XNOR2_X1 U685 ( .A(KEYINPUT28), .B(n598), .ZN(n599) );
  AND2_X1 U686 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U687 ( .A(n601), .B(KEYINPUT106), .ZN(n627) );
  INV_X1 U688 ( .A(KEYINPUT105), .ZN(n603) );
  NOR2_X1 U689 ( .A1(n604), .A2(n777), .ZN(n605) );
  NAND2_X1 U690 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U691 ( .A1(n622), .A2(n607), .ZN(n608) );
  AND2_X1 U692 ( .A1(n608), .A2(n616), .ZN(n648) );
  INV_X1 U693 ( .A(n609), .ZN(n610) );
  NAND2_X1 U694 ( .A1(n648), .A2(n610), .ZN(n612) );
  INV_X1 U695 ( .A(KEYINPUT36), .ZN(n611) );
  NOR2_X1 U696 ( .A1(n742), .A2(n622), .ZN(n613) );
  AND2_X1 U697 ( .A1(n617), .A2(n616), .ZN(n630) );
  INV_X1 U698 ( .A(n618), .ZN(n619) );
  NOR2_X1 U699 ( .A1(n619), .A2(n609), .ZN(n620) );
  AND2_X1 U700 ( .A1(n630), .A2(n620), .ZN(n665) );
  XNOR2_X1 U701 ( .A(n621), .B(KEYINPUT72), .ZN(n640) );
  NAND2_X1 U702 ( .A1(n728), .A2(n504), .ZN(n624) );
  INV_X1 U703 ( .A(KEYINPUT107), .ZN(n623) );
  XNOR2_X1 U704 ( .A(n624), .B(n623), .ZN(n726) );
  INV_X1 U705 ( .A(n625), .ZN(n729) );
  OR2_X1 U706 ( .A1(n726), .A2(n729), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n627), .A2(n750), .ZN(n629) );
  INV_X1 U708 ( .A(KEYINPUT42), .ZN(n628) );
  XNOR2_X1 U709 ( .A(n629), .B(n628), .ZN(n670) );
  NAND2_X1 U710 ( .A1(n630), .A2(n728), .ZN(n632) );
  INV_X1 U711 ( .A(KEYINPUT39), .ZN(n631) );
  XNOR2_X1 U712 ( .A(n632), .B(n631), .ZN(n644) );
  INV_X1 U713 ( .A(KEYINPUT40), .ZN(n634) );
  INV_X1 U714 ( .A(KEYINPUT82), .ZN(n636) );
  XNOR2_X1 U715 ( .A(n636), .B(KEYINPUT46), .ZN(n637) );
  XNOR2_X1 U716 ( .A(n638), .B(n637), .ZN(n639) );
  INV_X1 U717 ( .A(KEYINPUT48), .ZN(n641) );
  OR2_X1 U718 ( .A1(n644), .A2(n643), .ZN(n646) );
  INV_X1 U719 ( .A(KEYINPUT108), .ZN(n645) );
  XNOR2_X1 U720 ( .A(n646), .B(n645), .ZN(n805) );
  NAND2_X1 U721 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U722 ( .A(n649), .B(KEYINPUT43), .ZN(n650) );
  AND2_X1 U723 ( .A1(n609), .A2(n650), .ZN(n666) );
  NOR2_X1 U724 ( .A1(n805), .A2(n666), .ZN(n651) );
  INV_X1 U725 ( .A(n720), .ZN(n719) );
  NAND2_X1 U726 ( .A1(n366), .A2(G210), .ZN(n659) );
  XNOR2_X1 U727 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n656) );
  XNOR2_X1 U728 ( .A(n659), .B(n658), .ZN(n662) );
  INV_X1 U729 ( .A(G952), .ZN(n660) );
  NAND2_X1 U730 ( .A1(n662), .A2(n706), .ZN(n664) );
  XNOR2_X1 U731 ( .A(n664), .B(n663), .ZN(G51) );
  XOR2_X1 U732 ( .A(G143), .B(n665), .Z(G45) );
  XOR2_X1 U733 ( .A(G140), .B(n666), .Z(G42) );
  NOR2_X1 U734 ( .A1(n767), .A2(n777), .ZN(n667) );
  XOR2_X1 U735 ( .A(G104), .B(n667), .Z(G6) );
  XNOR2_X1 U736 ( .A(n668), .B(G119), .ZN(G21) );
  XNOR2_X1 U737 ( .A(n367), .B(G101), .ZN(G3) );
  XOR2_X1 U738 ( .A(G137), .B(n670), .Z(G39) );
  XNOR2_X1 U739 ( .A(n671), .B(KEYINPUT125), .ZN(n674) );
  BUF_X1 U740 ( .A(n672), .Z(n673) );
  XOR2_X1 U741 ( .A(n674), .B(n673), .Z(n677) );
  XOR2_X1 U742 ( .A(KEYINPUT126), .B(n677), .Z(n675) );
  XOR2_X1 U743 ( .A(n675), .B(n720), .Z(n676) );
  NAND2_X1 U744 ( .A1(n676), .A2(n449), .ZN(n683) );
  INV_X1 U745 ( .A(n677), .ZN(n678) );
  XOR2_X1 U746 ( .A(G227), .B(n678), .Z(n679) );
  NAND2_X1 U747 ( .A1(n679), .A2(G900), .ZN(n680) );
  XOR2_X1 U748 ( .A(KEYINPUT127), .B(n680), .Z(n681) );
  NAND2_X1 U749 ( .A1(G953), .A2(n681), .ZN(n682) );
  NAND2_X1 U750 ( .A1(n683), .A2(n682), .ZN(G72) );
  XNOR2_X1 U751 ( .A(n684), .B(G110), .ZN(G12) );
  BUF_X1 U752 ( .A(n685), .Z(n686) );
  XNOR2_X1 U753 ( .A(n686), .B(G122), .ZN(G24) );
  NAND2_X1 U754 ( .A1(n366), .A2(G472), .ZN(n690) );
  XNOR2_X1 U755 ( .A(KEYINPUT109), .B(KEYINPUT62), .ZN(n687) );
  XNOR2_X1 U756 ( .A(n690), .B(n689), .ZN(n691) );
  NAND2_X1 U757 ( .A1(n691), .A2(n706), .ZN(n692) );
  XNOR2_X1 U758 ( .A(n692), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U759 ( .A1(n701), .A2(G217), .ZN(n694) );
  XNOR2_X1 U760 ( .A(n694), .B(n693), .ZN(n695) );
  NAND2_X1 U761 ( .A1(n695), .A2(n706), .ZN(n696) );
  XNOR2_X1 U762 ( .A(n696), .B(KEYINPUT121), .ZN(G66) );
  BUF_X1 U763 ( .A(n701), .Z(n710) );
  NAND2_X1 U764 ( .A1(n710), .A2(G478), .ZN(n699) );
  XOR2_X1 U765 ( .A(KEYINPUT120), .B(n697), .Z(n698) );
  XNOR2_X1 U766 ( .A(n699), .B(n698), .ZN(n700) );
  INV_X1 U767 ( .A(n706), .ZN(n717) );
  NOR2_X1 U768 ( .A1(n700), .A2(n717), .ZN(G63) );
  NAND2_X1 U769 ( .A1(n366), .A2(G475), .ZN(n705) );
  XOR2_X1 U770 ( .A(KEYINPUT69), .B(KEYINPUT59), .Z(n702) );
  XNOR2_X1 U771 ( .A(n705), .B(n704), .ZN(n707) );
  NAND2_X1 U772 ( .A1(n707), .A2(n706), .ZN(n709) );
  XNOR2_X1 U773 ( .A(KEYINPUT119), .B(KEYINPUT60), .ZN(n708) );
  XNOR2_X1 U774 ( .A(n709), .B(n708), .ZN(G60) );
  NAND2_X1 U775 ( .A1(n710), .A2(G469), .ZN(n716) );
  XOR2_X1 U776 ( .A(KEYINPUT118), .B(KEYINPUT57), .Z(n712) );
  XNOR2_X1 U777 ( .A(n712), .B(KEYINPUT58), .ZN(n713) );
  XNOR2_X1 U778 ( .A(n714), .B(n713), .ZN(n715) );
  XNOR2_X1 U779 ( .A(n716), .B(n715), .ZN(n718) );
  NOR2_X1 U780 ( .A1(n718), .A2(n717), .ZN(G54) );
  NAND2_X1 U781 ( .A1(n720), .A2(KEYINPUT2), .ZN(n721) );
  NAND2_X1 U782 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U783 ( .A(n723), .B(KEYINPUT81), .ZN(n765) );
  XNOR2_X1 U784 ( .A(KEYINPUT116), .B(KEYINPUT52), .ZN(n755) );
  INV_X1 U785 ( .A(n725), .ZN(n727) );
  NOR2_X1 U786 ( .A1(n727), .A2(n726), .ZN(n732) );
  NOR2_X1 U787 ( .A1(n728), .A2(n504), .ZN(n730) );
  NOR2_X1 U788 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U789 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U790 ( .A1(n760), .A2(n733), .ZN(n753) );
  NOR2_X1 U791 ( .A1(n734), .A2(n553), .ZN(n736) );
  XNOR2_X1 U792 ( .A(KEYINPUT114), .B(KEYINPUT50), .ZN(n735) );
  XNOR2_X1 U793 ( .A(n736), .B(n735), .ZN(n745) );
  NAND2_X1 U794 ( .A1(n738), .A2(n737), .ZN(n741) );
  XNOR2_X1 U795 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n739) );
  XNOR2_X1 U796 ( .A(n739), .B(KEYINPUT49), .ZN(n740) );
  XNOR2_X1 U797 ( .A(n741), .B(n740), .ZN(n743) );
  NAND2_X1 U798 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U799 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U800 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U801 ( .A(n748), .B(KEYINPUT51), .ZN(n749) );
  XNOR2_X1 U802 ( .A(KEYINPUT115), .B(n749), .ZN(n751) );
  INV_X1 U803 ( .A(n750), .ZN(n759) );
  NOR2_X1 U804 ( .A1(n751), .A2(n759), .ZN(n752) );
  NOR2_X1 U805 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U806 ( .A(n755), .B(n754), .ZN(n757) );
  NOR2_X1 U807 ( .A1(n757), .A2(n756), .ZN(n758) );
  XOR2_X1 U808 ( .A(KEYINPUT117), .B(n758), .Z(n763) );
  OR2_X1 U809 ( .A1(n760), .A2(n759), .ZN(n761) );
  INV_X1 U810 ( .A(G953), .ZN(n789) );
  NAND2_X1 U811 ( .A1(n761), .A2(n789), .ZN(n762) );
  NOR2_X1 U812 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U813 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U814 ( .A(KEYINPUT53), .B(n766), .Z(G75) );
  NOR2_X1 U815 ( .A1(n767), .A2(n781), .ZN(n769) );
  XNOR2_X1 U816 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n768) );
  XNOR2_X1 U817 ( .A(n769), .B(n768), .ZN(n770) );
  XNOR2_X1 U818 ( .A(G107), .B(n770), .ZN(G9) );
  XOR2_X1 U819 ( .A(G128), .B(KEYINPUT29), .Z(n774) );
  INV_X1 U820 ( .A(n781), .ZN(n772) );
  NAND2_X1 U821 ( .A1(n771), .A2(n772), .ZN(n773) );
  XNOR2_X1 U822 ( .A(n774), .B(n773), .ZN(G30) );
  INV_X1 U823 ( .A(n777), .ZN(n775) );
  NAND2_X1 U824 ( .A1(n771), .A2(n775), .ZN(n776) );
  XNOR2_X1 U825 ( .A(n776), .B(G146), .ZN(G48) );
  NOR2_X1 U826 ( .A1(n777), .A2(n780), .ZN(n778) );
  XOR2_X1 U827 ( .A(KEYINPUT110), .B(n778), .Z(n779) );
  XNOR2_X1 U828 ( .A(G113), .B(n779), .ZN(G15) );
  NOR2_X1 U829 ( .A1(n781), .A2(n780), .ZN(n782) );
  XOR2_X1 U830 ( .A(G116), .B(n782), .Z(G18) );
  XOR2_X1 U831 ( .A(KEYINPUT111), .B(KEYINPUT37), .Z(n785) );
  XNOR2_X1 U832 ( .A(G125), .B(n783), .ZN(n784) );
  XNOR2_X1 U833 ( .A(n785), .B(n784), .ZN(G27) );
  NAND2_X1 U834 ( .A1(G953), .A2(G224), .ZN(n786) );
  XOR2_X1 U835 ( .A(KEYINPUT61), .B(n786), .Z(n787) );
  NOR2_X1 U836 ( .A1(n788), .A2(n787), .ZN(n793) );
  NAND2_X1 U837 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U838 ( .A(KEYINPUT122), .B(n791), .Z(n792) );
  NOR2_X1 U839 ( .A1(n793), .A2(n792), .ZN(n803) );
  BUF_X1 U840 ( .A(n794), .Z(n795) );
  XNOR2_X1 U841 ( .A(G101), .B(KEYINPUT123), .ZN(n796) );
  XNOR2_X1 U842 ( .A(n797), .B(n796), .ZN(n798) );
  XNOR2_X1 U843 ( .A(n795), .B(n798), .ZN(n800) );
  NAND2_X1 U844 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U845 ( .A(n801), .B(KEYINPUT124), .ZN(n802) );
  XNOR2_X1 U846 ( .A(n803), .B(n802), .ZN(G69) );
  XOR2_X1 U847 ( .A(G131), .B(n804), .Z(G33) );
  XOR2_X1 U848 ( .A(G134), .B(n805), .Z(G36) );
endmodule

