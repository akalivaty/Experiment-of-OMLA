//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1227, new_n1228, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G20), .ZN(new_n218));
  INV_X1    g0018(.A(new_n202), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT65), .Z(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n212), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n215), .B1(new_n218), .B2(new_n220), .C1(new_n227), .C2(KEYINPUT1), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  NAND2_X1  g0044(.A1(G33), .A2(G41), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n217), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(G33), .A2(G97), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  AND2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G1698), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n248), .B1(new_n253), .B2(G232), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G226), .A3(new_n252), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n246), .B1(new_n254), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT66), .B(G45), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n209), .A2(G274), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G45), .ZN(new_n267));
  AOI21_X1  g0067(.A(G1), .B1(new_n263), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n216), .B1(KEYINPUT67), .B2(new_n245), .ZN(new_n269));
  OR2_X1    g0069(.A1(new_n245), .A2(KEYINPUT67), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G238), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n266), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(KEYINPUT13), .B1(new_n261), .B2(new_n274), .ZN(new_n275));
  AND2_X1   g0075(.A1(new_n264), .A2(new_n265), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n276), .B1(G238), .B2(new_n271), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n259), .A2(G1698), .ZN(new_n278));
  INV_X1    g0078(.A(G232), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n260), .B(new_n247), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n246), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT13), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n277), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n275), .A2(new_n284), .A3(KEYINPUT69), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT69), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n286), .B(KEYINPUT13), .C1(new_n261), .C2(new_n274), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n285), .A2(G169), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(KEYINPUT14), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT70), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n284), .B(new_n290), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n275), .A2(G179), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT14), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n285), .A2(new_n295), .A3(G169), .A4(new_n287), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(KEYINPUT74), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(KEYINPUT74), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n294), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n216), .ZN(new_n302));
  NOR2_X1   g0102(.A1(G20), .A2(G33), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G50), .ZN(new_n305));
  OAI22_X1  g0105(.A1(new_n304), .A2(new_n305), .B1(new_n210), .B2(G68), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n210), .A2(G33), .ZN(new_n307));
  INV_X1    g0107(.A(G77), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n302), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT72), .ZN(new_n311));
  OR2_X1    g0111(.A1(new_n311), .A2(KEYINPUT11), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(KEYINPUT11), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n314));
  OAI22_X1  g0114(.A1(new_n314), .A2(G68), .B1(KEYINPUT73), .B2(KEYINPUT12), .ZN(new_n315));
  NAND2_X1  g0115(.A1(KEYINPUT73), .A2(KEYINPUT12), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(new_n316), .ZN(new_n318));
  INV_X1    g0118(.A(new_n314), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(new_n302), .ZN(new_n320));
  INV_X1    g0120(.A(G68), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n321), .B1(new_n209), .B2(G20), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n317), .A2(new_n318), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n312), .A2(new_n313), .A3(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n300), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n285), .A2(G200), .A3(new_n287), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n275), .A2(G190), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n291), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT71), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT71), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n291), .A2(new_n332), .A3(new_n329), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n328), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n302), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n203), .A2(G20), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT8), .B(G58), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n307), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n338), .A2(new_n339), .B1(G150), .B2(new_n303), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n335), .B1(new_n336), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n209), .A2(G20), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n320), .A2(G50), .A3(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(G50), .B2(new_n314), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  OR2_X1    g0145(.A1(new_n345), .A2(KEYINPUT9), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n259), .A2(G222), .A3(new_n252), .ZN(new_n347));
  INV_X1    g0147(.A(G223), .ZN(new_n348));
  OAI221_X1 g0148(.A(new_n347), .B1(new_n308), .B2(new_n259), .C1(new_n348), .C2(new_n278), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n281), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n276), .B1(G226), .B2(new_n271), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(G200), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n350), .A2(G190), .A3(new_n351), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n345), .A2(KEYINPUT9), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n346), .A2(new_n353), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  XNOR2_X1  g0156(.A(new_n356), .B(KEYINPUT10), .ZN(new_n357));
  INV_X1    g0157(.A(G169), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n345), .B1(new_n352), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G179), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n350), .A2(new_n360), .A3(new_n351), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n357), .A2(new_n363), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n338), .A2(new_n303), .B1(G20), .B2(G77), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT15), .B(G87), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n339), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n335), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n320), .A2(G77), .A3(new_n342), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(G77), .B2(new_n314), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n276), .B1(G244), .B2(new_n271), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n259), .A2(G232), .A3(new_n252), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n251), .A2(G107), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n375), .B(new_n376), .C1(new_n278), .C2(new_n273), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n281), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  OAI211_X1 g0180(.A(KEYINPUT68), .B(new_n373), .C1(new_n380), .C2(G169), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT68), .ZN(new_n382));
  AOI21_X1  g0182(.A(G169), .B1(new_n374), .B2(new_n378), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n382), .B1(new_n383), .B2(new_n372), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n380), .A2(new_n360), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n381), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n373), .B1(new_n380), .B2(G190), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n379), .A2(G200), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NOR4_X1   g0190(.A1(new_n326), .A2(new_n334), .A3(new_n364), .A4(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(G159), .ZN(new_n392));
  NOR3_X1   g0192(.A1(new_n392), .A2(G20), .A3(G33), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G58), .A2(G68), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT76), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(KEYINPUT76), .A2(G58), .A3(G68), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n219), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n393), .B1(new_n398), .B2(G20), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n258), .A2(new_n210), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT7), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT75), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n256), .ZN(new_n404));
  NAND2_X1  g0204(.A1(KEYINPUT75), .A2(G33), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n255), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n401), .B1(new_n400), .B2(new_n250), .ZN(new_n408));
  AND2_X1   g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n399), .B1(new_n409), .B2(new_n321), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT16), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI211_X1 g0212(.A(new_n411), .B(new_n393), .C1(new_n398), .C2(G20), .ZN(new_n413));
  XNOR2_X1  g0213(.A(KEYINPUT75), .B(G33), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n250), .B1(new_n414), .B2(KEYINPUT3), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n401), .B1(new_n415), .B2(new_n210), .ZN(new_n416));
  AND2_X1   g0216(.A1(KEYINPUT75), .A2(G33), .ZN(new_n417));
  NOR2_X1   g0217(.A1(KEYINPUT75), .A2(G33), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT3), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n419), .A2(new_n401), .A3(new_n210), .A4(new_n257), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(G68), .ZN(new_n421));
  OAI211_X1 g0221(.A(KEYINPUT77), .B(new_n413), .C1(new_n416), .C2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n419), .A2(new_n210), .A3(new_n257), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT7), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n425), .A2(G68), .A3(new_n420), .ZN(new_n426));
  AOI21_X1  g0226(.A(KEYINPUT77), .B1(new_n426), .B2(new_n413), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n412), .B(new_n302), .C1(new_n423), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n338), .A2(new_n342), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n335), .A2(new_n314), .ZN(new_n430));
  OAI22_X1  g0230(.A1(new_n429), .A2(new_n430), .B1(new_n314), .B2(new_n338), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  OR2_X1    g0232(.A1(G223), .A2(G1698), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(G226), .B2(new_n252), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(new_n257), .B2(new_n419), .ZN(new_n435));
  INV_X1    g0235(.A(G87), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n256), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n281), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n271), .A2(G232), .B1(new_n264), .B2(new_n265), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(G200), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(G190), .B2(new_n440), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n428), .A2(new_n432), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT17), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n428), .A2(KEYINPUT17), .A3(new_n443), .A4(new_n432), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT78), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n440), .A2(G169), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n438), .A2(G179), .A3(new_n439), .ZN(new_n452));
  AND2_X1   g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n453), .B1(new_n428), .B2(new_n432), .ZN(new_n454));
  XNOR2_X1  g0254(.A(new_n454), .B(KEYINPUT18), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n446), .A2(KEYINPUT78), .A3(new_n447), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n450), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n391), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  AOI211_X1 g0260(.A(new_n302), .B(new_n319), .C1(new_n209), .C2(G33), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT25), .B1(new_n319), .B2(new_n206), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n319), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n461), .A2(G107), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n206), .A2(G20), .ZN(new_n466));
  XNOR2_X1  g0266(.A(new_n466), .B(KEYINPUT23), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT84), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n417), .A2(new_n418), .ZN(new_n470));
  INV_X1    g0270(.A(G116), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n469), .B1(new_n472), .B2(new_n210), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n414), .A2(new_n210), .A3(G116), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(KEYINPUT84), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n468), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n255), .B1(new_n404), .B2(new_n405), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n210), .B(G87), .C1(new_n477), .C2(new_n250), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT83), .ZN(new_n479));
  AOI21_X1  g0279(.A(G20), .B1(new_n419), .B2(new_n257), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT83), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n480), .A2(new_n481), .A3(G87), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n479), .A2(new_n482), .A3(KEYINPUT22), .ZN(new_n483));
  NOR4_X1   g0283(.A1(new_n251), .A2(KEYINPUT22), .A3(G20), .A4(new_n436), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n476), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT85), .ZN(new_n487));
  OAI21_X1  g0287(.A(KEYINPUT24), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(KEYINPUT22), .B1(new_n478), .B2(KEYINPUT83), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n481), .B1(new_n480), .B2(G87), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n485), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n476), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(new_n487), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT24), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT22), .ZN(new_n497));
  AOI211_X1 g0297(.A(G20), .B(new_n436), .C1(new_n419), .C2(new_n257), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n497), .B1(new_n498), .B2(new_n481), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n484), .B1(new_n499), .B2(new_n479), .ZN(new_n500));
  OAI211_X1 g0300(.A(KEYINPUT85), .B(new_n496), .C1(new_n500), .C2(new_n476), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n302), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n465), .B1(new_n495), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(G257), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G1698), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(G250), .B2(G1698), .ZN(new_n506));
  INV_X1    g0306(.A(G294), .ZN(new_n507));
  OAI22_X1  g0307(.A1(new_n415), .A2(new_n506), .B1(new_n507), .B2(new_n470), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n281), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n269), .A2(new_n270), .ZN(new_n510));
  XNOR2_X1  g0310(.A(KEYINPUT5), .B(G41), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n267), .A2(G1), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n510), .A2(G274), .A3(new_n511), .A4(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n512), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n510), .A2(new_n514), .A3(G264), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n509), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(KEYINPUT86), .A3(G169), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n360), .B2(new_n516), .ZN(new_n518));
  AOI21_X1  g0318(.A(KEYINPUT86), .B1(new_n516), .B2(G169), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n503), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n465), .ZN(new_n523));
  OAI21_X1  g0323(.A(KEYINPUT85), .B1(new_n500), .B2(new_n476), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n524), .A2(KEYINPUT24), .A3(new_n493), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n487), .B1(new_n491), .B2(new_n492), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n335), .B1(new_n526), .B2(new_n496), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n523), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(G190), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n516), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n530), .B1(G200), .B2(new_n516), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n522), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT81), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n535), .A2(KEYINPUT19), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT19), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n537), .A2(KEYINPUT81), .ZN(new_n538));
  OAI22_X1  g0338(.A1(new_n536), .A2(new_n538), .B1(new_n307), .B2(new_n205), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n436), .A2(new_n205), .A3(new_n206), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n247), .A2(new_n210), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n537), .A2(KEYINPUT81), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n535), .A2(KEYINPUT19), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n540), .A2(new_n541), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n210), .B(G68), .C1(new_n477), .C2(new_n250), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n335), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n367), .A2(new_n314), .ZN(new_n548));
  OAI21_X1  g0348(.A(KEYINPUT82), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI211_X1 g0349(.A(G20), .B(new_n321), .C1(new_n419), .C2(new_n257), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n539), .A2(new_n544), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n302), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT82), .ZN(new_n553));
  INV_X1    g0353(.A(new_n548), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n461), .A2(new_n367), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n273), .A2(new_n252), .ZN(new_n559));
  INV_X1    g0359(.A(G244), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G1698), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n562), .B1(new_n419), .B2(new_n257), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n281), .B1(new_n563), .B2(new_n472), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n512), .A2(G274), .ZN(new_n565));
  INV_X1    g0365(.A(G250), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n565), .B1(new_n512), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n510), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n358), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(G179), .B2(new_n569), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n558), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n461), .A2(G87), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n564), .A2(G190), .A3(new_n568), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n441), .B1(new_n564), .B2(new_n568), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n556), .A2(new_n574), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n461), .A2(G116), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n319), .A2(new_n471), .ZN(new_n581));
  NAND2_X1  g0381(.A1(G33), .A2(G283), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT80), .ZN(new_n583));
  XNOR2_X1  g0383(.A(new_n582), .B(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(G20), .B1(new_n256), .B2(G97), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n301), .A2(new_n216), .B1(G20), .B2(new_n471), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n586), .A2(KEYINPUT20), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT20), .B1(new_n586), .B2(new_n587), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n580), .B(new_n581), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n510), .A2(new_n514), .A3(G270), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n513), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n504), .A2(new_n252), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(G264), .B2(new_n252), .ZN(new_n595));
  INV_X1    g0395(.A(G303), .ZN(new_n596));
  OAI22_X1  g0396(.A1(new_n415), .A2(new_n595), .B1(new_n596), .B2(new_n259), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n281), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G200), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n591), .B(new_n600), .C1(new_n529), .C2(new_n599), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n590), .A2(G169), .A3(new_n599), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT21), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n590), .A2(new_n599), .A3(KEYINPUT21), .A4(G169), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n599), .A2(new_n360), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n590), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n601), .A2(new_n604), .A3(new_n605), .A4(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n510), .A2(new_n514), .A3(G257), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n513), .A2(new_n609), .ZN(new_n610));
  OAI211_X1 g0410(.A(G250), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n611));
  AND2_X1   g0411(.A1(KEYINPUT4), .A2(G244), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n252), .B(new_n612), .C1(new_n249), .C2(new_n250), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n584), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n419), .A2(new_n257), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n615), .A2(G244), .A3(new_n252), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT4), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n614), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n610), .B1(new_n618), .B2(new_n246), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(G200), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n303), .A2(G77), .ZN(new_n621));
  XNOR2_X1  g0421(.A(new_n621), .B(KEYINPUT79), .ZN(new_n622));
  NAND2_X1  g0422(.A1(G97), .A2(G107), .ZN(new_n623));
  AOI21_X1  g0423(.A(KEYINPUT6), .B1(new_n207), .B2(new_n623), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n206), .A2(KEYINPUT6), .A3(G97), .ZN(new_n625));
  OAI21_X1  g0425(.A(G20), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n206), .B1(new_n407), .B2(new_n408), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n302), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n314), .A2(G97), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n630), .B1(new_n461), .B2(G97), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n620), .B(new_n633), .C1(new_n529), .C2(new_n619), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n252), .A2(G244), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n617), .B1(new_n415), .B2(new_n635), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n584), .A2(new_n611), .A3(new_n613), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n246), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n513), .A2(new_n609), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n358), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n610), .B(new_n360), .C1(new_n618), .C2(new_n246), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(new_n641), .A3(new_n632), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n634), .A2(new_n642), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n579), .A2(new_n608), .A3(new_n643), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n460), .A2(new_n534), .A3(new_n644), .ZN(G372));
  NAND2_X1  g0445(.A1(new_n331), .A2(new_n333), .ZN(new_n646));
  INV_X1    g0446(.A(new_n328), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n386), .ZN(new_n649));
  INV_X1    g0449(.A(new_n299), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n289), .B(new_n293), .C1(new_n650), .C2(new_n297), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n648), .A2(new_n649), .B1(new_n651), .B2(new_n324), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n446), .A2(KEYINPUT78), .A3(new_n447), .ZN(new_n653));
  AOI21_X1  g0453(.A(KEYINPUT78), .B1(new_n446), .B2(new_n447), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n455), .B1(new_n652), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n362), .B1(new_n657), .B2(new_n357), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n503), .A2(KEYINPUT87), .A3(new_n521), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT87), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n528), .B2(new_n520), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n659), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n579), .A2(new_n643), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n532), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT89), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n640), .A2(new_n641), .A3(new_n632), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n549), .A2(new_n555), .B1(new_n367), .B2(new_n461), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n578), .B(new_n667), .C1(new_n668), .C2(new_n571), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT26), .ZN(new_n670));
  XOR2_X1   g0470(.A(KEYINPUT88), .B(KEYINPUT26), .Z(new_n671));
  NAND4_X1  g0471(.A1(new_n573), .A2(new_n667), .A3(new_n578), .A4(new_n671), .ZN(new_n672));
  AND4_X1   g0472(.A1(new_n666), .A2(new_n670), .A3(new_n573), .A4(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n668), .A2(new_n571), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n674), .B1(new_n669), .B2(KEYINPUT26), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n666), .B1(new_n675), .B2(new_n672), .ZN(new_n676));
  OAI22_X1  g0476(.A1(new_n663), .A2(new_n665), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n658), .B1(new_n678), .B2(new_n459), .ZN(G369));
  NAND3_X1  g0479(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G213), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT90), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G343), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n590), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT91), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n659), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n608), .B2(new_n688), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G330), .ZN(new_n691));
  XOR2_X1   g0491(.A(new_n691), .B(KEYINPUT92), .Z(new_n692));
  NOR2_X1   g0492(.A1(new_n528), .A2(new_n685), .ZN(new_n693));
  OAI22_X1  g0493(.A1(new_n533), .A2(new_n693), .B1(new_n522), .B2(new_n685), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n660), .A2(new_n662), .A3(new_n685), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n659), .A2(new_n685), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n534), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(G399));
  INV_X1    g0499(.A(new_n213), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n540), .A2(G116), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G1), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n220), .B2(new_n702), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n528), .A2(new_n520), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n532), .B(new_n664), .C1(new_n707), .C2(new_n659), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n573), .B1(new_n669), .B2(KEYINPUT26), .ZN(new_n709));
  INV_X1    g0509(.A(new_n671), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n709), .B1(new_n669), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n686), .B1(new_n708), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT29), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n665), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n660), .A2(new_n662), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n715), .B1(new_n716), .B2(new_n659), .ZN(new_n717));
  OR2_X1    g0517(.A1(new_n673), .A2(new_n676), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n686), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n714), .B1(new_n719), .B2(new_n713), .ZN(new_n720));
  INV_X1    g0520(.A(G330), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n509), .A2(new_n515), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n638), .A2(new_n639), .ZN(new_n723));
  INV_X1    g0523(.A(new_n569), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n606), .A2(new_n722), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT30), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n722), .A2(new_n724), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n728), .A2(KEYINPUT30), .A3(new_n606), .A4(new_n723), .ZN(new_n729));
  AND3_X1   g0529(.A1(new_n599), .A2(new_n360), .A3(new_n569), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(new_n516), .A3(new_n619), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n727), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  AND3_X1   g0532(.A1(new_n732), .A2(KEYINPUT31), .A3(new_n686), .ZN(new_n733));
  AOI21_X1  g0533(.A(KEYINPUT31), .B1(new_n732), .B2(new_n686), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n644), .A2(new_n522), .A3(new_n532), .A4(new_n685), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n721), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n720), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n706), .B1(new_n740), .B2(G1), .ZN(G364));
  INV_X1    g0541(.A(new_n692), .ZN(new_n742));
  INV_X1    g0542(.A(G13), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n209), .B1(new_n744), .B2(G45), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n701), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n742), .B(new_n748), .C1(G330), .C2(new_n690), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n216), .B1(G20), .B2(new_n358), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n210), .A2(G179), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(G190), .A3(G200), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n210), .A2(new_n360), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT93), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G190), .A2(G200), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G311), .ZN(new_n759));
  OAI221_X1 g0559(.A(new_n251), .B1(new_n596), .B2(new_n753), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n529), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n760), .B1(G322), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n752), .A2(new_n529), .A3(G200), .ZN(new_n765));
  INV_X1    g0565(.A(G283), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n752), .A2(new_n757), .ZN(new_n767));
  INV_X1    g0567(.A(G329), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n765), .A2(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT94), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n210), .B1(new_n761), .B2(new_n360), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n507), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n754), .A2(G200), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G190), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OR2_X1    g0575(.A1(KEYINPUT33), .A2(G317), .ZN(new_n776));
  NAND2_X1  g0576(.A1(KEYINPUT33), .A2(G317), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n773), .A2(new_n529), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n772), .B(new_n778), .C1(G326), .C2(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n764), .A2(new_n770), .A3(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n758), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n782), .A2(G77), .B1(new_n763), .B2(G58), .ZN(new_n783));
  INV_X1    g0583(.A(new_n779), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n305), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n753), .A2(new_n436), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n765), .A2(new_n206), .ZN(new_n787));
  NOR4_X1   g0587(.A1(new_n785), .A2(new_n251), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n771), .A2(new_n205), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n789), .B1(G68), .B2(new_n774), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n767), .A2(new_n392), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT32), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n783), .A2(new_n788), .A3(new_n790), .A4(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n751), .B1(new_n781), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G13), .A2(G33), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(G20), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n750), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n700), .A2(new_n615), .ZN(new_n799));
  INV_X1    g0599(.A(new_n262), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n799), .B1(new_n220), .B2(new_n800), .C1(new_n243), .C2(new_n267), .ZN(new_n801));
  INV_X1    g0601(.A(G355), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n213), .A2(new_n259), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n801), .B1(G116), .B2(new_n213), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n748), .B(new_n794), .C1(new_n798), .C2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n797), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n805), .B1(new_n690), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n749), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(G396));
  NAND2_X1  g0609(.A1(new_n386), .A2(KEYINPUT96), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n387), .A2(new_n388), .B1(new_n373), .B2(new_n686), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT97), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT96), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n381), .A2(new_n384), .A3(new_n813), .A4(new_n385), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n810), .A2(new_n811), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n649), .A2(new_n373), .A3(new_n686), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n810), .A2(new_n814), .A3(new_n811), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(KEYINPUT97), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n719), .B(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n747), .B1(new_n823), .B2(new_n738), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n738), .B2(new_n823), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n751), .A2(new_n796), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n747), .B1(new_n826), .B2(G77), .ZN(new_n827));
  INV_X1    g0627(.A(new_n767), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n415), .B1(G132), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(G58), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n771), .A2(new_n830), .B1(new_n765), .B2(new_n321), .ZN(new_n831));
  INV_X1    g0631(.A(new_n753), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n831), .B1(G50), .B2(new_n832), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n774), .A2(G150), .B1(new_n779), .B2(G137), .ZN(new_n834));
  INV_X1    g0634(.A(G143), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n834), .B1(new_n762), .B2(new_n835), .C1(new_n392), .C2(new_n758), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT34), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n829), .B(new_n833), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n251), .B1(new_n767), .B2(new_n759), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n789), .B(new_n840), .C1(new_n782), .C2(G116), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n507), .B2(new_n762), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n765), .A2(new_n436), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(G303), .B2(new_n779), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n774), .A2(KEYINPUT95), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n774), .A2(KEYINPUT95), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n844), .B1(new_n206), .B2(new_n753), .C1(new_n847), .C2(new_n766), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n838), .A2(new_n839), .B1(new_n842), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n827), .B1(new_n849), .B2(new_n750), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n820), .B2(new_n796), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n825), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(G384));
  NOR2_X1   g0653(.A1(new_n744), .A2(new_n209), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT104), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n413), .B1(new_n416), .B2(new_n421), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT77), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n335), .B1(new_n858), .B2(new_n422), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n399), .B1(new_n416), .B2(new_n421), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT101), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n426), .A2(KEYINPUT101), .A3(new_n399), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n862), .A2(new_n411), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n431), .B1(new_n859), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n684), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n457), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n444), .B1(new_n865), .B2(new_n866), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n865), .A2(new_n453), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT37), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT102), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g0673(.A(KEYINPUT102), .B(KEYINPUT37), .C1(new_n869), .C2(new_n870), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n428), .A2(new_n432), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n684), .ZN(new_n876));
  XNOR2_X1  g0676(.A(KEYINPUT103), .B(KEYINPUT37), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n428), .A2(new_n432), .A3(new_n443), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n880), .A2(new_n454), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n873), .A2(new_n874), .A3(new_n882), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n868), .A2(new_n883), .A3(KEYINPUT38), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT38), .B1(new_n868), .B2(new_n883), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n855), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n873), .A2(new_n874), .A3(new_n882), .ZN(new_n888));
  INV_X1    g0688(.A(new_n867), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n655), .B2(new_n455), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n887), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n868), .A2(new_n883), .A3(KEYINPUT38), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n891), .A2(KEYINPUT104), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n886), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n324), .A2(new_n686), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n648), .B(new_n895), .C1(new_n300), .C2(new_n325), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n324), .B(new_n686), .C1(new_n651), .C2(new_n334), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n735), .A2(new_n736), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n898), .A2(new_n899), .A3(new_n820), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT40), .B1(new_n894), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT106), .B1(new_n880), .B2(new_n454), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT106), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n431), .B1(new_n859), .B2(new_n412), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n444), .B(new_n904), .C1(new_n905), .C2(new_n453), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n903), .A2(new_n876), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n877), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n881), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT107), .B1(new_n910), .B2(new_n878), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT107), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n879), .A2(new_n912), .A3(new_n881), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n909), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n455), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n875), .B(new_n684), .C1(new_n915), .C2(new_n448), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n887), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n892), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT40), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n900), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n902), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n459), .B1(new_n736), .B2(new_n735), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n721), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n922), .B2(new_n923), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT108), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n896), .A2(new_n897), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n677), .A2(new_n685), .A3(new_n820), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n810), .A2(new_n814), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n930), .A2(new_n686), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n928), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n894), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT39), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT38), .B1(new_n914), .B2(new_n916), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n935), .B1(new_n884), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n326), .A2(new_n685), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n938), .B(KEYINPUT105), .Z(new_n939));
  NAND3_X1  g0739(.A1(new_n891), .A2(KEYINPUT39), .A3(new_n892), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n915), .A2(new_n866), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n934), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n658), .B1(new_n720), .B2(new_n459), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n943), .B(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n854), .B1(new_n927), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n927), .B2(new_n945), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n624), .A2(new_n625), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT35), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n471), .B(new_n218), .C1(new_n948), .C2(new_n949), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n950), .B1(new_n952), .B2(KEYINPUT98), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(KEYINPUT98), .B2(new_n952), .ZN(new_n954));
  XOR2_X1   g0754(.A(KEYINPUT99), .B(KEYINPUT36), .Z(new_n955));
  XNOR2_X1  g0755(.A(new_n954), .B(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n396), .A2(new_n397), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n220), .A2(new_n957), .A3(new_n308), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT100), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n958), .A2(new_n959), .B1(G68), .B2(new_n201), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n959), .B2(new_n958), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n961), .A2(G1), .A3(new_n743), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n947), .A2(new_n956), .A3(new_n962), .ZN(G367));
  INV_X1    g0763(.A(new_n799), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n798), .B1(new_n213), .B2(new_n366), .C1(new_n964), .C2(new_n236), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n965), .A2(new_n747), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n685), .B1(new_n556), .B2(new_n574), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n674), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n579), .B2(new_n967), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n832), .A2(KEYINPUT46), .A3(G116), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n970), .B1(new_n762), .B2(new_n596), .C1(new_n766), .C2(new_n758), .ZN(new_n971));
  AOI21_X1  g0771(.A(KEYINPUT46), .B1(new_n832), .B2(G116), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n615), .B(new_n972), .C1(G317), .C2(new_n828), .ZN(new_n973));
  INV_X1    g0773(.A(new_n771), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n779), .A2(G311), .B1(new_n974), .B2(G107), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n973), .B(new_n975), .C1(new_n205), .C2(new_n765), .ZN(new_n976));
  INV_X1    g0776(.A(new_n847), .ZN(new_n977));
  AOI211_X1 g0777(.A(new_n971), .B(new_n976), .C1(G294), .C2(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n765), .A2(new_n308), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n259), .B1(new_n784), .B2(new_n835), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n979), .B(new_n980), .C1(G68), .C2(new_n974), .ZN(new_n981));
  INV_X1    g0781(.A(G150), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n981), .B1(new_n982), .B2(new_n762), .C1(new_n201), .C2(new_n758), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT112), .ZN(new_n984));
  INV_X1    g0784(.A(G137), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n753), .A2(new_n830), .B1(new_n767), .B2(new_n985), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n977), .A2(G159), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n984), .B2(new_n986), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n983), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n978), .A2(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(KEYINPUT113), .B(KEYINPUT47), .Z(new_n991));
  XNOR2_X1  g0791(.A(new_n990), .B(new_n991), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n966), .B1(new_n806), .B2(new_n969), .C1(new_n992), .C2(new_n751), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n698), .A2(new_n696), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n634), .B(new_n642), .C1(new_n633), .C2(new_n685), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n667), .A2(new_n686), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n994), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT45), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n994), .A2(new_n998), .ZN(new_n1001));
  XOR2_X1   g0801(.A(KEYINPUT110), .B(KEYINPUT44), .Z(new_n1002));
  XNOR2_X1  g0802(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n695), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1000), .A2(new_n695), .A3(new_n1003), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1004), .A2(KEYINPUT111), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n698), .B1(new_n694), .B2(new_n697), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n692), .B(new_n1011), .Z(new_n1012));
  NOR2_X1   g0812(.A1(new_n1012), .A2(new_n739), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n1009), .B2(new_n1005), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n740), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(KEYINPUT109), .B(KEYINPUT41), .Z(new_n1016));
  XNOR2_X1  g0816(.A(new_n701), .B(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n746), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n534), .A2(new_n697), .A3(new_n997), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1019), .A2(KEYINPUT42), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n642), .B1(new_n522), .B2(new_n995), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1019), .A2(KEYINPUT42), .B1(new_n685), .B2(new_n1021), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n1020), .A2(new_n1022), .B1(KEYINPUT43), .B2(new_n969), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1005), .A2(new_n997), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n993), .B1(new_n1018), .B2(new_n1027), .ZN(G387));
  INV_X1    g0828(.A(new_n1013), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1012), .A2(new_n739), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1029), .A2(new_n701), .A3(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n799), .B1(new_n233), .B2(new_n262), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n703), .B2(new_n803), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n337), .A2(G50), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT50), .ZN(new_n1035));
  AOI21_X1  g0835(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1035), .A2(new_n703), .A3(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1033), .A2(new_n1037), .B1(new_n206), .B2(new_n700), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n798), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n747), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n771), .A2(new_n366), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n775), .A2(new_n337), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1041), .B(new_n1042), .C1(G159), .C2(new_n779), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n782), .A2(G68), .B1(new_n763), .B2(G50), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n308), .A2(new_n753), .B1(new_n765), .B2(new_n205), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n415), .B(new_n1045), .C1(G150), .C2(new_n828), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n615), .B1(G326), .B2(new_n828), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n771), .A2(new_n766), .B1(new_n753), .B2(new_n507), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n782), .A2(G303), .B1(G322), .B2(new_n779), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n763), .A2(G317), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1050), .B(new_n1051), .C1(new_n759), .C2(new_n847), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT48), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1049), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n1053), .B2(new_n1052), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT49), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1048), .B1(new_n471), .B2(new_n765), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  AND2_X1   g0857(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1047), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1040), .B1(new_n1059), .B2(new_n750), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n694), .B2(new_n806), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT114), .Z(new_n1062));
  OAI211_X1 g0862(.A(new_n1031), .B(new_n1062), .C1(new_n745), .C2(new_n1012), .ZN(G393));
  INV_X1    g0863(.A(new_n1008), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n701), .B1(new_n1064), .B2(new_n1013), .C1(new_n1010), .C2(new_n1014), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n998), .A2(new_n797), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n798), .B1(new_n205), .B2(new_n213), .C1(new_n964), .C2(new_n240), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n747), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n763), .A2(G311), .B1(G317), .B2(new_n779), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1069), .B(new_n1070), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n259), .B(new_n787), .C1(G322), .C2(new_n828), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n974), .A2(G116), .B1(new_n832), .B2(G283), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1074), .B1(new_n507), .B2(new_n758), .C1(new_n596), .C2(new_n847), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n762), .A2(new_n392), .B1(new_n982), .B2(new_n784), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT51), .Z(new_n1077));
  INV_X1    g0877(.A(new_n201), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n977), .A2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n753), .A2(new_n321), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n843), .B(new_n1080), .C1(G77), .C2(new_n974), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n782), .A2(new_n338), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n415), .B1(G143), .B2(new_n828), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n1071), .A2(new_n1075), .B1(new_n1077), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1068), .B1(new_n1085), .B2(new_n750), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1064), .A2(new_n746), .B1(new_n1066), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1065), .A2(new_n1087), .ZN(G390));
  NAND3_X1  g0888(.A1(new_n898), .A2(new_n737), .A3(new_n820), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n929), .A2(new_n932), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n898), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n938), .B(KEYINPUT105), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1092), .A2(new_n1093), .B1(new_n937), .B2(new_n940), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n712), .A2(new_n820), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n898), .B1(new_n1095), .B2(new_n931), .ZN(new_n1096));
  AND3_X1   g0896(.A1(new_n1096), .A2(new_n919), .A3(new_n1093), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1090), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1096), .A2(new_n919), .A3(new_n1093), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n937), .A2(new_n940), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n933), .A2(new_n939), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1089), .B(new_n1099), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1098), .A2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1103), .A2(new_n745), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n747), .B1(new_n826), .B2(new_n338), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1100), .A2(new_n796), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(KEYINPUT54), .B(G143), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT118), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n782), .A2(new_n1108), .B1(new_n763), .B2(G132), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n779), .A2(G128), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n974), .A2(G159), .B1(new_n828), .B2(G125), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n259), .B1(new_n201), .B2(new_n765), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT119), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n753), .A2(new_n982), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT53), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1114), .B(new_n1116), .C1(new_n985), .C2(new_n847), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n259), .B(new_n786), .C1(G294), .C2(new_n828), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1118), .B1(new_n205), .B2(new_n758), .C1(new_n471), .C2(new_n762), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n765), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n974), .A2(G77), .B1(new_n1120), .B2(G68), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1121), .B1(new_n766), .B2(new_n784), .C1(new_n847), .C2(new_n206), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1112), .A2(new_n1117), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1105), .B(new_n1106), .C1(new_n750), .C2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1104), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT116), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n820), .B1(new_n737), .B2(new_n1126), .ZN(new_n1127));
  AOI211_X1 g0927(.A(KEYINPUT116), .B(new_n721), .C1(new_n735), .C2(new_n736), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n928), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n931), .B1(new_n712), .B2(new_n820), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1089), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n899), .A2(new_n820), .A3(G330), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n928), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n1089), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1129), .A2(new_n1131), .B1(new_n1134), .B2(new_n1091), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n391), .A2(new_n458), .A3(new_n737), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n658), .B(new_n1136), .C1(new_n720), .C2(new_n459), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n702), .B1(new_n1103), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1098), .A2(new_n1102), .A3(new_n1138), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1140), .A2(KEYINPUT117), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(KEYINPUT117), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1125), .B1(new_n1142), .B2(new_n1143), .ZN(G378));
  INV_X1    g0944(.A(new_n1137), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1141), .A2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n866), .A2(new_n345), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n364), .B(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1148), .B(new_n1149), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(new_n884), .A2(new_n885), .A3(new_n855), .ZN(new_n1151));
  AOI21_X1  g0951(.A(KEYINPUT104), .B1(new_n891), .B2(new_n892), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n901), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n920), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n721), .B1(new_n921), .B2(new_n919), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1150), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n900), .B1(new_n886), .B2(new_n893), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1155), .B(new_n1150), .C1(new_n1157), .C2(KEYINPUT40), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n943), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1150), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1155), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1161), .B1(new_n902), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n943), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1163), .A2(new_n1164), .A3(new_n1158), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1146), .A2(new_n1160), .A3(KEYINPUT57), .A4(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n943), .A2(KEYINPUT121), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1163), .A2(KEYINPUT121), .A3(new_n943), .A4(new_n1158), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n1168), .A2(new_n1169), .B1(new_n1145), .B2(new_n1141), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1166), .B(new_n701), .C1(new_n1170), .C2(KEYINPUT57), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n745), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1150), .A2(new_n795), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n747), .B1(new_n826), .B2(new_n1078), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n206), .A2(new_n762), .B1(new_n758), .B2(new_n366), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n774), .A2(G97), .B1(new_n1120), .B2(G58), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n471), .B2(new_n784), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n415), .B(new_n263), .C1(new_n766), .C2(new_n767), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n771), .A2(new_n321), .B1(new_n753), .B2(new_n308), .ZN(new_n1179));
  NOR4_X1   g0979(.A1(new_n1175), .A2(new_n1177), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n263), .B1(new_n419), .B2(new_n256), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1180), .A2(KEYINPUT58), .B1(new_n305), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1108), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1183), .A2(new_n753), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT120), .Z(new_n1185));
  NAND2_X1  g0985(.A1(new_n974), .A2(G150), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n774), .A2(G132), .B1(new_n779), .B2(G125), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n782), .A2(G137), .B1(new_n763), .B2(G128), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(KEYINPUT59), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1120), .A2(G159), .ZN(new_n1191));
  AOI211_X1 g0991(.A(G33), .B(G41), .C1(new_n828), .C2(G124), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1189), .A2(KEYINPUT59), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1182), .B1(KEYINPUT58), .B2(new_n1180), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1174), .B1(new_n1195), .B2(new_n750), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1172), .B1(new_n1173), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT122), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n1171), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1198), .B1(new_n1171), .B2(new_n1197), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1199), .A2(new_n1200), .ZN(G375));
  NAND2_X1  g1001(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1139), .A2(new_n1017), .A3(new_n1202), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT123), .Z(new_n1204));
  INV_X1    g1004(.A(new_n1135), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n928), .A2(new_n795), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n747), .B1(new_n826), .B2(G68), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n259), .B(new_n979), .C1(G303), .C2(new_n828), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n206), .B2(new_n758), .C1(new_n766), .C2(new_n762), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1041), .B1(G294), .B2(new_n779), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1210), .B1(new_n205), .B2(new_n753), .C1(new_n847), .C2(new_n471), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n415), .B1(G128), .B2(new_n828), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1212), .B1(new_n762), .B2(new_n985), .C1(new_n982), .C2(new_n758), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n974), .A2(G50), .B1(new_n1120), .B2(G58), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n779), .A2(G132), .B1(new_n832), .B2(G159), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1214), .B(new_n1215), .C1(new_n847), .C2(new_n1183), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n1209), .A2(new_n1211), .B1(new_n1213), .B2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1207), .B1(new_n1217), .B2(new_n750), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1205), .A2(new_n746), .B1(new_n1206), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1204), .A2(new_n1219), .ZN(G381));
  OR4_X1    g1020(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n1221), .A2(G387), .A3(G381), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1125), .A2(new_n1223), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(G375), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1222), .A2(new_n1225), .ZN(G407));
  INV_X1    g1026(.A(G343), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1225), .B1(new_n1222), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(G213), .ZN(G409));
  NAND2_X1  g1029(.A1(new_n1227), .A2(G213), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1171), .A2(new_n1197), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n1232), .A2(G378), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1160), .A2(new_n746), .A3(new_n1165), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1173), .A2(new_n1196), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT124), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n1017), .B2(new_n1170), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1234), .A2(KEYINPUT124), .A3(new_n1235), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1224), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1230), .B1(new_n1233), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1139), .A2(KEYINPUT60), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1241), .A2(new_n1202), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n701), .B1(new_n1241), .B2(new_n1202), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1219), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1244), .A2(new_n852), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n852), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1227), .A2(G213), .A3(G2897), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1247), .B(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(KEYINPUT61), .B1(new_n1240), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1239), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1232), .A2(G378), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1251), .A2(new_n1252), .B1(G213), .B2(new_n1227), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1247), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1253), .A2(KEYINPUT63), .A3(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(G387), .A2(new_n1065), .A3(new_n1087), .ZN(new_n1256));
  OAI211_X1 g1056(.A(G390), .B(new_n993), .C1(new_n1018), .C2(new_n1027), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(G393), .B(new_n808), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1258), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1230), .B(new_n1254), .C1(new_n1233), .C2(new_n1239), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT63), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1250), .A2(new_n1255), .A3(new_n1261), .A4(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT125), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(KEYINPUT62), .ZN(new_n1267));
  OR2_X1    g1067(.A1(new_n1266), .A2(KEYINPUT62), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1253), .A2(new_n1267), .A3(new_n1268), .A4(new_n1254), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1262), .A2(new_n1266), .A3(KEYINPUT62), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1269), .A2(new_n1270), .A3(new_n1250), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1265), .B1(new_n1271), .B2(new_n1261), .ZN(G405));
  INV_X1    g1072(.A(KEYINPUT126), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1224), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1273), .B1(G375), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1231), .A2(KEYINPUT122), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1171), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1276), .A2(new_n1273), .A3(new_n1277), .A4(new_n1274), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1252), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1247), .B1(new_n1275), .B2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1276), .A2(new_n1277), .A3(new_n1274), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(KEYINPUT126), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1282), .A2(new_n1252), .A3(new_n1254), .A4(new_n1278), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1280), .A2(new_n1261), .A3(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(KEYINPUT127), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT127), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1280), .A2(new_n1261), .A3(new_n1286), .A4(new_n1283), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1261), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1285), .A2(new_n1287), .A3(new_n1290), .ZN(G402));
endmodule


