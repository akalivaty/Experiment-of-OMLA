//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 0 1 0 0 1 1 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1282, new_n1283, new_n1284, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  INV_X1    g0004(.A(KEYINPUT64), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  NOR2_X1   g0007(.A1(G58), .A2(G68), .ZN(new_n208));
  NAND3_X1  g0008(.A1(new_n208), .A2(KEYINPUT64), .A3(new_n201), .ZN(new_n209));
  AND3_X1   g0009(.A1(new_n206), .A2(new_n207), .A3(new_n209), .ZN(G353));
  OAI21_X1  g0010(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  OR3_X1    g0012(.A1(new_n212), .A2(KEYINPUT65), .A3(G13), .ZN(new_n213));
  OAI21_X1  g0013(.A(KEYINPUT65), .B1(new_n212), .B2(G13), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT0), .ZN(new_n217));
  AND2_X1   g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G20), .ZN(new_n219));
  OAI21_X1  g0019(.A(G50), .B1(G58), .B2(G68), .ZN(new_n220));
  OAI22_X1  g0020(.A1(new_n216), .A2(new_n217), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(new_n217), .B2(new_n216), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT66), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT67), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n212), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT1), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n223), .A2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G226), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XNOR2_X1  g0041(.A(G68), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n201), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n202), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT69), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n245), .B(new_n249), .ZN(G351));
  NAND2_X1  g0050(.A1(G1), .A2(G13), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n251), .B1(G33), .B2(G41), .ZN(new_n252));
  INV_X1    g0052(.A(G41), .ZN(new_n253));
  INV_X1    g0053(.A(G45), .ZN(new_n254));
  AOI21_X1  g0054(.A(G1), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT71), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT71), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G41), .A2(G45), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n257), .B1(new_n258), .B2(G1), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n252), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  XOR2_X1   g0060(.A(KEYINPUT70), .B(G226), .Z(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G274), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n263), .B1(new_n218), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n255), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G77), .ZN(new_n271));
  AND2_X1   g0071(.A1(KEYINPUT72), .A2(G1698), .ZN(new_n272));
  NOR2_X1   g0072(.A1(KEYINPUT72), .A2(G1698), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n274), .A2(G222), .B1(G223), .B2(G1698), .ZN(new_n275));
  OAI211_X1 g0075(.A(KEYINPUT73), .B(new_n271), .C1(new_n275), .C2(new_n270), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT73), .ZN(new_n277));
  OR2_X1    g0077(.A1(KEYINPUT72), .A2(G1698), .ZN(new_n278));
  NAND2_X1  g0078(.A1(KEYINPUT72), .A2(G1698), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n278), .A2(G222), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G223), .A2(G1698), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n270), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT3), .ZN(new_n283));
  INV_X1    g0083(.A(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(new_n207), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n277), .B1(new_n282), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n276), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n267), .B1(new_n290), .B2(new_n252), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT76), .ZN(new_n292));
  AND3_X1   g0092(.A1(new_n291), .A2(new_n292), .A3(G190), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n292), .B1(new_n291), .B2(G190), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n251), .ZN(new_n297));
  INV_X1    g0097(.A(G20), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n298), .B1(new_n206), .B2(new_n209), .ZN(new_n299));
  XNOR2_X1  g0099(.A(KEYINPUT8), .B(G58), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(G33), .ZN(new_n301));
  INV_X1    g0101(.A(G150), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n298), .A2(new_n284), .ZN(new_n303));
  OAI22_X1  g0103(.A1(new_n300), .A2(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n297), .B1(new_n299), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT75), .ZN(new_n306));
  INV_X1    g0106(.A(G13), .ZN(new_n307));
  NOR3_X1   g0107(.A1(new_n307), .A2(new_n298), .A3(G1), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(new_n297), .ZN(new_n309));
  INV_X1    g0109(.A(G1), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n201), .B1(new_n310), .B2(G20), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n309), .A2(new_n311), .B1(new_n201), .B2(new_n308), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n305), .A2(new_n306), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n306), .B1(new_n305), .B2(new_n312), .ZN(new_n315));
  NOR3_X1   g0115(.A1(new_n314), .A2(KEYINPUT9), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT9), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n305), .A2(new_n312), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT75), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n317), .B1(new_n319), .B2(new_n313), .ZN(new_n320));
  INV_X1    g0120(.A(G200), .ZN(new_n321));
  OAI22_X1  g0121(.A1(new_n316), .A2(new_n320), .B1(new_n321), .B2(new_n291), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT10), .B1(new_n295), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(KEYINPUT9), .B1(new_n314), .B2(new_n315), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n319), .A2(new_n317), .A3(new_n313), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n290), .A2(new_n252), .ZN(new_n326));
  INV_X1    g0126(.A(new_n267), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n324), .A2(new_n325), .B1(new_n328), .B2(G200), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT10), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n329), .B(new_n330), .C1(new_n293), .C2(new_n294), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n323), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G169), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G179), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n291), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n318), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n298), .A2(G33), .A3(G77), .ZN(new_n339));
  OAI221_X1 g0139(.A(new_n339), .B1(new_n298), .B2(G68), .C1(new_n303), .C2(new_n201), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n297), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT11), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n340), .A2(KEYINPUT11), .A3(new_n297), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n307), .A2(G1), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT12), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n298), .A2(G68), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n345), .A2(G20), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n348), .A2(new_n349), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n343), .A2(new_n344), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n297), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n353), .A2(new_n350), .A3(KEYINPUT74), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT74), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(new_n308), .B2(new_n297), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n310), .A2(G20), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n354), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n203), .B1(new_n358), .B2(KEYINPUT12), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n352), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n360), .B(KEYINPUT79), .ZN(new_n361));
  INV_X1    g0161(.A(new_n266), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n362), .B1(new_n260), .B2(G238), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n287), .A2(G232), .A3(G1698), .ZN(new_n364));
  NAND2_X1  g0164(.A1(G33), .A2(G97), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n287), .A2(new_n274), .A3(G226), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT77), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n287), .A2(new_n274), .A3(KEYINPUT77), .A4(G226), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n366), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n218), .A2(new_n264), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n363), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT13), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT13), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n375), .B(new_n363), .C1(new_n371), .C2(new_n372), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT14), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n378), .A3(G169), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n373), .A2(KEYINPUT78), .A3(KEYINPUT13), .ZN(new_n380));
  NAND2_X1  g0180(.A1(KEYINPUT78), .A2(KEYINPUT13), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n363), .B(new_n381), .C1(new_n371), .C2(new_n372), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n380), .A2(new_n382), .A3(G179), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n378), .B1(new_n377), .B2(G169), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n361), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n380), .A2(new_n382), .A3(G190), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n321), .B1(new_n374), .B2(new_n376), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n387), .A2(new_n361), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  OR2_X1    g0191(.A1(new_n358), .A2(new_n207), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G20), .A2(G77), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT15), .B(G87), .ZN(new_n394));
  OAI221_X1 g0194(.A(new_n393), .B1(new_n300), .B2(new_n303), .C1(new_n301), .C2(new_n394), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n395), .A2(new_n297), .B1(new_n207), .B2(new_n308), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G238), .A2(G1698), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n278), .A2(new_n279), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n287), .B(new_n399), .C1(new_n400), .C2(new_n236), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n401), .B(new_n252), .C1(G107), .C2(new_n287), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n260), .A2(G244), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(new_n266), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(G200), .ZN(new_n405));
  INV_X1    g0205(.A(G190), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n398), .B(new_n405), .C1(new_n406), .C2(new_n404), .ZN(new_n407));
  OR2_X1    g0207(.A1(new_n404), .A2(G179), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n404), .A2(new_n333), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(new_n397), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  NOR3_X1   g0211(.A1(new_n338), .A2(new_n391), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n309), .ZN(new_n413));
  INV_X1    g0213(.A(new_n300), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n357), .ZN(new_n415));
  OAI22_X1  g0215(.A1(new_n413), .A2(new_n415), .B1(new_n350), .B2(new_n414), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT82), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n202), .A2(new_n203), .ZN(new_n418));
  OAI21_X1  g0218(.A(G20), .B1(new_n418), .B2(new_n208), .ZN(new_n419));
  NOR2_X1   g0219(.A1(G20), .A2(G33), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(G159), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT16), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT80), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n268), .B2(new_n269), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n285), .A2(KEYINPUT80), .A3(new_n286), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n426), .A2(new_n427), .A3(new_n298), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT7), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n268), .A2(new_n269), .A3(G20), .ZN(new_n431));
  XOR2_X1   g0231(.A(KEYINPUT81), .B(KEYINPUT7), .Z(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n424), .B1(new_n434), .B2(G68), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n285), .A2(KEYINPUT7), .A3(new_n298), .A4(new_n286), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n431), .B2(new_n432), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n422), .B1(new_n437), .B2(G68), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n297), .B1(new_n438), .B2(KEYINPUT16), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n417), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT16), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n422), .A2(new_n441), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n428), .A2(new_n429), .B1(new_n431), .B2(new_n432), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n442), .B1(new_n443), .B2(new_n203), .ZN(new_n444));
  XNOR2_X1  g0244(.A(KEYINPUT81), .B(KEYINPUT7), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n445), .B1(new_n287), .B2(G20), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n203), .B1(new_n446), .B2(new_n436), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n441), .B1(new_n447), .B2(new_n422), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n444), .A2(KEYINPUT82), .A3(new_n448), .A4(new_n297), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n416), .B1(new_n440), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G1698), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n451), .B1(new_n285), .B2(new_n286), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G226), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT83), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT83), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n452), .A2(new_n455), .A3(G226), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n287), .A2(G223), .ZN(new_n458));
  INV_X1    g0258(.A(G87), .ZN(new_n459));
  OAI22_X1  g0259(.A1(new_n458), .A2(new_n400), .B1(new_n284), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n372), .B1(new_n457), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n362), .B1(new_n260), .B2(G232), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n321), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n460), .B1(new_n456), .B2(new_n454), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n463), .B1(new_n466), .B2(new_n372), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n465), .B1(G190), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g0268(.A(KEYINPUT85), .B(KEYINPUT17), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n450), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n450), .A2(new_n468), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT17), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT85), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n470), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n416), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n437), .A2(G68), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n423), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n353), .B1(new_n477), .B2(new_n441), .ZN(new_n478));
  AOI21_X1  g0278(.A(KEYINPUT82), .B1(new_n478), .B2(new_n444), .ZN(new_n479));
  INV_X1    g0279(.A(new_n449), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n475), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(G169), .B1(new_n462), .B2(new_n464), .ZN(new_n482));
  OAI211_X1 g0282(.A(G179), .B(new_n463), .C1(new_n466), .C2(new_n372), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n481), .A2(KEYINPUT18), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT18), .B1(new_n481), .B2(new_n484), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT84), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n482), .A2(new_n483), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT18), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n450), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n490), .B1(new_n450), .B2(new_n489), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT84), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n474), .B1(new_n488), .B2(new_n493), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n412), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT5), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(G41), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n254), .A2(G1), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n496), .A2(G41), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n265), .A2(new_n498), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n310), .B(G45), .C1(new_n253), .C2(KEYINPUT5), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n372), .B(G264), .C1(new_n502), .C2(new_n497), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(G257), .B(G1698), .C1(new_n268), .C2(new_n269), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G33), .A2(G294), .ZN(new_n507));
  OAI21_X1  g0307(.A(G250), .B1(new_n268), .B2(new_n269), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n506), .B(new_n507), .C1(new_n508), .C2(new_n400), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n252), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n505), .A2(new_n510), .A3(G179), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n506), .A2(new_n507), .ZN(new_n512));
  INV_X1    g0312(.A(G250), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n513), .B1(new_n285), .B2(new_n286), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n274), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n372), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n516), .A2(new_n504), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n511), .B1(new_n517), .B2(new_n333), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT23), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(new_n298), .B2(G107), .ZN(new_n520));
  INV_X1    g0320(.A(G107), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n521), .A2(KEYINPUT23), .A3(G20), .ZN(new_n522));
  INV_X1    g0322(.A(G116), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n284), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n520), .A2(new_n522), .B1(new_n524), .B2(new_n298), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n298), .B(G87), .C1(new_n268), .C2(new_n269), .ZN(new_n526));
  AND2_X1   g0326(.A1(new_n526), .A2(KEYINPUT22), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n526), .A2(KEYINPUT22), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(KEYINPUT24), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT24), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n531), .B(new_n525), .C1(new_n527), .C2(new_n528), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n353), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n309), .B1(G1), .B2(new_n284), .ZN(new_n534));
  AOI21_X1  g0334(.A(KEYINPUT25), .B1(new_n308), .B2(new_n521), .ZN(new_n535));
  AND3_X1   g0335(.A1(new_n308), .A2(KEYINPUT25), .A3(new_n521), .ZN(new_n536));
  OAI22_X1  g0336(.A1(new_n534), .A2(new_n521), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n518), .B1(new_n533), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n530), .A2(new_n532), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n537), .B1(new_n539), .B2(new_n297), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n505), .A2(new_n510), .A3(new_n406), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT91), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n505), .A2(new_n510), .A3(KEYINPUT91), .A4(new_n406), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n321), .B1(new_n516), .B2(new_n504), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n540), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT4), .ZN(new_n548));
  OAI21_X1  g0348(.A(G244), .B1(new_n268), .B2(new_n269), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n548), .B1(new_n549), .B2(new_n400), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n287), .A2(new_n274), .A3(KEYINPUT4), .A4(G244), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G33), .A2(G283), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n514), .A2(G1698), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n550), .A2(new_n551), .A3(new_n552), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n252), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n372), .B(G257), .C1(new_n502), .C2(new_n497), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n501), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(G169), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(KEYINPUT6), .A2(G97), .ZN(new_n561));
  OR3_X1    g0361(.A1(new_n561), .A2(KEYINPUT87), .A3(G107), .ZN(new_n562));
  OAI21_X1  g0362(.A(KEYINPUT87), .B1(new_n561), .B2(G107), .ZN(new_n563));
  INV_X1    g0363(.A(G97), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n564), .A2(new_n521), .ZN(new_n565));
  NOR2_X1   g0365(.A1(G97), .A2(G107), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n562), .B(new_n563), .C1(new_n567), .C2(KEYINPUT6), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G20), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n437), .A2(G107), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n420), .A2(G77), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT86), .ZN(new_n572));
  XNOR2_X1  g0372(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n569), .A2(new_n570), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n297), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n350), .A2(G97), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n534), .B2(new_n564), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  AOI211_X1 g0381(.A(G179), .B(new_n557), .C1(new_n554), .C2(new_n252), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n560), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n579), .B1(new_n575), .B2(new_n297), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n557), .B1(new_n554), .B2(new_n252), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G190), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n585), .B(new_n587), .C1(new_n321), .C2(new_n586), .ZN(new_n588));
  AND4_X1   g0388(.A1(new_n538), .A2(new_n547), .A3(new_n584), .A4(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n523), .B1(new_n310), .B2(G33), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n354), .A2(new_n356), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n345), .A2(G20), .A3(new_n523), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n552), .B(new_n298), .C1(G33), .C2(new_n564), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT90), .ZN(new_n594));
  AOI21_X1  g0394(.A(G20), .B1(new_n284), .B2(G97), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT90), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n596), .A3(new_n552), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n296), .A2(new_n251), .B1(G20), .B2(new_n523), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(KEYINPUT20), .A3(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(KEYINPUT20), .B1(new_n598), .B2(new_n599), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n591), .B(new_n592), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n372), .B(G270), .C1(new_n502), .C2(new_n497), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n501), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT89), .ZN(new_n606));
  INV_X1    g0406(.A(G257), .ZN(new_n607));
  NOR3_X1   g0407(.A1(new_n272), .A2(new_n273), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(G264), .A2(G1698), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n268), .B2(new_n269), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n252), .B1(new_n287), .B2(G303), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n606), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n287), .B(new_n609), .C1(new_n400), .C2(new_n607), .ZN(new_n614));
  INV_X1    g0414(.A(G303), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n372), .B1(new_n270), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(new_n616), .A3(KEYINPUT89), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n605), .B1(new_n613), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n603), .A2(G179), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(G190), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n591), .A2(new_n592), .ZN(new_n621));
  INV_X1    g0421(.A(new_n602), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n621), .B1(new_n622), .B2(new_n600), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n620), .B(new_n623), .C1(new_n321), .C2(new_n618), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n613), .A2(new_n617), .ZN(new_n625));
  INV_X1    g0425(.A(new_n605), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n333), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT21), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n627), .A2(new_n603), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n628), .B1(new_n627), .B2(new_n603), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n619), .B(new_n624), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n459), .A2(new_n564), .A3(new_n521), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n365), .A2(new_n298), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(new_n634), .A3(KEYINPUT19), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n298), .B(G68), .C1(new_n268), .C2(new_n269), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT19), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(new_n301), .B2(new_n564), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n635), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n639), .A2(new_n297), .B1(new_n308), .B2(new_n394), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n309), .B(G87), .C1(G1), .C2(new_n284), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n278), .A2(G238), .A3(new_n279), .ZN(new_n643));
  NAND2_X1  g0443(.A1(G244), .A2(G1698), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n270), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(KEYINPUT88), .B1(new_n645), .B2(new_n524), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT88), .ZN(new_n647));
  INV_X1    g0447(.A(new_n524), .ZN(new_n648));
  INV_X1    g0448(.A(new_n644), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(new_n274), .B2(G238), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n647), .B(new_n648), .C1(new_n650), .C2(new_n270), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n646), .A2(new_n651), .A3(new_n252), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n499), .A2(new_n263), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n513), .B1(new_n254), .B2(G1), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(new_n372), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n652), .A2(G190), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n655), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n648), .B1(new_n650), .B2(new_n270), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n372), .B1(new_n658), .B2(KEYINPUT88), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n657), .B1(new_n659), .B2(new_n651), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n642), .B(new_n656), .C1(new_n660), .C2(new_n321), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n652), .A2(new_n335), .A3(new_n655), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n640), .B1(new_n394), .B2(new_n534), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n662), .B(new_n663), .C1(new_n660), .C2(G169), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  AND4_X1   g0465(.A1(new_n495), .A2(new_n589), .A3(new_n632), .A4(new_n665), .ZN(G372));
  INV_X1    g0466(.A(new_n664), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n640), .A2(KEYINPUT92), .A3(new_n641), .ZN(new_n668));
  AOI21_X1  g0468(.A(KEYINPUT92), .B1(new_n640), .B2(new_n641), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n652), .A2(new_n655), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(G200), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n670), .A2(new_n672), .A3(new_n656), .ZN(new_n673));
  AND4_X1   g0473(.A1(new_n547), .A2(new_n673), .A3(new_n584), .A4(new_n588), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n538), .B(new_n619), .C1(new_n629), .C2(new_n630), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n667), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n585), .A2(new_n559), .A3(new_n582), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n678), .A2(new_n661), .A3(new_n664), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(KEYINPUT26), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT26), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n673), .A2(new_n678), .A3(new_n664), .A4(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n495), .B1(new_n677), .B2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n337), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n485), .A2(new_n492), .ZN(new_n686));
  INV_X1    g0486(.A(new_n410), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n377), .A2(G169), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(KEYINPUT14), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n689), .A2(new_n383), .A3(new_n379), .ZN(new_n690));
  AOI22_X1  g0490(.A1(new_n390), .A2(new_n687), .B1(new_n690), .B2(new_n361), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n686), .B1(new_n691), .B2(new_n474), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n685), .B1(new_n692), .B2(new_n332), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n684), .A2(new_n693), .ZN(G369));
  OR2_X1    g0494(.A1(new_n629), .A2(new_n630), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n619), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n346), .A2(KEYINPUT27), .A3(G20), .ZN(new_n697));
  INV_X1    g0497(.A(G213), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT27), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n699), .B1(new_n345), .B2(new_n298), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n697), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(G343), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n623), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n696), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n631), .B2(new_n703), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G330), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n547), .A2(new_n538), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n540), .B2(new_n702), .ZN(new_n709));
  INV_X1    g0509(.A(new_n538), .ZN(new_n710));
  INV_X1    g0510(.A(new_n702), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n707), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n711), .B1(new_n695), .B2(new_n619), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n715), .A2(new_n708), .B1(new_n710), .B2(new_n702), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n714), .A2(new_n716), .ZN(G399));
  INV_X1    g0517(.A(new_n215), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G41), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n633), .A2(G116), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n719), .A2(new_n310), .A3(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n220), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(new_n719), .ZN(new_n723));
  XOR2_X1   g0523(.A(new_n723), .B(KEYINPUT28), .Z(new_n724));
  NAND2_X1  g0524(.A1(new_n679), .A2(new_n681), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n673), .A2(new_n678), .A3(new_n664), .A4(KEYINPUT26), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI211_X1 g0527(.A(KEYINPUT95), .B(new_n711), .C1(new_n676), .C2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT95), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n321), .B1(new_n555), .B2(new_n558), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n573), .B1(G107), .B2(new_n437), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n353), .B1(new_n731), .B2(new_n569), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n730), .A2(new_n732), .A3(new_n579), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n559), .A2(new_n582), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n733), .A2(new_n587), .B1(new_n734), .B2(new_n581), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n675), .A2(new_n735), .A3(new_n547), .A4(new_n673), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n727), .A2(new_n664), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n729), .B1(new_n737), .B2(new_n702), .ZN(new_n738));
  OAI21_X1  g0538(.A(KEYINPUT29), .B1(new_n728), .B2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT96), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI211_X1 g0541(.A(KEYINPUT96), .B(KEYINPUT29), .C1(new_n728), .C2(new_n738), .ZN(new_n742));
  INV_X1    g0542(.A(new_n683), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n711), .B1(new_n743), .B2(new_n676), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n744), .A2(KEYINPUT29), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n741), .A2(new_n742), .A3(new_n745), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n589), .A2(new_n632), .A3(new_n665), .A4(new_n702), .ZN(new_n747));
  INV_X1    g0547(.A(new_n586), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n625), .A2(new_n626), .ZN(new_n749));
  AOI21_X1  g0549(.A(G179), .B1(new_n505), .B2(new_n510), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n671), .A2(new_n748), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT94), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT30), .ZN(new_n754));
  INV_X1    g0554(.A(new_n604), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n755), .B1(new_n613), .B2(new_n617), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n517), .A2(new_n586), .A3(new_n756), .A4(G179), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n754), .B1(new_n757), .B2(new_n671), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n611), .A2(new_n612), .A3(new_n606), .ZN(new_n759));
  AOI21_X1  g0559(.A(KEYINPUT89), .B1(new_n614), .B2(new_n616), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n604), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n511), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n762), .A2(KEYINPUT30), .A3(new_n660), .A4(new_n586), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n335), .B1(new_n516), .B2(new_n504), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n618), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n765), .A2(KEYINPUT94), .A3(new_n748), .A4(new_n671), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n753), .A2(new_n758), .A3(new_n763), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n711), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT31), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n758), .A2(new_n763), .A3(new_n751), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n702), .A2(new_n769), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n771), .A2(KEYINPUT93), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT93), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n747), .A2(new_n770), .A3(new_n773), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G330), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n746), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n724), .B1(new_n779), .B2(G1), .ZN(G364));
  NOR2_X1   g0580(.A1(new_n307), .A2(G20), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n310), .B1(new_n781), .B2(G45), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n719), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n707), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(G330), .B2(new_n705), .ZN(new_n786));
  XOR2_X1   g0586(.A(new_n784), .B(KEYINPUT97), .Z(new_n787));
  NOR2_X1   g0587(.A1(new_n298), .A2(new_n335), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n788), .A2(G190), .A3(new_n321), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(G200), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(G190), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n287), .B1(new_n202), .B2(new_n789), .C1(new_n792), .C2(new_n203), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n406), .A2(G179), .A3(G200), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n298), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n564), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n298), .A2(G179), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n797), .A2(G190), .A3(G200), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n459), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n790), .A2(new_n406), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n797), .A2(new_n406), .A3(G200), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n800), .B1(new_n201), .B2(new_n802), .C1(new_n521), .C2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(G190), .A2(G200), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n788), .A2(new_n805), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n806), .A2(KEYINPUT98), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(KEYINPUT98), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n793), .B(new_n804), .C1(G77), .C2(new_n810), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n797), .A2(new_n805), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n812), .A2(KEYINPUT99), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(KEYINPUT99), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G159), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT32), .ZN(new_n818));
  INV_X1    g0618(.A(new_n789), .ZN(new_n819));
  INV_X1    g0619(.A(new_n806), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n819), .A2(G322), .B1(new_n820), .B2(G311), .ZN(new_n821));
  INV_X1    g0621(.A(G294), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n822), .B2(new_n795), .ZN(new_n823));
  INV_X1    g0623(.A(G317), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(KEYINPUT33), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n824), .A2(KEYINPUT33), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n791), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(G283), .ZN(new_n828));
  INV_X1    g0628(.A(G326), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n827), .B1(new_n828), .B2(new_n803), .C1(new_n829), .C2(new_n802), .ZN(new_n830));
  INV_X1    g0630(.A(new_n815), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n823), .B(new_n830), .C1(G329), .C2(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n270), .B1(new_n798), .B2(new_n615), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT100), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n811), .A2(new_n818), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n251), .B1(G20), .B2(new_n333), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n787), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(G13), .A2(G33), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(G20), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n841), .A2(new_n836), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n426), .A2(new_n427), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n718), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(new_n254), .B2(new_n722), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n245), .B2(new_n254), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n718), .A2(new_n270), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n848), .A2(G355), .B1(new_n523), .B2(new_n718), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n838), .B1(new_n842), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n841), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n851), .B1(new_n705), .B2(new_n852), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n786), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(G396));
  OAI21_X1  g0655(.A(new_n407), .B1(new_n398), .B2(new_n702), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n410), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n687), .A2(new_n702), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n744), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n744), .A2(new_n860), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n784), .B1(new_n863), .B2(new_n778), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n778), .B2(new_n863), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n836), .A2(new_n839), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT101), .ZN(new_n867));
  AOI22_X1  g0667(.A1(G150), .A2(new_n791), .B1(new_n819), .B2(G143), .ZN(new_n868));
  INV_X1    g0668(.A(G137), .ZN(new_n869));
  OAI221_X1 g0669(.A(new_n868), .B1(new_n869), .B2(new_n802), .C1(new_n809), .C2(new_n816), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT34), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n843), .B1(new_n201), .B2(new_n798), .ZN(new_n872));
  OAI22_X1  g0672(.A1(new_n795), .A2(new_n202), .B1(new_n803), .B2(new_n203), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n872), .B(new_n873), .C1(new_n831), .C2(G132), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n803), .A2(new_n459), .ZN(new_n875));
  OAI22_X1  g0675(.A1(new_n792), .A2(new_n828), .B1(new_n802), .B2(new_n615), .ZN(new_n876));
  INV_X1    g0676(.A(new_n798), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n875), .B(new_n876), .C1(G107), .C2(new_n877), .ZN(new_n878));
  OAI221_X1 g0678(.A(new_n270), .B1(new_n789), .B2(new_n822), .C1(new_n564), .C2(new_n795), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n809), .A2(new_n523), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n879), .B(new_n880), .C1(G311), .C2(new_n831), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n871), .A2(new_n874), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n787), .B1(G77), .B2(new_n867), .C1(new_n882), .C2(new_n837), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n883), .A2(KEYINPUT102), .B1(new_n839), .B2(new_n859), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(KEYINPUT102), .B2(new_n883), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n865), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(G384));
  AOI211_X1 g0687(.A(new_n523), .B(new_n219), .C1(new_n568), .C2(KEYINPUT35), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(KEYINPUT35), .B2(new_n568), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(KEYINPUT36), .ZN(new_n890));
  OAI21_X1  g0690(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n891));
  OAI22_X1  g0691(.A1(new_n891), .A2(new_n220), .B1(G50), .B2(new_n203), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n892), .A2(G1), .A3(new_n307), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n894), .B(KEYINPUT103), .Z(new_n895));
  NAND2_X1  g0695(.A1(new_n481), .A2(new_n484), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n481), .A2(new_n701), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT37), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n450), .A2(new_n468), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n896), .A2(new_n897), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n444), .A2(new_n297), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n423), .B1(new_n443), .B2(new_n203), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT104), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT16), .B1(new_n902), .B2(new_n903), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n901), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n701), .B1(new_n906), .B2(new_n416), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n484), .B1(new_n906), .B2(new_n416), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n907), .A2(new_n908), .A3(new_n899), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n900), .B1(new_n909), .B2(new_n898), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n494), .B2(new_n907), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT38), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI211_X1 g0713(.A(KEYINPUT38), .B(new_n910), .C1(new_n494), .C2(new_n907), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n361), .A2(new_n711), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n386), .A2(new_n390), .A3(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n361), .B(new_n711), .C1(new_n690), .C2(new_n389), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n859), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n767), .A2(KEYINPUT106), .A3(new_n711), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT106), .B1(new_n767), .B2(new_n711), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n920), .A2(new_n921), .A3(KEYINPUT31), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n767), .A2(new_n772), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n747), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n919), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT40), .B1(new_n915), .B2(new_n926), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n919), .B(KEYINPUT40), .C1(new_n922), .C2(new_n924), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n896), .A2(new_n897), .A3(new_n899), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT37), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n900), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n473), .B1(new_n450), .B2(new_n468), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n471), .B2(new_n469), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n897), .B1(new_n933), .B2(new_n686), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT105), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n931), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AOI211_X1 g0736(.A(KEYINPUT105), .B(new_n897), .C1(new_n933), .C2(new_n686), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n912), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n928), .B1(new_n938), .B2(new_n914), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n927), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n922), .A2(new_n924), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n495), .A2(new_n942), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT107), .Z(new_n944));
  OAI21_X1  g0744(.A(G330), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n944), .B2(new_n941), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n917), .A2(new_n918), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n744), .A2(new_n857), .B1(new_n687), .B2(new_n702), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n915), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n686), .B2(new_n701), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n690), .A2(new_n361), .A3(new_n702), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n491), .B1(KEYINPUT84), .B2(new_n492), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n896), .A2(new_n487), .A3(new_n490), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n933), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n907), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(KEYINPUT38), .B1(new_n957), .B2(new_n910), .ZN(new_n958));
  INV_X1    g0758(.A(new_n914), .ZN(new_n959));
  OAI21_X1  g0759(.A(KEYINPUT39), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT39), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n938), .A2(new_n961), .A3(new_n914), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n952), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n951), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n741), .A2(new_n495), .A3(new_n742), .A4(new_n745), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n693), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n964), .B(new_n966), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n946), .A2(new_n967), .B1(new_n310), .B2(new_n781), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n946), .A2(new_n967), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n895), .B1(new_n968), .B2(new_n969), .ZN(G367));
  INV_X1    g0770(.A(KEYINPUT108), .ZN(new_n971));
  INV_X1    g0771(.A(new_n714), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n735), .B1(new_n585), .B2(new_n702), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n678), .A2(new_n711), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n716), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT45), .ZN(new_n977));
  OR3_X1    g0777(.A1(new_n716), .A2(KEYINPUT44), .A3(new_n975), .ZN(new_n978));
  OAI21_X1  g0778(.A(KEYINPUT44), .B1(new_n716), .B2(new_n975), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OR3_X1    g0780(.A1(new_n972), .A2(new_n977), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n972), .B1(new_n977), .B2(new_n980), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n715), .A2(new_n708), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n713), .B2(new_n715), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n706), .B(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n779), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n719), .B(KEYINPUT41), .Z(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n990), .A2(new_n783), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n973), .A2(new_n538), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n711), .B1(new_n992), .B2(new_n584), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n975), .A2(new_n708), .A3(new_n715), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n993), .B1(new_n994), .B2(KEYINPUT42), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(KEYINPUT42), .B2(new_n994), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n711), .B1(new_n668), .B2(new_n669), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n673), .A2(new_n664), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n664), .B2(new_n997), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n714), .B1(new_n973), .B2(new_n974), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n971), .B1(new_n991), .B2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1003), .B(new_n1004), .Z(new_n1007));
  OAI211_X1 g0807(.A(new_n1007), .B(KEYINPUT108), .C1(new_n783), .C2(new_n990), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n845), .A2(new_n240), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n842), .B1(new_n215), .B2(new_n394), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n787), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n803), .A2(new_n207), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n801), .A2(G143), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n202), .B2(new_n798), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1013), .B(new_n1015), .C1(G159), .C2(new_n791), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n287), .B1(new_n789), .B2(new_n302), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n795), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1017), .B1(G68), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n831), .A2(G137), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n810), .A2(G50), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1016), .A2(new_n1019), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n843), .B1(G303), .B2(new_n819), .ZN(new_n1023));
  XOR2_X1   g0823(.A(KEYINPUT110), .B(G317), .Z(new_n1024));
  OAI221_X1 g0824(.A(new_n1023), .B1(new_n809), .B2(new_n828), .C1(new_n815), .C2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(KEYINPUT109), .B1(new_n798), .B2(new_n523), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1026), .A2(KEYINPUT46), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n791), .A2(G294), .B1(new_n801), .B2(G311), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1026), .A2(KEYINPUT46), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n803), .A2(new_n564), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G107), .B2(new_n1018), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .A4(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1022), .B1(new_n1025), .B2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT47), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1012), .B1(new_n1034), .B2(new_n836), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n999), .B2(new_n852), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1009), .A2(new_n1036), .ZN(G387));
  INV_X1    g0837(.A(new_n986), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n779), .A2(new_n1038), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1039), .A2(new_n719), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n779), .B2(new_n1038), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1038), .A2(new_n783), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n787), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n845), .B1(new_n237), .B2(G45), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n720), .B2(new_n848), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n414), .A2(new_n201), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT50), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n254), .B1(new_n203), .B2(new_n207), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n1047), .A2(new_n720), .A3(new_n1048), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n1045), .A2(new_n1049), .B1(G107), .B2(new_n215), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1043), .B1(new_n1050), .B2(new_n842), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n816), .A2(new_n802), .B1(new_n792), .B2(new_n300), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1030), .B(new_n1052), .C1(G77), .C2(new_n877), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n795), .A2(new_n394), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G50), .B2(new_n819), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT111), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n831), .A2(G150), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n843), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G68), .B2(new_n820), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1053), .A2(new_n1056), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n803), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n843), .B1(G116), .B2(new_n1061), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n795), .A2(new_n828), .B1(new_n798), .B2(new_n822), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1024), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G322), .A2(new_n801), .B1(new_n819), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n791), .A2(G311), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(new_n809), .C2(new_n615), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT48), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1063), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n1068), .B2(new_n1067), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT49), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1062), .B1(new_n829), .B2(new_n815), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1060), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n836), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1051), .B(new_n1075), .C1(new_n713), .C2(new_n852), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n1042), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1041), .A2(new_n1077), .ZN(G393));
  INV_X1    g0878(.A(new_n983), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n783), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n845), .A2(new_n248), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n842), .B1(new_n215), .B2(new_n564), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n787), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1058), .B(new_n875), .C1(new_n831), .C2(G143), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n798), .A2(new_n203), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n795), .A2(new_n207), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(G50), .C2(new_n791), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1084), .B(new_n1087), .C1(new_n300), .C2(new_n809), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G150), .A2(new_n801), .B1(new_n819), .B2(G159), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT51), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G317), .A2(new_n801), .B1(new_n819), .B2(G311), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT52), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n831), .A2(G322), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n877), .A2(G283), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(G116), .A2(new_n1018), .B1(new_n791), .B2(G303), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n270), .B1(new_n806), .B2(new_n822), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(G107), .B2(new_n1061), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .A4(new_n1097), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n1088), .A2(new_n1090), .B1(new_n1092), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1083), .B1(new_n1099), .B2(new_n836), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n975), .B2(new_n852), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1080), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1079), .A2(new_n779), .A3(new_n1038), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1039), .A2(new_n983), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1103), .A2(new_n1104), .A3(new_n719), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT112), .ZN(new_n1106));
  OR2_X1    g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1102), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(G390));
  NAND2_X1  g0910(.A1(new_n737), .A2(new_n702), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(KEYINPUT95), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n737), .A2(new_n729), .A3(new_n702), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1112), .A2(new_n1113), .A3(new_n858), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n857), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n947), .A2(new_n777), .A3(G330), .A4(new_n860), .ZN(new_n1116));
  OAI211_X1 g0916(.A(G330), .B(new_n860), .C1(new_n922), .C2(new_n924), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n947), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1115), .A2(new_n1116), .A3(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n919), .B(G330), .C1(new_n922), .C2(new_n924), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n777), .A2(G330), .A3(new_n860), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n1118), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n949), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1120), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n495), .A2(G330), .A3(new_n942), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1126), .A2(new_n693), .A3(new_n965), .A4(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n952), .B1(new_n948), .B2(new_n1118), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n960), .A2(new_n962), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1116), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n1121), .B2(KEYINPUT113), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n938), .A2(new_n914), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1114), .A2(new_n857), .A3(new_n947), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1133), .A2(new_n1134), .A3(new_n952), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n1130), .A2(new_n1132), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT113), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1121), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n1130), .B2(new_n1135), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1128), .B1(new_n1136), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1130), .A2(new_n1135), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n1138), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n965), .A2(new_n693), .A3(new_n1127), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n948), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1131), .B1(new_n857), .B2(new_n1114), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1145), .B1(new_n1146), .B2(new_n1119), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1130), .A2(new_n1132), .A3(new_n1135), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1143), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1141), .A2(new_n1150), .A3(new_n719), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT114), .ZN(new_n1152));
  OR2_X1    g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NOR3_X1   g0953(.A1(new_n1136), .A2(new_n1140), .A3(new_n782), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n960), .A2(new_n962), .A3(new_n839), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n787), .B1(new_n414), .B2(new_n867), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n287), .B(new_n799), .C1(G116), .C2(new_n819), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1157), .B1(new_n564), .B2(new_n809), .C1(new_n822), .C2(new_n815), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1086), .B1(G68), .B2(new_n1061), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1159), .B1(new_n521), .B2(new_n792), .C1(new_n828), .C2(new_n802), .ZN(new_n1160));
  INV_X1    g0960(.A(G132), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n287), .B1(new_n789), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(G137), .B2(new_n791), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(G159), .A2(new_n1018), .B1(new_n801), .B2(G128), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1061), .A2(G50), .ZN(new_n1165));
  OAI21_X1  g0965(.A(KEYINPUT53), .B1(new_n798), .B2(new_n302), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  OR3_X1    g0967(.A1(new_n798), .A2(KEYINPUT53), .A3(new_n302), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT54), .B(G143), .ZN(new_n1169));
  INV_X1    g0969(.A(G125), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1168), .B1(new_n809), .B2(new_n1169), .C1(new_n815), .C2(new_n1170), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n1158), .A2(new_n1160), .B1(new_n1167), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1156), .B1(new_n1172), .B2(new_n836), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1154), .B1(new_n1155), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1153), .A2(new_n1174), .A3(new_n1175), .ZN(G378));
  INV_X1    g0976(.A(KEYINPUT57), .ZN(new_n1177));
  OR2_X1    g0977(.A1(new_n951), .A2(new_n963), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n701), .B1(new_n314), .B2(new_n315), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n332), .B2(new_n337), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1179), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n685), .B(new_n1182), .C1(new_n323), .C2(new_n331), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT119), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1181), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1187));
  OAI21_X1  g0987(.A(KEYINPUT119), .B1(new_n1180), .B2(new_n1183), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1187), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n940), .B2(G330), .ZN(new_n1193));
  INV_X1    g0993(.A(G330), .ZN(new_n1194));
  NOR4_X1   g0994(.A1(new_n927), .A2(new_n1191), .A3(new_n939), .A4(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1178), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n939), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n925), .B1(new_n913), .B2(new_n914), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1197), .B(G330), .C1(KEYINPUT40), .C2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n1191), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n940), .A2(G330), .A3(new_n1192), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1200), .A2(new_n964), .A3(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1177), .B1(new_n1196), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT121), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1144), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n1150), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1204), .B1(new_n1150), .B2(new_n1205), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1203), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT122), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1203), .B(KEYINPUT122), .C1(new_n1206), .C2(new_n1207), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1136), .A2(new_n1128), .A3(new_n1140), .ZN(new_n1213));
  OAI21_X1  g1013(.A(KEYINPUT121), .B1(new_n1213), .B2(new_n1144), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1150), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1215));
  OAI21_X1  g1015(.A(KEYINPUT120), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n964), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1178), .B(KEYINPUT120), .C1(new_n1193), .C2(new_n1195), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1214), .A2(new_n1215), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n719), .B1(new_n1219), .B2(KEYINPUT57), .ZN(new_n1220));
  OR2_X1    g1020(.A1(new_n1212), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n782), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n866), .A2(new_n201), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n784), .A2(new_n1223), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n803), .A2(new_n202), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n802), .A2(new_n523), .B1(new_n798), .B2(new_n207), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1225), .B(new_n1226), .C1(G97), .C2(new_n791), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n253), .B1(new_n806), .B2(new_n394), .C1(new_n521), .C2(new_n789), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n843), .B(new_n1228), .C1(G68), .C2(new_n1018), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1227), .B(new_n1229), .C1(new_n828), .C2(new_n815), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT58), .ZN(new_n1231));
  AOI21_X1  g1031(.A(G41), .B1(new_n843), .B2(G33), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1169), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(G128), .A2(new_n819), .B1(new_n877), .B2(new_n1233), .ZN(new_n1234));
  XOR2_X1   g1034(.A(new_n1234), .B(KEYINPUT115), .Z(new_n1235));
  AOI22_X1  g1035(.A1(new_n1018), .A2(G150), .B1(new_n820), .B2(G137), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n791), .A2(G132), .B1(new_n801), .B2(G125), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  XOR2_X1   g1038(.A(new_n1238), .B(KEYINPUT59), .Z(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(KEYINPUT116), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n831), .A2(G124), .ZN(new_n1241));
  AOI211_X1 g1041(.A(G33), .B(G41), .C1(new_n1061), .C2(G159), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1239), .A2(KEYINPUT116), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1231), .B1(G50), .B2(new_n1232), .C1(new_n1243), .C2(new_n1244), .ZN(new_n1245));
  XOR2_X1   g1045(.A(new_n1245), .B(KEYINPUT117), .Z(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n836), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT118), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1224), .B(new_n1248), .C1(new_n839), .C2(new_n1191), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1222), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1221), .A2(new_n1250), .ZN(G375));
  NAND2_X1  g1051(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1128), .A2(new_n1252), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1253), .A2(new_n988), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1254), .B(KEYINPUT123), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1118), .A2(new_n839), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n787), .B1(G68), .B2(new_n867), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n802), .A2(new_n822), .B1(new_n798), .B2(new_n564), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n1054), .B(new_n1258), .C1(G116), .C2(new_n791), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n810), .A2(G107), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n831), .A2(G303), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n287), .B(new_n1013), .C1(G283), .C2(new_n819), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .A4(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n843), .B1(new_n302), .B2(new_n806), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1225), .B1(G50), .B2(new_n1018), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n816), .B2(new_n798), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n1264), .B(new_n1266), .C1(G128), .C2(new_n831), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT124), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n802), .A2(new_n1161), .B1(new_n869), .B2(new_n789), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(new_n791), .B2(new_n1233), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1267), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1271));
  AND2_X1   g1071(.A1(new_n1270), .A2(new_n1268), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1263), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1257), .B1(new_n1273), .B2(new_n836), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n1126), .A2(new_n783), .B1(new_n1256), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1255), .A2(new_n1275), .ZN(G381));
  NAND3_X1  g1076(.A1(new_n1009), .A2(new_n1036), .A3(new_n1109), .ZN(new_n1277));
  AND2_X1   g1077(.A1(new_n1174), .A2(new_n1151), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(G393), .A2(G396), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1278), .A2(new_n1279), .A3(new_n886), .ZN(new_n1280));
  OR4_X1    g1080(.A1(G375), .A2(G381), .A3(new_n1277), .A4(new_n1280), .ZN(G407));
  INV_X1    g1081(.A(G375), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n698), .A2(G343), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1282), .A2(new_n1278), .A3(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(G407), .A2(G213), .A3(new_n1284), .ZN(G409));
  OAI211_X1 g1085(.A(G378), .B(new_n1250), .C1(new_n1212), .C2(new_n1220), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1219), .A2(new_n989), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n782), .B1(new_n1196), .B2(new_n1202), .ZN(new_n1288));
  OR2_X1    g1088(.A1(new_n1249), .A2(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1278), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1286), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT127), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1283), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1253), .A2(KEYINPUT60), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT60), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1252), .A2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1294), .A2(new_n719), .A3(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1275), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n886), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1297), .A2(G384), .A3(new_n1275), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT126), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1299), .A2(KEYINPUT126), .A3(new_n1300), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n1303), .A2(new_n1304), .A3(KEYINPUT63), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1291), .A2(new_n1292), .A3(new_n1293), .A4(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n854), .B1(new_n1041), .B2(new_n1077), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1279), .A2(new_n1307), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1009), .A2(new_n1036), .A3(new_n1109), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1109), .B1(new_n1009), .B2(new_n1036), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1308), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(G387), .A2(G390), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1308), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1312), .A2(new_n1277), .A3(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT61), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1311), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1306), .A2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1283), .B1(new_n1286), .B2(new_n1290), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1292), .B1(new_n1318), .B2(new_n1305), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1317), .A2(new_n1319), .ZN(new_n1320));
  AND3_X1   g1120(.A1(new_n1286), .A2(KEYINPUT125), .A3(new_n1290), .ZN(new_n1321));
  AOI21_X1  g1121(.A(KEYINPUT125), .B1(new_n1286), .B2(new_n1290), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1293), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1283), .A2(G2897), .ZN(new_n1325));
  AND2_X1   g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1301), .A2(new_n1325), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1323), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1324), .ZN(new_n1329));
  OAI211_X1 g1129(.A(new_n1293), .B(new_n1329), .C1(new_n1321), .C2(new_n1322), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT63), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1320), .A2(new_n1328), .A3(new_n1332), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1315), .B1(new_n1334), .B2(new_n1318), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT62), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1330), .A2(new_n1336), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1318), .A2(KEYINPUT62), .A3(new_n1329), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1335), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1311), .A2(new_n1314), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1340), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1333), .B1(new_n1339), .B2(new_n1341), .ZN(G405));
  INV_X1    g1142(.A(new_n1278), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1286), .B1(new_n1282), .B2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1344), .A2(new_n1329), .ZN(new_n1345));
  OAI211_X1 g1145(.A(new_n1301), .B(new_n1286), .C1(new_n1282), .C2(new_n1343), .ZN(new_n1346));
  AND3_X1   g1146(.A1(new_n1345), .A2(new_n1340), .A3(new_n1346), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1340), .B1(new_n1345), .B2(new_n1346), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(new_n1347), .A2(new_n1348), .ZN(G402));
endmodule


