//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 0 1 0 0 1 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 1 1 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 0 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1269, new_n1270, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1339, new_n1340;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n204), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G77), .ZN(new_n208));
  INV_X1    g0008(.A(G244), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G68), .A2(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G107), .ZN(new_n213));
  INV_X1    g0013(.A(G264), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n211), .B(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n210), .B(new_n215), .C1(G116), .C2(G270), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G58), .A2(G232), .ZN(new_n217));
  INV_X1    g0017(.A(G50), .ZN(new_n218));
  INV_X1    g0018(.A(G226), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n216), .B(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G1), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n220), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT1), .Z(new_n226));
  NAND2_X1  g0026(.A1(new_n204), .A2(new_n205), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n227), .A2(new_n218), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n228), .A2(G20), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n224), .A2(G13), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n232), .B(G250), .C1(G257), .C2(G264), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT0), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n226), .A2(new_n231), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT65), .ZN(G361));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n214), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(KEYINPUT66), .B(G50), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G58), .ZN(new_n246));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G97), .B(G107), .Z(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(KEYINPUT73), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT68), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT68), .ZN(new_n256));
  NAND4_X1  g0056(.A1(new_n256), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(new_n229), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT69), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n255), .A2(new_n257), .A3(KEYINPUT69), .A4(new_n229), .ZN(new_n261));
  AND2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n222), .B1(new_n227), .B2(new_n218), .ZN(new_n263));
  XOR2_X1   g0063(.A(KEYINPUT8), .B(G58), .Z(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n222), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(G150), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G20), .A2(G33), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  OAI22_X1  g0069(.A1(new_n265), .A2(new_n266), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n262), .B1(new_n263), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n221), .A2(G13), .A3(G20), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT70), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n221), .A2(KEYINPUT70), .A3(G13), .A4(G20), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n271), .B1(G50), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n260), .A2(new_n261), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n221), .A2(G20), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n278), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(new_n218), .ZN(new_n281));
  OR2_X1    g0081(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT3), .B(G33), .ZN(new_n283));
  INV_X1    g0083(.A(G223), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  AND2_X1   g0085(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n286));
  NOR2_X1   g0086(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G222), .ZN(new_n289));
  OAI221_X1 g0089(.A(new_n283), .B1(new_n284), .B2(new_n285), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(G1), .A3(G13), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n290), .B(new_n293), .C1(G77), .C2(new_n283), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n221), .B(G274), .C1(G41), .C2(G45), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n221), .B1(G41), .B2(G45), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G226), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n294), .A2(new_n295), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G169), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n299), .ZN(new_n302));
  INV_X1    g0102(.A(G179), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n282), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  OAI22_X1  g0105(.A1(new_n265), .A2(new_n269), .B1(new_n222), .B2(new_n208), .ZN(new_n306));
  XOR2_X1   g0106(.A(KEYINPUT15), .B(G87), .Z(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(new_n266), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n258), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n276), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n208), .ZN(new_n312));
  AND3_X1   g0112(.A1(new_n255), .A2(new_n229), .A3(new_n257), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n313), .A2(new_n276), .A3(new_n279), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n310), .B(new_n312), .C1(new_n208), .C2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G33), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT3), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT3), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G33), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G107), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT67), .B(G1698), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n322), .A2(G232), .B1(G238), .B2(G1698), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n321), .B1(new_n323), .B2(new_n320), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT71), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n292), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(new_n325), .B2(new_n324), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n297), .A2(G244), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n327), .A2(new_n295), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n315), .B1(new_n329), .B2(G190), .ZN(new_n330));
  INV_X1    g0130(.A(G200), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n330), .B1(new_n331), .B2(new_n329), .ZN(new_n332));
  OR3_X1    g0132(.A1(new_n277), .A2(KEYINPUT9), .A3(new_n281), .ZN(new_n333));
  OAI21_X1  g0133(.A(KEYINPUT9), .B1(new_n277), .B2(new_n281), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT72), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(new_n302), .B2(new_n331), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n299), .A2(KEYINPUT72), .A3(G200), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n337), .A2(new_n338), .B1(G190), .B2(new_n302), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT10), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n335), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n340), .B1(new_n335), .B2(new_n339), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n305), .B(new_n332), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n329), .A2(new_n303), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n327), .A2(new_n295), .A3(new_n328), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n300), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n345), .A2(new_n347), .A3(new_n315), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n253), .B1(new_n344), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n305), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n335), .A2(new_n339), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT10), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n351), .B1(new_n353), .B2(new_n341), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n354), .A2(KEYINPUT73), .A3(new_n348), .A4(new_n332), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n322), .A2(G226), .B1(G232), .B2(G1698), .ZN(new_n356));
  INV_X1    g0156(.A(G97), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n356), .A2(new_n320), .B1(new_n316), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n293), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n297), .A2(G238), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(new_n360), .A3(new_n295), .ZN(new_n361));
  XNOR2_X1  g0161(.A(KEYINPUT74), .B(KEYINPUT13), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  AND3_X1   g0164(.A1(new_n359), .A2(new_n360), .A3(new_n295), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n365), .A2(KEYINPUT75), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT75), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT13), .B1(new_n361), .B2(new_n367), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n364), .B(G190), .C1(new_n366), .C2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n203), .A2(G20), .ZN(new_n370));
  OAI221_X1 g0170(.A(new_n370), .B1(new_n266), .B2(new_n208), .C1(new_n269), .C2(new_n218), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n262), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g0172(.A(KEYINPUT76), .B(KEYINPUT11), .ZN(new_n373));
  XNOR2_X1  g0173(.A(new_n372), .B(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n311), .A2(new_n203), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n375), .B(KEYINPUT12), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(new_n203), .B2(new_n314), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n361), .A2(new_n362), .ZN(new_n379));
  OAI21_X1  g0179(.A(G200), .B1(new_n379), .B2(new_n363), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n369), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(G169), .B1(new_n379), .B2(new_n363), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT14), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n364), .B(G179), .C1(new_n366), .C2(new_n368), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT14), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n386), .B(G169), .C1(new_n379), .C2(new_n363), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n378), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n382), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI22_X1  g0190(.A1(new_n288), .A2(new_n284), .B1(new_n219), .B2(new_n285), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n318), .A2(G33), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT77), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(new_n316), .B2(KEYINPUT3), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n318), .A2(KEYINPUT77), .A3(G33), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n392), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n391), .A2(new_n396), .B1(G33), .B2(G87), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT78), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n292), .A2(G232), .A3(new_n296), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n398), .B1(new_n399), .B2(new_n295), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n399), .A2(new_n398), .A3(new_n295), .ZN(new_n401));
  OAI22_X1  g0201(.A1(new_n397), .A2(new_n292), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n402), .A2(G179), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n322), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n404));
  AND3_X1   g0204(.A1(new_n318), .A2(KEYINPUT77), .A3(G33), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT77), .B1(new_n318), .B2(G33), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n317), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(G87), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n404), .A2(new_n407), .B1(new_n316), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n293), .ZN(new_n410));
  INV_X1    g0210(.A(new_n400), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n399), .A2(new_n398), .A3(new_n295), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(G169), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT79), .B1(new_n403), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n402), .A2(new_n300), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT79), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n410), .A2(new_n413), .A3(new_n303), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT7), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n407), .A2(new_n420), .A3(new_n222), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT7), .B1(new_n396), .B2(G20), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n422), .A3(G68), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n204), .B(new_n205), .C1(new_n202), .C2(new_n203), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n424), .A2(G20), .B1(G159), .B2(new_n268), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(KEYINPUT16), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT16), .ZN(new_n427));
  INV_X1    g0227(.A(new_n425), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n420), .B1(new_n283), .B2(G20), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n320), .A2(KEYINPUT7), .A3(new_n222), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n203), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n427), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n426), .A2(new_n432), .A3(new_n258), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n280), .A2(new_n264), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n265), .A2(new_n276), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n415), .A2(new_n419), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT18), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n415), .A2(new_n437), .A3(KEYINPUT18), .A4(new_n419), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n402), .A2(G200), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n410), .A2(new_n413), .A3(G190), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n433), .A2(new_n436), .A3(new_n443), .A4(new_n444), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n445), .B(KEYINPUT17), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n350), .A2(new_n355), .A3(new_n390), .A4(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT22), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n222), .A2(G87), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n450), .B1(new_n320), .B2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n396), .A2(KEYINPUT22), .A3(new_n222), .A4(G87), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G116), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT83), .B1(new_n454), .B2(G20), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT83), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n456), .A2(new_n222), .A3(G33), .A4(G116), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT84), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT23), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(new_n222), .B2(G107), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n213), .A2(KEYINPUT23), .A3(G20), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n458), .A2(new_n459), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n459), .B1(new_n458), .B2(new_n463), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n452), .B(new_n453), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT24), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n458), .A2(new_n463), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT84), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n458), .A2(new_n459), .A3(new_n463), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n472), .A2(KEYINPUT24), .A3(new_n452), .A4(new_n453), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n468), .A2(new_n473), .A3(new_n258), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n221), .A2(G33), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n278), .A2(new_n276), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G107), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n276), .A2(G107), .ZN(new_n478));
  XNOR2_X1  g0278(.A(new_n478), .B(KEYINPUT25), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n474), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n221), .A2(G45), .ZN(new_n481));
  OR2_X1    g0281(.A1(KEYINPUT5), .A2(G41), .ZN(new_n482));
  NAND2_X1  g0282(.A1(KEYINPUT5), .A2(G41), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(new_n293), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G264), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(G274), .ZN(new_n487));
  INV_X1    g0287(.A(G294), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n316), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(G250), .B1(new_n286), .B2(new_n287), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G257), .A2(G1698), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n489), .B1(new_n492), .B2(new_n396), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n486), .B(new_n487), .C1(new_n493), .C2(new_n292), .ZN(new_n494));
  OR3_X1    g0294(.A1(new_n494), .A2(KEYINPUT86), .A3(G190), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n331), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT87), .ZN(new_n497));
  OAI21_X1  g0297(.A(KEYINPUT86), .B1(new_n494), .B2(G190), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT87), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n494), .A2(new_n499), .A3(new_n331), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n495), .A2(new_n497), .A3(new_n498), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n480), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n474), .A2(new_n477), .A3(new_n479), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n494), .A2(G169), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT85), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n492), .A2(new_n396), .ZN(new_n507));
  INV_X1    g0307(.A(new_n489), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n509), .A2(new_n293), .B1(G264), .B2(new_n485), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(G179), .A3(new_n487), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n494), .A2(KEYINPUT85), .A3(G169), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n506), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n503), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n502), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT88), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT88), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n502), .A2(new_n517), .A3(new_n514), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NOR3_X1   g0319(.A1(new_n283), .A2(new_n420), .A3(G20), .ZN(new_n520));
  AOI21_X1  g0320(.A(KEYINPUT7), .B1(new_n320), .B2(new_n222), .ZN(new_n521));
  OAI21_X1  g0321(.A(G107), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n213), .A2(KEYINPUT6), .A3(G97), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n357), .A2(new_n213), .ZN(new_n524));
  NOR2_X1   g0324(.A1(G97), .A2(G107), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n523), .B1(new_n526), .B2(KEYINPUT6), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G20), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n268), .A2(G77), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n522), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  AOI22_X1  g0330(.A1(G97), .A2(new_n476), .B1(new_n530), .B2(new_n258), .ZN(new_n531));
  OAI211_X1 g0331(.A(KEYINPUT4), .B(G244), .C1(new_n286), .C2(new_n287), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G250), .A2(G1698), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n534), .A2(new_n283), .B1(G33), .B2(G283), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT4), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n322), .A2(G244), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n536), .B1(new_n407), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n293), .ZN(new_n540));
  INV_X1    g0340(.A(G45), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n541), .A2(G1), .ZN(new_n542));
  INV_X1    g0342(.A(new_n483), .ZN(new_n543));
  NOR2_X1   g0343(.A1(KEYINPUT5), .A2(G41), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n545), .A2(G257), .A3(new_n292), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT80), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n546), .A2(new_n487), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n547), .B1(new_n546), .B2(new_n487), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n540), .A2(G190), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n546), .A2(new_n487), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT80), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n546), .A2(new_n487), .A3(new_n547), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n292), .B1(new_n535), .B2(new_n538), .ZN(new_n556));
  OAI21_X1  g0356(.A(G200), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n311), .A2(new_n357), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n531), .A2(new_n551), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n530), .A2(new_n258), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n278), .A2(G97), .A3(new_n276), .A4(new_n475), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n300), .B1(new_n555), .B2(new_n556), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n540), .A2(new_n303), .A3(new_n550), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n559), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(G257), .ZN(new_n567));
  OR2_X1    g0367(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n568));
  NAND2_X1  g0368(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n214), .A2(new_n285), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n396), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n320), .A2(G303), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n292), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n545), .A2(G270), .A3(new_n292), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n487), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G190), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n331), .B2(new_n577), .ZN(new_n579));
  AOI21_X1  g0379(.A(G20), .B1(new_n316), .B2(G97), .ZN(new_n580));
  INV_X1    g0380(.A(G283), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n580), .B1(new_n316), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(G116), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(G20), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n258), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT20), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n258), .A2(new_n582), .A3(KEYINPUT20), .A4(new_n584), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n274), .A2(new_n583), .A3(new_n275), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n583), .B1(new_n221), .B2(G33), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n313), .A2(new_n276), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n579), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(G190), .ZN(new_n595));
  OR2_X1    g0395(.A1(new_n481), .A2(G274), .ZN(new_n596));
  INV_X1    g0396(.A(G250), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n481), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n596), .A2(new_n292), .A3(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n454), .ZN(new_n600));
  OAI21_X1  g0400(.A(G238), .B1(new_n286), .B2(new_n287), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n209), .A2(new_n285), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n600), .B1(new_n604), .B2(new_n396), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n595), .B(new_n599), .C1(new_n605), .C2(new_n292), .ZN(new_n606));
  INV_X1    g0406(.A(new_n599), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n602), .B1(new_n322), .B2(G238), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n454), .B1(new_n608), .B2(new_n407), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n607), .B1(new_n609), .B2(new_n293), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n606), .B1(new_n610), .B2(G200), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n394), .A2(new_n395), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n612), .A2(new_n222), .A3(G68), .A4(new_n317), .ZN(new_n613));
  XOR2_X1   g0413(.A(KEYINPUT81), .B(KEYINPUT19), .Z(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(new_n357), .B2(new_n266), .ZN(new_n615));
  XNOR2_X1  g0415(.A(KEYINPUT82), .B(G87), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n616), .A2(G97), .A3(G107), .ZN(new_n617));
  XNOR2_X1  g0417(.A(KEYINPUT81), .B(KEYINPUT19), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n316), .A2(new_n357), .ZN(new_n619));
  AOI21_X1  g0419(.A(G20), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n613), .B(new_n615), .C1(new_n617), .C2(new_n620), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n621), .A2(new_n258), .B1(new_n311), .B2(new_n308), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n476), .A2(G87), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n611), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n621), .A2(new_n258), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n278), .A2(new_n276), .A3(new_n475), .A4(new_n307), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n311), .A2(new_n308), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n610), .A2(new_n303), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n599), .B1(new_n605), .B2(new_n292), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n300), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n628), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n624), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT21), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n592), .A2(new_n590), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n635), .B1(new_n587), .B2(new_n588), .ZN(new_n636));
  OAI21_X1  g0436(.A(G169), .B1(new_n574), .B2(new_n576), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n634), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n571), .B1(new_n322), .B2(G257), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n573), .B1(new_n639), .B2(new_n407), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n293), .ZN(new_n641));
  INV_X1    g0441(.A(new_n576), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n300), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n643), .A2(new_n593), .A3(KEYINPUT21), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n593), .A2(G179), .A3(new_n577), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n638), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NOR4_X1   g0446(.A1(new_n566), .A2(new_n594), .A3(new_n633), .A4(new_n646), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n449), .A2(new_n519), .A3(new_n647), .ZN(G372));
  AOI22_X1  g0448(.A1(new_n388), .A2(new_n389), .B1(new_n349), .B2(new_n381), .ZN(new_n649));
  INV_X1    g0449(.A(new_n446), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n442), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n353), .A2(new_n341), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n351), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  INV_X1    g0454(.A(new_n565), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n624), .A2(new_n632), .A3(KEYINPUT89), .ZN(new_n656));
  AOI21_X1  g0456(.A(KEYINPUT89), .B1(new_n624), .B2(new_n632), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n654), .B(new_n655), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT26), .B1(new_n633), .B2(new_n565), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n658), .A2(new_n632), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n566), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT89), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n633), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n624), .A2(new_n632), .A3(KEYINPUT89), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n663), .A2(new_n664), .B1(new_n480), .B2(new_n501), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT90), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n646), .B(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n514), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n661), .B(new_n665), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n660), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n653), .B1(new_n448), .B2(new_n671), .ZN(G369));
  NAND3_X1  g0472(.A1(new_n221), .A2(new_n222), .A3(G13), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n503), .A2(new_n678), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n502), .A2(new_n517), .A3(new_n514), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n517), .B1(new_n502), .B2(new_n514), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n668), .A2(new_n678), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n678), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n636), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n667), .A2(new_n687), .ZN(new_n688));
  OR3_X1    g0488(.A1(new_n594), .A2(new_n646), .A3(new_n687), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G330), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n638), .A2(new_n644), .A3(new_n645), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(new_n678), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n696), .B1(new_n516), .B2(new_n518), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n514), .A2(new_n678), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n693), .A2(new_n699), .ZN(G399));
  INV_X1    g0500(.A(new_n232), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G41), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G1), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n617), .A2(new_n583), .ZN(new_n705));
  INV_X1    g0505(.A(new_n228), .ZN(new_n706));
  OAI22_X1  g0506(.A1(new_n704), .A2(new_n705), .B1(new_n706), .B2(new_n703), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT28), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n663), .A2(new_n664), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n514), .A2(new_n694), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(new_n502), .A3(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT93), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n566), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n559), .A2(new_n565), .A3(KEYINPUT93), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n655), .A2(new_n654), .A3(new_n632), .A4(new_n624), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n565), .B1(new_n663), .B2(new_n664), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n632), .B(new_n717), .C1(new_n718), .C2(new_n654), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n686), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(KEYINPUT94), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT94), .ZN(new_n722));
  OAI211_X1 g0522(.A(new_n722), .B(new_n686), .C1(new_n716), .C2(new_n719), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n721), .A2(KEYINPUT29), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n678), .B1(new_n660), .B2(new_n669), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT29), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT92), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n555), .A2(new_n556), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n577), .A2(G179), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n730), .A2(new_n731), .A3(new_n494), .A4(new_n630), .ZN(new_n732));
  NOR4_X1   g0532(.A1(new_n630), .A2(new_n574), .A3(new_n303), .A4(new_n576), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n733), .A2(new_n729), .A3(KEYINPUT30), .A4(new_n510), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT30), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n540), .A2(new_n510), .A3(new_n550), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n577), .A2(G179), .A3(new_n610), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n732), .A2(new_n734), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n739), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n733), .A2(new_n729), .A3(new_n510), .ZN(new_n741));
  AOI21_X1  g0541(.A(KEYINPUT91), .B1(new_n741), .B2(new_n735), .ZN(new_n742));
  OAI211_X1 g0542(.A(KEYINPUT91), .B(new_n735), .C1(new_n736), .C2(new_n737), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n732), .A2(new_n734), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n686), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n728), .B(new_n740), .C1(new_n747), .C2(KEYINPUT31), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT91), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n738), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n750), .A2(new_n734), .A3(new_n732), .A4(new_n743), .ZN(new_n751));
  AOI21_X1  g0551(.A(KEYINPUT31), .B1(new_n751), .B2(new_n678), .ZN(new_n752));
  INV_X1    g0552(.A(new_n740), .ZN(new_n753));
  OAI21_X1  g0553(.A(KEYINPUT92), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n647), .B(new_n686), .C1(new_n680), .C2(new_n681), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n748), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G330), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n724), .A2(new_n727), .A3(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n708), .B1(new_n759), .B2(G1), .ZN(G364));
  INV_X1    g0560(.A(new_n691), .ZN(new_n761));
  INV_X1    g0561(.A(G13), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n704), .B1(G45), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(G330), .B2(new_n690), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n229), .B1(G20), .B2(new_n300), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G179), .A2(G200), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n222), .B1(new_n769), .B2(G190), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n488), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n303), .A2(new_n331), .ZN(new_n772));
  NAND2_X1  g0572(.A1(G20), .A2(G190), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(KEYINPUT97), .B(G326), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n595), .A2(G20), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(new_n772), .ZN(new_n779));
  XOR2_X1   g0579(.A(KEYINPUT33), .B(G317), .Z(new_n780));
  OAI221_X1 g0580(.A(new_n320), .B1(new_n775), .B2(new_n776), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n777), .A2(new_n303), .A3(G200), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n771), .B(new_n781), .C1(G311), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n778), .A2(new_n769), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n773), .A2(new_n303), .A3(G200), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n785), .A2(G329), .B1(G322), .B2(new_n786), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n331), .A2(G179), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n778), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G303), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n789), .A2(new_n774), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n788), .B1(new_n581), .B2(new_n790), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n770), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G97), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n203), .B2(new_n779), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(KEYINPUT96), .ZN(new_n797));
  INV_X1    g0597(.A(new_n792), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n320), .B1(new_n798), .B2(new_n616), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(new_n213), .B2(new_n790), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n782), .A2(G77), .B1(new_n786), .B2(G58), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT95), .ZN(new_n803));
  INV_X1    g0603(.A(new_n775), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n796), .A2(KEYINPUT96), .B1(G50), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G159), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n784), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT32), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n801), .A2(new_n803), .A3(new_n805), .A4(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n768), .B1(new_n793), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n228), .A2(new_n541), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n701), .A2(new_n396), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n811), .B(new_n812), .C1(new_n248), .C2(new_n541), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n232), .A2(G355), .A3(new_n283), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n813), .B(new_n814), .C1(G116), .C2(new_n232), .ZN(new_n815));
  NOR2_X1   g0615(.A1(G13), .A2(G33), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(G20), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(new_n767), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n818), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n820), .B(new_n764), .C1(new_n690), .C2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n766), .B1(new_n810), .B2(new_n822), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT98), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(G396));
  NOR2_X1   g0625(.A1(new_n767), .A2(new_n816), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n782), .A2(G159), .B1(new_n786), .B2(G143), .ZN(new_n828));
  INV_X1    g0628(.A(G137), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n828), .B1(new_n829), .B2(new_n775), .C1(new_n267), .C2(new_n779), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT34), .Z(new_n831));
  AOI211_X1 g0631(.A(new_n407), .B(new_n831), .C1(G132), .C2(new_n785), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n794), .A2(G58), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n798), .A2(G50), .ZN(new_n834));
  INV_X1    g0634(.A(new_n790), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(G68), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n832), .A2(new_n833), .A3(new_n834), .A4(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(G311), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n795), .B1(new_n581), .B2(new_n779), .C1(new_n838), .C2(new_n784), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n835), .A2(G87), .ZN(new_n840));
  INV_X1    g0640(.A(new_n782), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n583), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n320), .B1(new_n792), .B2(new_n213), .ZN(new_n843));
  NOR3_X1   g0643(.A1(new_n839), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n786), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n844), .B1(new_n488), .B2(new_n845), .C1(new_n791), .C2(new_n775), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n837), .A2(new_n846), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n764), .B1(G77), .B2(new_n827), .C1(new_n847), .C2(new_n768), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT99), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n315), .A2(new_n678), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT100), .Z(new_n851));
  NAND2_X1  g0651(.A1(new_n332), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n348), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n348), .A2(new_n678), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n849), .B1(new_n816), .B2(new_n856), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT101), .Z(new_n858));
  XNOR2_X1  g0658(.A(new_n725), .B(new_n856), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(new_n757), .ZN(new_n860));
  INV_X1    g0660(.A(new_n764), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n858), .A2(new_n862), .ZN(G384));
  NAND2_X1  g0663(.A1(new_n724), .A2(new_n727), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n449), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT104), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n864), .A2(KEYINPUT104), .A3(new_n449), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n653), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n388), .A2(new_n389), .A3(new_n686), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT39), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT38), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n423), .A2(new_n425), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n278), .B1(new_n875), .B2(new_n427), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n876), .A2(new_n426), .B1(new_n434), .B2(new_n435), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n403), .A2(new_n414), .A3(KEYINPUT79), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n417), .B1(new_n416), .B2(new_n418), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n445), .B1(new_n877), .B2(new_n676), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT37), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT37), .ZN(new_n883));
  INV_X1    g0683(.A(new_n676), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n437), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n438), .A2(new_n883), .A3(new_n445), .A4(new_n885), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  OR2_X1    g0687(.A1(new_n877), .A2(new_n676), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n442), .B2(new_n446), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n874), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n882), .A2(new_n886), .ZN(new_n891));
  OAI211_X1 g0691(.A(KEYINPUT38), .B(new_n891), .C1(new_n447), .C2(new_n888), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n438), .A2(new_n445), .A3(new_n885), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT37), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n895), .A2(new_n886), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n885), .B1(new_n442), .B2(new_n446), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n874), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT103), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n873), .B1(new_n893), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT103), .ZN(new_n901));
  AND4_X1   g0701(.A1(new_n901), .A2(new_n898), .A3(new_n892), .A4(new_n873), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n872), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n440), .A2(new_n441), .A3(new_n676), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT102), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n854), .B1(new_n852), .B2(new_n348), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n854), .B1(new_n725), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n388), .A2(new_n389), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n389), .A2(new_n678), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n908), .A2(new_n381), .A3(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n389), .B(new_n678), .C1(new_n382), .C2(new_n388), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n905), .B1(new_n907), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n670), .A2(new_n686), .A3(new_n906), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n855), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n916), .A2(KEYINPUT102), .A3(new_n912), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n890), .A2(new_n892), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n914), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n903), .A2(new_n904), .A3(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n870), .B(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT106), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n856), .B1(new_n910), .B2(new_n911), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n751), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n925), .A2(new_n752), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT105), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n926), .A2(new_n927), .A3(new_n755), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n927), .B1(new_n926), .B2(new_n755), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n918), .B(new_n924), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT40), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n912), .A2(new_n906), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n747), .A2(KEYINPUT31), .ZN(new_n933));
  INV_X1    g0733(.A(new_n752), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n755), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT105), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n926), .A2(new_n927), .A3(new_n755), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n932), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n931), .B1(new_n898), .B2(new_n892), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n930), .A2(new_n931), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n928), .A2(new_n929), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n941), .A2(new_n448), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n940), .B(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(G330), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n923), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n921), .B(KEYINPUT106), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n946), .B1(new_n221), .B2(new_n763), .C1(new_n947), .C2(new_n945), .ZN(new_n948));
  OAI211_X1 g0748(.A(G20), .B(new_n230), .C1(new_n527), .C2(KEYINPUT35), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n583), .B(new_n949), .C1(KEYINPUT35), .C2(new_n527), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT36), .Z(new_n951));
  OAI21_X1  g0751(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n706), .A2(new_n952), .B1(G50), .B2(new_n203), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(G1), .A3(new_n762), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n948), .A2(new_n951), .A3(new_n954), .ZN(G367));
  INV_X1    g0755(.A(new_n812), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n819), .B1(new_n232), .B2(new_n308), .C1(new_n243), .C2(new_n956), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n784), .A2(new_n829), .B1(new_n792), .B2(new_n202), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT109), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n845), .A2(new_n267), .B1(new_n790), .B2(new_n208), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(G68), .B2(new_n794), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n320), .B1(new_n804), .B2(G143), .ZN(new_n962));
  AND3_X1   g0762(.A1(new_n959), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n963), .B1(new_n218), .B2(new_n841), .C1(new_n806), .C2(new_n779), .ZN(new_n964));
  INV_X1    g0764(.A(G317), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n784), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n798), .A2(G116), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT46), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n407), .B1(new_n357), .B2(new_n790), .ZN(new_n969));
  INV_X1    g0769(.A(new_n779), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n969), .B1(G294), .B2(new_n970), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n782), .A2(G283), .B1(new_n786), .B2(G303), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n804), .A2(G311), .B1(new_n794), .B2(G107), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n968), .A2(new_n971), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n964), .B1(new_n966), .B2(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT47), .Z(new_n976));
  OAI211_X1 g0776(.A(new_n764), .B(new_n957), .C1(new_n976), .C2(new_n768), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n623), .A2(new_n622), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n678), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n709), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n632), .B2(new_n979), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n977), .B1(new_n982), .B2(new_n818), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n221), .B1(new_n763), .B2(G45), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT44), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n713), .A2(new_n714), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n562), .A2(new_n678), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n988), .A2(new_n989), .B1(new_n655), .B2(new_n678), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT108), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n990), .B(new_n991), .C1(new_n697), .C2(new_n698), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n695), .B1(new_n680), .B2(new_n681), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n514), .B2(new_n678), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n991), .B1(new_n995), .B2(new_n990), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n987), .B1(new_n993), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n990), .ZN(new_n998));
  OAI21_X1  g0798(.A(KEYINPUT108), .B1(new_n699), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n999), .A2(KEYINPUT44), .A3(new_n992), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT45), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n995), .B2(new_n990), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n699), .A2(new_n998), .A3(KEYINPUT45), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n997), .A2(new_n1000), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n692), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n997), .A2(new_n1000), .A3(new_n693), .A4(new_n1004), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n682), .A2(new_n683), .A3(new_n696), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n994), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(new_n691), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n758), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1006), .A2(new_n1007), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n759), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n702), .B(KEYINPUT41), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n986), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n692), .A2(new_n998), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n715), .B1(new_n562), .B2(new_n678), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1017), .A2(new_n519), .A3(new_n679), .A4(new_n695), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(KEYINPUT42), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n988), .A2(new_n989), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n565), .B1(new_n1020), .B2(new_n514), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n686), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(KEYINPUT107), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1018), .A2(KEYINPUT42), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT107), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1019), .A2(new_n1022), .A3(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1024), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1016), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1028), .A2(new_n1016), .A3(new_n1029), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1032), .ZN(new_n1035));
  AND3_X1   g0835(.A1(new_n1028), .A2(new_n1016), .A3(new_n1029), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1035), .B1(new_n1036), .B2(new_n1030), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1034), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n984), .B1(new_n1015), .B2(new_n1038), .ZN(G387));
  NAND2_X1  g0839(.A1(new_n758), .A2(new_n1010), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(KEYINPUT112), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1010), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n759), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT112), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n758), .A2(new_n1010), .A3(new_n1044), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1041), .A2(new_n1043), .A3(new_n702), .A4(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n861), .B1(new_n685), .B2(new_n818), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n804), .A2(G159), .B1(new_n782), .B2(G68), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n798), .A2(G77), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n794), .A2(new_n307), .ZN(new_n1050));
  AND3_X1   g0850(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n785), .A2(G150), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n407), .B1(G50), .B2(new_n786), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n970), .A2(new_n264), .B1(new_n835), .B2(G97), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n970), .A2(G311), .B1(new_n804), .B2(G322), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1056), .B1(new_n791), .B2(new_n841), .C1(new_n965), .C2(new_n845), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT48), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n581), .B2(new_n770), .C1(new_n488), .C2(new_n792), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(KEYINPUT111), .B(KEYINPUT49), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1059), .B(new_n1060), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n407), .B1(new_n790), .B2(new_n583), .C1(new_n776), .C2(new_n784), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1055), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n767), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n264), .A2(new_n218), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT50), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n203), .A2(new_n208), .ZN(new_n1067));
  NOR4_X1   g0867(.A1(new_n1066), .A2(G45), .A3(new_n1067), .A4(new_n705), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n812), .B1(new_n240), .B2(new_n541), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n705), .A2(new_n232), .A3(new_n283), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1068), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n232), .A2(G107), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n819), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1047), .A2(new_n1064), .A3(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1042), .A2(KEYINPUT110), .A3(new_n986), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT110), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n1010), .B2(new_n985), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1046), .A2(new_n1074), .A3(new_n1078), .ZN(G393));
  NAND2_X1  g0879(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n703), .B1(new_n1080), .B2(new_n1043), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n1012), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1006), .A2(new_n986), .A3(new_n1007), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n990), .A2(new_n818), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n792), .A2(new_n581), .B1(new_n770), .B2(new_n583), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n283), .B(new_n1085), .C1(G294), .C2(new_n782), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n845), .A2(new_n838), .B1(new_n775), .B2(new_n965), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n1088));
  XNOR2_X1  g0888(.A(new_n1087), .B(new_n1088), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n779), .A2(new_n791), .B1(new_n790), .B2(new_n213), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G322), .B2(new_n785), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1086), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n804), .A2(G150), .B1(G159), .B2(new_n786), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT51), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n779), .A2(new_n218), .B1(new_n770), .B2(new_n208), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n407), .B1(new_n785), .B2(G143), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n798), .A2(G68), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1096), .A2(new_n840), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n841), .A2(new_n265), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1092), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n767), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n819), .B1(new_n357), .B2(new_n232), .C1(new_n956), .C2(new_n251), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1084), .A2(new_n764), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1082), .A2(new_n1083), .A3(new_n1104), .ZN(G390));
  OAI211_X1 g0905(.A(G330), .B(new_n906), .C1(new_n928), .C2(new_n929), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n913), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n721), .A2(new_n723), .A3(new_n855), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n853), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n756), .A2(G330), .A3(new_n906), .A4(new_n912), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1107), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n756), .A2(G330), .A3(new_n906), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n913), .ZN(new_n1113));
  OAI211_X1 g0913(.A(G330), .B(new_n924), .C1(new_n928), .C2(new_n929), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n916), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1111), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n942), .A2(G330), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n869), .A2(new_n1117), .A3(new_n653), .A4(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1108), .A2(new_n853), .A3(new_n912), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n898), .A2(new_n892), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1121), .A2(new_n872), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n871), .B1(new_n907), .B2(new_n913), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n895), .A2(new_n886), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n447), .B2(new_n885), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n901), .B1(new_n1126), .B2(new_n874), .ZN(new_n1127));
  OAI21_X1  g0927(.A(KEYINPUT39), .B1(new_n1127), .B2(new_n918), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1121), .A2(new_n901), .A3(new_n873), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1124), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1110), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n1123), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1114), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(new_n1123), .B2(new_n1130), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n702), .B1(new_n1119), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(KEYINPUT114), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1119), .A2(new_n1135), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT114), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1139), .B(new_n702), .C1(new_n1119), .C2(new_n1135), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1137), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1128), .A2(new_n1129), .A3(new_n816), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n798), .A2(G150), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT53), .ZN(new_n1144));
  INV_X1    g0944(.A(G128), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n775), .A2(new_n1145), .B1(new_n770), .B2(new_n806), .ZN(new_n1146));
  XOR2_X1   g0946(.A(KEYINPUT54), .B(G143), .Z(new_n1147));
  AND2_X1   g0947(.A1(new_n782), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(G125), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n283), .B1(new_n784), .B2(new_n1149), .C1(new_n829), .C2(new_n779), .ZN(new_n1150));
  NOR4_X1   g0950(.A1(new_n1144), .A2(new_n1146), .A3(new_n1148), .A4(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(G132), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1151), .B1(new_n218), .B2(new_n790), .C1(new_n1152), .C2(new_n845), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n836), .B1(new_n357), .B2(new_n841), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n283), .B(new_n1154), .C1(G107), .C2(new_n970), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n845), .A2(new_n583), .B1(new_n770), .B2(new_n208), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT115), .ZN(new_n1157));
  AND2_X1   g0957(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1158), .B1(new_n408), .B2(new_n792), .C1(new_n581), .C2(new_n775), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n784), .A2(new_n488), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1153), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n767), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1142), .A2(new_n764), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n265), .B2(new_n826), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1164), .B1(new_n1165), .B2(new_n986), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1141), .A2(new_n1166), .ZN(G378));
  AOI211_X1 g0967(.A(new_n866), .B(new_n448), .C1(new_n724), .C2(new_n727), .ZN(new_n1168));
  AOI21_X1  g0968(.A(KEYINPUT104), .B1(new_n864), .B2(new_n449), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n653), .B(new_n1118), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(KEYINPUT117), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT117), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n869), .A2(new_n1172), .A3(new_n653), .A4(new_n1118), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1171), .B(new_n1173), .C1(new_n1119), .C2(new_n1135), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n930), .A2(new_n931), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n938), .A2(new_n939), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1175), .A2(G330), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n652), .A2(new_n305), .ZN(new_n1178));
  XOR2_X1   g0978(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1179));
  OR2_X1    g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n282), .A2(new_n884), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1180), .A2(new_n282), .A3(new_n884), .A4(new_n1181), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1177), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n940), .A2(G330), .A3(new_n1186), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n920), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(KEYINPUT118), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n903), .A2(new_n904), .A3(new_n919), .ZN(new_n1192));
  AND4_X1   g0992(.A1(G330), .A2(new_n1186), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1186), .B1(new_n940), .B2(G330), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1192), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT118), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1188), .A2(new_n920), .A3(new_n1189), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1174), .A2(KEYINPUT57), .A3(new_n1191), .A4(new_n1198), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1188), .A2(new_n920), .A3(new_n1189), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1200), .A2(new_n1190), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n1111), .A2(new_n1116), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1170), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n1165), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1201), .B1(new_n1202), .B2(new_n1205), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1199), .B(new_n702), .C1(new_n1206), .C2(KEYINPUT57), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1187), .A2(new_n817), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n612), .A2(G33), .ZN(new_n1209));
  INV_X1    g1009(.A(G41), .ZN(new_n1210));
  AOI21_X1  g1010(.A(G50), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT116), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1212), .A2(G124), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(G124), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n785), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n770), .A2(new_n267), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n841), .A2(new_n829), .B1(new_n1145), .B2(new_n845), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(new_n798), .C2(new_n1147), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(new_n1149), .B2(new_n775), .C1(new_n1152), .C2(new_n779), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1210), .B(new_n1215), .C1(new_n1219), .C2(KEYINPUT59), .ZN(new_n1220));
  AOI211_X1 g1020(.A(G33), .B(new_n1220), .C1(G159), .C2(new_n835), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1219), .A2(KEYINPUT59), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1211), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(G41), .B1(new_n804), .B2(G116), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n782), .A2(new_n307), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1224), .A2(new_n407), .A3(new_n1049), .A4(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n835), .A2(G58), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1227), .B1(new_n203), .B2(new_n770), .C1(new_n581), .C2(new_n784), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1226), .B(new_n1228), .C1(G107), .C2(new_n786), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n357), .B2(new_n779), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT58), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n768), .B1(new_n1223), .B2(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n827), .A2(G50), .ZN(new_n1233));
  NOR4_X1   g1033(.A1(new_n1208), .A2(new_n861), .A3(new_n1232), .A4(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1234), .B1(new_n1235), .B2(new_n986), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1207), .A2(new_n1236), .ZN(G375));
  NAND2_X1  g1037(.A1(new_n1170), .A2(new_n1203), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1238), .A2(new_n1119), .A3(new_n1014), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n912), .A2(new_n817), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n827), .A2(G68), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n970), .A2(new_n1147), .B1(new_n804), .B2(G132), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(new_n829), .B2(new_n845), .ZN(new_n1243));
  XOR2_X1   g1043(.A(new_n1243), .B(KEYINPUT119), .Z(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G128), .B2(new_n785), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n794), .A2(G50), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1227), .A2(KEYINPUT120), .A3(new_n396), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n841), .A2(new_n267), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT120), .B1(new_n1227), .B2(new_n396), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n1248), .B(new_n1249), .C1(G159), .C2(new_n798), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .A4(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1050), .B1(new_n488), .B2(new_n775), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n841), .A2(new_n213), .B1(new_n790), .B2(new_n208), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n784), .A2(new_n791), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n320), .B1(new_n792), .B2(new_n357), .ZN(new_n1255));
  NOR4_X1   g1055(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n1256), .B1(new_n583), .B2(new_n779), .C1(new_n581), .C2(new_n845), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n768), .B1(new_n1251), .B2(new_n1257), .ZN(new_n1258));
  NOR4_X1   g1058(.A1(new_n1240), .A2(new_n861), .A3(new_n1241), .A4(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n1117), .B2(new_n986), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1239), .A2(new_n1260), .ZN(G381));
  XNOR2_X1  g1061(.A(G375), .B(KEYINPUT121), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1262), .A2(G378), .ZN(new_n1263));
  INV_X1    g1063(.A(G384), .ZN(new_n1264));
  INV_X1    g1064(.A(G387), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1046), .A2(new_n824), .A3(new_n1074), .A4(new_n1078), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(G381), .A2(G390), .A3(new_n1266), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1263), .A2(new_n1264), .A3(new_n1265), .A4(new_n1267), .ZN(G407));
  INV_X1    g1068(.A(G213), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(new_n1263), .B2(new_n677), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(G407), .ZN(G409));
  INV_X1    g1071(.A(new_n1014), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(new_n1012), .B2(new_n759), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1034), .B(new_n1037), .C1(new_n1273), .C2(new_n986), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(G390), .A2(new_n1274), .A3(new_n984), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(G393), .A2(G396), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1266), .ZN(new_n1277));
  NOR3_X1   g1077(.A1(new_n1275), .A2(new_n1277), .A3(KEYINPUT122), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1276), .A2(new_n1266), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n1082), .A2(new_n1083), .A3(new_n1104), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1279), .A2(G387), .A3(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(G390), .B1(new_n1274), .B2(new_n984), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1277), .A2(KEYINPUT122), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1281), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1278), .B1(new_n1284), .B2(new_n1275), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT62), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT60), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n702), .B(new_n1119), .C1(new_n1238), .C2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(KEYINPUT60), .B1(new_n1170), .B2(new_n1203), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1260), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1264), .ZN(new_n1291));
  OAI211_X1 g1091(.A(G384), .B(new_n1260), .C1(new_n1288), .C2(new_n1289), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1269), .A2(G343), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1207), .A2(G378), .A3(new_n1236), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1174), .A2(new_n1014), .A3(new_n1235), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1198), .A2(new_n986), .A3(new_n1191), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1166), .B(new_n1141), .C1(new_n1298), .C2(new_n1234), .ZN(new_n1299));
  AOI211_X1 g1099(.A(new_n1293), .B(new_n1294), .C1(new_n1295), .C2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT126), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1286), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1294), .B1(new_n1295), .B2(new_n1299), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1293), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1305), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1302), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT61), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1294), .A2(G2897), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1293), .A2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1291), .A2(new_n1292), .A3(new_n1309), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1308), .B1(new_n1303), .B2(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1285), .B1(new_n1307), .B2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(KEYINPUT63), .B1(new_n1303), .B2(new_n1313), .ZN(new_n1316));
  OAI21_X1  g1116(.A(KEYINPUT123), .B1(new_n1285), .B2(KEYINPUT61), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT123), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1275), .ZN(new_n1319));
  OAI22_X1  g1119(.A1(new_n1265), .A2(G390), .B1(KEYINPUT122), .B2(new_n1277), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1319), .B1(new_n1320), .B2(new_n1281), .ZN(new_n1321));
  OAI211_X1 g1121(.A(new_n1318), .B(new_n1308), .C1(new_n1321), .C2(new_n1278), .ZN(new_n1322));
  AOI22_X1  g1122(.A1(new_n1316), .A2(new_n1305), .B1(new_n1317), .B2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1295), .A2(new_n1299), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1294), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1324), .A2(KEYINPUT63), .A3(new_n1304), .A4(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT124), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1303), .A2(KEYINPUT124), .A3(KEYINPUT63), .A4(new_n1304), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT125), .ZN(new_n1331));
  AND3_X1   g1131(.A1(new_n1323), .A2(new_n1330), .A3(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1331), .B1(new_n1323), .B2(new_n1330), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1315), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(KEYINPUT127), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT127), .ZN(new_n1336));
  OAI211_X1 g1136(.A(new_n1315), .B(new_n1336), .C1(new_n1332), .C2(new_n1333), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1335), .A2(new_n1337), .ZN(G405));
  XNOR2_X1  g1138(.A(G375), .B(G378), .ZN(new_n1339));
  XNOR2_X1  g1139(.A(new_n1339), .B(new_n1293), .ZN(new_n1340));
  XNOR2_X1  g1140(.A(new_n1340), .B(new_n1285), .ZN(G402));
endmodule


