//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 1 0 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 1 0 1 0 0 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n822, new_n823, new_n824, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937;
  INV_X1    g000(.A(KEYINPUT97), .ZN(new_n202));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203));
  INV_X1    g002(.A(KEYINPUT15), .ZN(new_n204));
  OR2_X1    g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT14), .ZN(new_n206));
  INV_X1    g005(.A(G29gat), .ZN(new_n207));
  INV_X1    g006(.A(G36gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n210));
  AOI22_X1  g009(.A1(new_n209), .A2(new_n210), .B1(G29gat), .B2(G36gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n203), .A2(new_n204), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n205), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n210), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n215), .B1(KEYINPUT83), .B2(new_n209), .ZN(new_n216));
  OR2_X1    g015(.A1(new_n209), .A2(KEYINPUT83), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n216), .A2(new_n217), .B1(G29gat), .B2(G36gat), .ZN(new_n218));
  OR3_X1    g017(.A1(new_n218), .A2(KEYINPUT84), .A3(new_n205), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT84), .B1(new_n218), .B2(new_n205), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n214), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(KEYINPUT95), .A2(G85gat), .A3(G92gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT7), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g023(.A1(KEYINPUT95), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(G99gat), .A2(G106gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT8), .ZN(new_n227));
  INV_X1    g026(.A(G85gat), .ZN(new_n228));
  INV_X1    g027(.A(G92gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n224), .A2(new_n225), .A3(new_n227), .A4(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G99gat), .B(G106gat), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  AOI22_X1  g033(.A1(KEYINPUT8), .A2(new_n226), .B1(new_n228), .B2(new_n229), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n235), .A2(new_n232), .A3(new_n225), .A4(new_n224), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT41), .ZN(new_n238));
  NAND2_X1  g037(.A1(G232gat), .A2(G233gat), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n239), .B(KEYINPUT93), .Z(new_n240));
  OAI22_X1  g039(.A1(new_n221), .A2(new_n237), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n237), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n219), .A2(new_n220), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(new_n213), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT17), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n242), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n221), .A2(KEYINPUT17), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n241), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G190gat), .B(G218gat), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n202), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n240), .A2(new_n238), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n252), .B1(new_n244), .B2(new_n242), .ZN(new_n253));
  INV_X1    g052(.A(new_n247), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n237), .B1(new_n221), .B2(KEYINPUT17), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n256), .A2(KEYINPUT97), .A3(new_n249), .ZN(new_n257));
  AND2_X1   g056(.A1(new_n251), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n240), .A2(new_n238), .ZN(new_n259));
  XNOR2_X1  g058(.A(G134gat), .B(G162gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n261), .B1(new_n248), .B2(new_n250), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT96), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n248), .A2(new_n264), .A3(new_n250), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n253), .B(new_n250), .C1(new_n254), .C2(new_n255), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT96), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n251), .A2(new_n265), .A3(new_n267), .A4(new_n257), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT98), .ZN(new_n269));
  XOR2_X1   g068(.A(new_n261), .B(KEYINPUT94), .Z(new_n270));
  AND3_X1   g069(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n269), .B1(new_n268), .B2(new_n270), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n263), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G15gat), .B(G22gat), .ZN(new_n274));
  OR2_X1    g073(.A1(new_n274), .A2(G1gat), .ZN(new_n275));
  INV_X1    g074(.A(G1gat), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n276), .A2(KEYINPUT85), .A3(KEYINPUT16), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT85), .B1(new_n276), .B2(KEYINPUT16), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n274), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(G8gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n275), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT87), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n275), .A2(new_n279), .A3(KEYINPUT86), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n284), .B(G8gat), .C1(KEYINPUT86), .C2(new_n275), .ZN(new_n285));
  AND2_X1   g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT21), .ZN(new_n287));
  OR2_X1    g086(.A1(G57gat), .A2(G64gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT90), .ZN(new_n289));
  NAND2_X1  g088(.A1(G57gat), .A2(G64gat), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AND2_X1   g090(.A1(G57gat), .A2(G64gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(G57gat), .A2(G64gat), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT90), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n291), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT89), .B1(G71gat), .B2(G78gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(KEYINPUT89), .A2(G71gat), .A3(G78gat), .ZN(new_n300));
  INV_X1    g099(.A(G71gat), .ZN(new_n301));
  INV_X1    g100(.A(G78gat), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n299), .A2(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n301), .A2(new_n302), .A3(KEYINPUT9), .ZN(new_n305));
  NAND2_X1  g104(.A1(G71gat), .A2(G78gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n292), .A2(new_n293), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n286), .B1(new_n287), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n311), .B(KEYINPUT92), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n287), .ZN(new_n313));
  NAND2_X1  g112(.A1(G231gat), .A2(G233gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n313), .B(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(G127gat), .B(G155gat), .Z(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(KEYINPUT20), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n315), .B(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n312), .B(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(G183gat), .B(G211gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n321));
  XOR2_X1   g120(.A(new_n320), .B(new_n321), .Z(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  OR2_X1    g123(.A1(new_n312), .A2(new_n318), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n312), .A2(new_n318), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(new_n322), .A3(new_n326), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(G230gat), .A2(G233gat), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n300), .ZN(new_n331));
  OAI22_X1  g130(.A1(new_n331), .A2(new_n298), .B1(G71gat), .B2(G78gat), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n295), .B1(new_n308), .B2(new_n289), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n332), .B1(new_n333), .B2(new_n294), .ZN(new_n334));
  INV_X1    g133(.A(new_n309), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n237), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT10), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n304), .A2(new_n309), .A3(new_n236), .A4(new_n234), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT99), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n336), .A2(new_n338), .A3(KEYINPUT99), .A4(new_n337), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n338), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT10), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n330), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n329), .B1(new_n336), .B2(new_n338), .ZN(new_n347));
  XOR2_X1   g146(.A(G120gat), .B(G148gat), .Z(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(KEYINPUT100), .ZN(new_n349));
  XNOR2_X1  g148(.A(G176gat), .B(G204gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  OR3_X1    g151(.A1(new_n346), .A2(new_n347), .A3(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n352), .B1(new_n346), .B2(new_n347), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NOR3_X1   g154(.A1(new_n273), .A2(new_n328), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT88), .ZN(new_n357));
  XNOR2_X1  g156(.A(G8gat), .B(G36gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(G64gat), .B(G92gat), .ZN(new_n359));
  XOR2_X1   g158(.A(new_n358), .B(new_n359), .Z(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G197gat), .B(G204gat), .ZN(new_n362));
  INV_X1    g161(.A(G211gat), .ZN(new_n363));
  INV_X1    g162(.A(G218gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n362), .B1(KEYINPUT22), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G211gat), .B(G218gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT70), .ZN(new_n369));
  AND2_X1   g168(.A1(G183gat), .A2(G190gat), .ZN(new_n370));
  INV_X1    g169(.A(G169gat), .ZN(new_n371));
  INV_X1    g170(.A(G176gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NOR2_X1   g172(.A1(G169gat), .A2(G176gat), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n373), .A2(KEYINPUT26), .A3(new_n374), .ZN(new_n375));
  AOI211_X1 g174(.A(new_n370), .B(new_n375), .C1(KEYINPUT26), .C2(new_n374), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT27), .B(G183gat), .ZN(new_n377));
  INV_X1    g176(.A(G190gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT28), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(KEYINPUT66), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n373), .B1(KEYINPUT23), .B2(new_n374), .ZN(new_n384));
  OR2_X1    g183(.A1(new_n384), .A2(KEYINPUT65), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT24), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n386), .A2(G183gat), .A3(G190gat), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(new_n370), .B2(new_n386), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n388), .B1(G183gat), .B2(G190gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n374), .A2(KEYINPUT23), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT25), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n384), .A2(KEYINPUT65), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n385), .A2(new_n389), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n384), .B1(KEYINPUT23), .B2(new_n374), .ZN(new_n395));
  NOR2_X1   g194(.A1(G183gat), .A2(G190gat), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n396), .A2(KEYINPUT64), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(KEYINPUT64), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n388), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n391), .B1(new_n395), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n394), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n383), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT29), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(G226gat), .A2(G233gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n405), .B1(new_n401), .B2(new_n382), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n369), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n405), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n410), .B1(new_n402), .B2(new_n403), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n411), .A2(KEYINPUT70), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n368), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n401), .A2(new_n382), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n410), .A2(KEYINPUT29), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n416), .B1(new_n402), .B2(new_n405), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n418), .A2(new_n368), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n413), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n361), .B1(new_n421), .B2(KEYINPUT37), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n369), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT70), .B1(new_n411), .B2(new_n407), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n419), .B1(new_n425), .B2(new_n368), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT37), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT38), .B1(new_n422), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n360), .B1(new_n426), .B2(new_n427), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT38), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT78), .ZN(new_n432));
  INV_X1    g231(.A(new_n368), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n425), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n427), .B1(new_n417), .B2(new_n368), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n432), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n368), .B1(new_n423), .B2(new_n424), .ZN(new_n437));
  INV_X1    g236(.A(new_n435), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n437), .A2(KEYINPUT78), .A3(new_n438), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n430), .B(new_n431), .C1(new_n436), .C2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT71), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n441), .B1(new_n426), .B2(new_n360), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n433), .B1(new_n423), .B2(new_n424), .ZN(new_n443));
  NOR4_X1   g242(.A1(new_n443), .A2(KEYINPUT71), .A3(new_n361), .A4(new_n419), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(G1gat), .B(G29gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n446), .B(KEYINPUT0), .ZN(new_n447));
  XNOR2_X1  g246(.A(G57gat), .B(G85gat), .ZN(new_n448));
  XOR2_X1   g247(.A(new_n447), .B(new_n448), .Z(new_n449));
  XNOR2_X1  g248(.A(G155gat), .B(G162gat), .ZN(new_n450));
  XOR2_X1   g249(.A(G141gat), .B(G148gat), .Z(new_n451));
  AOI21_X1  g250(.A(new_n450), .B1(new_n451), .B2(KEYINPUT72), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT2), .ZN(new_n453));
  AND2_X1   g252(.A1(G155gat), .A2(G162gat), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  OAI221_X1 g255(.A(new_n451), .B1(new_n453), .B2(new_n454), .C1(new_n450), .C2(KEYINPUT72), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(KEYINPUT73), .ZN(new_n459));
  INV_X1    g258(.A(G127gat), .ZN(new_n460));
  OR3_X1    g259(.A1(new_n460), .A2(KEYINPUT67), .A3(G134gat), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT67), .B1(new_n460), .B2(G134gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(KEYINPUT68), .B(G127gat), .ZN(new_n463));
  INV_X1    g262(.A(G134gat), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n461), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(G113gat), .B(G120gat), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n465), .B1(KEYINPUT1), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT69), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(G120gat), .ZN(new_n470));
  OR3_X1    g269(.A1(new_n468), .A2(new_n470), .A3(G113gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n460), .A2(G134gat), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT1), .B1(new_n464), .B2(G127gat), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n469), .A2(new_n471), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n467), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n459), .A2(KEYINPUT4), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(G225gat), .A2(G233gat), .ZN(new_n478));
  INV_X1    g277(.A(new_n458), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(new_n475), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n476), .A2(new_n479), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT4), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n477), .A2(new_n478), .A3(new_n483), .A4(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT5), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n475), .B(new_n458), .ZN(new_n489));
  INV_X1    g288(.A(new_n478), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n488), .B1(new_n491), .B2(KEYINPUT74), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n487), .B(new_n492), .C1(KEYINPUT74), .C2(new_n491), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n459), .A2(new_n485), .A3(new_n476), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n484), .A2(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n496), .A2(new_n488), .A3(new_n478), .A4(new_n483), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n449), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT6), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT79), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n498), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT6), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n493), .A2(new_n449), .A3(new_n497), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n499), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT79), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n501), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n429), .A2(new_n440), .A3(new_n445), .A4(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n478), .B1(new_n496), .B2(new_n483), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT39), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT39), .B1(new_n489), .B2(new_n490), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n512), .B(new_n449), .C1(new_n510), .C2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT40), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n502), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n515), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT77), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n514), .A2(KEYINPUT77), .A3(new_n515), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n516), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR3_X1   g320(.A1(new_n442), .A2(new_n444), .A3(KEYINPUT30), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n413), .A2(KEYINPUT30), .A3(new_n360), .A4(new_n420), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n361), .B1(new_n443), .B2(new_n419), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n521), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n433), .B1(new_n481), .B2(new_n403), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n527), .B1(G228gat), .B2(G233gat), .ZN(new_n528));
  INV_X1    g327(.A(new_n459), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n480), .B1(new_n368), .B2(KEYINPUT29), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n530), .A2(new_n458), .ZN(new_n533));
  OAI211_X1 g332(.A(G228gat), .B(G233gat), .C1(new_n527), .C2(new_n533), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n532), .A2(G22gat), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(G22gat), .B1(new_n532), .B2(new_n534), .ZN(new_n536));
  XNOR2_X1  g335(.A(G78gat), .B(G106gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT31), .B(G50gat), .ZN(new_n538));
  XOR2_X1   g337(.A(new_n537), .B(new_n538), .Z(new_n539));
  XOR2_X1   g338(.A(new_n539), .B(KEYINPUT75), .Z(new_n540));
  OR3_X1    g339(.A1(new_n535), .A2(new_n536), .A3(new_n540), .ZN(new_n541));
  OAI22_X1  g340(.A1(new_n535), .A2(new_n536), .B1(KEYINPUT75), .B2(new_n539), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n509), .A2(new_n526), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n413), .A2(new_n360), .A3(new_n420), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT71), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT30), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n426), .A2(new_n441), .A3(new_n360), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n525), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n549), .A2(new_n506), .A3(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT76), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n543), .B(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT36), .ZN(new_n554));
  XOR2_X1   g353(.A(G15gat), .B(G43gat), .Z(new_n555));
  XNOR2_X1  g354(.A(G71gat), .B(G99gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n402), .A2(new_n476), .ZN(new_n559));
  AND2_X1   g358(.A1(G227gat), .A2(G233gat), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n383), .A2(new_n475), .A3(new_n401), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT33), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n558), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n560), .B1(new_n559), .B2(new_n561), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT34), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI211_X1 g366(.A(KEYINPUT34), .B(new_n560), .C1(new_n559), .C2(new_n561), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n564), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NOR3_X1   g369(.A1(new_n564), .A2(new_n567), .A3(new_n568), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n562), .A2(KEYINPUT32), .ZN(new_n572));
  NOR3_X1   g371(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n572), .ZN(new_n574));
  INV_X1    g373(.A(new_n567), .ZN(new_n575));
  INV_X1    g374(.A(new_n568), .ZN(new_n576));
  AND2_X1   g375(.A1(new_n562), .A2(new_n563), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n575), .B(new_n576), .C1(new_n577), .C2(new_n558), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n574), .B1(new_n578), .B2(new_n569), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n554), .B1(new_n573), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n572), .B1(new_n570), .B2(new_n571), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n578), .A2(new_n574), .A3(new_n569), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(new_n582), .A3(KEYINPUT36), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n551), .A2(new_n553), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n544), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n581), .A2(new_n582), .A3(new_n543), .ZN(new_n586));
  OAI21_X1  g385(.A(KEYINPUT35), .B1(new_n551), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n525), .B1(new_n445), .B2(new_n547), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT35), .ZN(new_n589));
  AND4_X1   g388(.A1(new_n589), .A2(new_n581), .A3(new_n582), .A4(new_n543), .ZN(new_n590));
  INV_X1    g389(.A(new_n508), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n585), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(KEYINPUT80), .B(KEYINPUT11), .Z(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT81), .ZN(new_n596));
  XOR2_X1   g395(.A(G113gat), .B(G141gat), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G169gat), .B(G197gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n244), .A2(new_n245), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n603), .A2(new_n286), .A3(new_n247), .ZN(new_n604));
  NAND2_X1  g403(.A1(G229gat), .A2(G233gat), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n286), .A2(new_n221), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT18), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n604), .A2(KEYINPUT18), .A3(new_n605), .A4(new_n606), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n286), .B(new_n221), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n605), .B(KEYINPUT13), .Z(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AND4_X1   g412(.A1(new_n602), .A2(new_n609), .A3(new_n610), .A4(new_n613), .ZN(new_n614));
  AOI22_X1  g413(.A1(new_n607), .A2(new_n608), .B1(new_n611), .B2(new_n612), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n602), .B1(new_n615), .B2(new_n610), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n357), .B1(new_n594), .B2(new_n618), .ZN(new_n619));
  AOI22_X1  g418(.A1(new_n544), .A2(new_n584), .B1(new_n587), .B2(new_n592), .ZN(new_n620));
  NOR3_X1   g419(.A1(new_n620), .A2(KEYINPUT88), .A3(new_n617), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n356), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT101), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n594), .A2(new_n357), .A3(new_n618), .ZN(new_n624));
  OAI21_X1  g423(.A(KEYINPUT88), .B1(new_n620), .B2(new_n617), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT101), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n626), .A2(new_n627), .A3(new_n356), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n506), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(G1gat), .ZN(G1324gat));
  INV_X1    g431(.A(new_n588), .ZN(new_n633));
  XOR2_X1   g432(.A(KEYINPUT16), .B(G8gat), .Z(new_n634));
  AOI21_X1  g433(.A(new_n627), .B1(new_n626), .B2(new_n356), .ZN(new_n635));
  INV_X1    g434(.A(new_n356), .ZN(new_n636));
  AOI211_X1 g435(.A(KEYINPUT101), .B(new_n636), .C1(new_n624), .C2(new_n625), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n633), .B(new_n634), .C1(new_n635), .C2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT42), .ZN(new_n639));
  OAI21_X1  g438(.A(KEYINPUT103), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n588), .B1(new_n623), .B2(new_n628), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT103), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n641), .A2(new_n642), .A3(KEYINPUT42), .A4(new_n634), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n635), .A2(new_n637), .ZN(new_n645));
  OAI21_X1  g444(.A(G8gat), .B1(new_n645), .B2(new_n588), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT102), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n638), .B2(new_n639), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n638), .A2(new_n647), .A3(new_n639), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n644), .B(new_n646), .C1(new_n648), .C2(new_n649), .ZN(G1325gat));
  NAND2_X1  g449(.A1(new_n580), .A2(new_n583), .ZN(new_n651));
  OAI21_X1  g450(.A(G15gat), .B1(new_n645), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n573), .A2(new_n579), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n654), .A2(G15gat), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n652), .B1(new_n645), .B2(new_n655), .ZN(G1326gat));
  XNOR2_X1  g455(.A(KEYINPUT43), .B(G22gat), .ZN(new_n657));
  INV_X1    g456(.A(new_n553), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n657), .B1(new_n645), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n660));
  INV_X1    g459(.A(new_n657), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n629), .A2(new_n553), .A3(new_n661), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n659), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n660), .B1(new_n659), .B2(new_n662), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(new_n664), .ZN(G1327gat));
  NAND2_X1  g464(.A1(new_n268), .A2(new_n270), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(KEYINPUT98), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n668));
  AOI22_X1  g467(.A1(new_n667), .A2(new_n668), .B1(new_n258), .B2(new_n262), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n620), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n670), .B(KEYINPUT44), .Z(new_n671));
  NAND2_X1  g470(.A1(new_n324), .A2(new_n327), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n672), .A2(new_n617), .A3(new_n355), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(G29gat), .B1(new_n674), .B2(new_n506), .ZN(new_n675));
  INV_X1    g474(.A(new_n355), .ZN(new_n676));
  AND4_X1   g475(.A1(new_n626), .A2(new_n328), .A3(new_n273), .A4(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n677), .A2(new_n207), .A3(new_n630), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n678), .A2(new_n680), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n675), .B1(new_n681), .B2(new_n682), .ZN(G1328gat));
  OAI21_X1  g482(.A(G36gat), .B1(new_n674), .B2(new_n588), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT46), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n677), .A2(new_n208), .A3(new_n633), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n677), .A2(new_n685), .A3(new_n208), .A4(new_n633), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT107), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  OAI221_X1 g489(.A(new_n684), .B1(new_n685), .B2(new_n686), .C1(new_n689), .C2(new_n690), .ZN(G1329gat));
  INV_X1    g490(.A(G43gat), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n674), .A2(new_n692), .A3(new_n651), .ZN(new_n693));
  AOI21_X1  g492(.A(G43gat), .B1(new_n677), .B2(new_n653), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  OR3_X1    g495(.A1(new_n693), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n696), .B1(new_n693), .B2(new_n694), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(G1330gat));
  OAI21_X1  g498(.A(G50gat), .B1(new_n674), .B2(new_n543), .ZN(new_n700));
  INV_X1    g499(.A(G50gat), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n677), .A2(new_n701), .A3(new_n553), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n700), .A2(KEYINPUT48), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(G50gat), .B1(new_n674), .B2(new_n658), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n704), .A2(new_n702), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n705), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g505(.A1(new_n669), .A2(new_n617), .A3(new_n672), .A4(new_n355), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n620), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n630), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g509(.A1(new_n620), .A2(new_n588), .A3(new_n707), .ZN(new_n711));
  NOR2_X1   g510(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n712));
  AND2_X1   g511(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n714), .B1(new_n711), .B2(new_n712), .ZN(G1333gat));
  INV_X1    g514(.A(new_n651), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n301), .B1(new_n708), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n654), .A2(G71gat), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n717), .B1(new_n708), .B2(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g519(.A1(new_n708), .A2(new_n553), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g521(.A1(new_n328), .A2(new_n617), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT109), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n724), .A2(new_n355), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n671), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(G85gat), .B1(new_n726), .B2(new_n506), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n670), .A2(new_n724), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n728), .B(KEYINPUT51), .Z(new_n729));
  AOI21_X1  g528(.A(new_n676), .B1(new_n729), .B2(KEYINPUT110), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(KEYINPUT110), .B2(new_n729), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n630), .A2(new_n228), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n727), .B1(new_n731), .B2(new_n732), .ZN(G1336gat));
  OAI21_X1  g532(.A(G92gat), .B1(new_n726), .B2(new_n588), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n729), .A2(new_n229), .A3(new_n633), .A4(new_n355), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT52), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT52), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n734), .A2(new_n735), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(G1337gat));
  OAI21_X1  g539(.A(G99gat), .B1(new_n726), .B2(new_n651), .ZN(new_n741));
  OR2_X1    g540(.A1(new_n654), .A2(G99gat), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n731), .B2(new_n742), .ZN(G1338gat));
  INV_X1    g542(.A(new_n543), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n671), .A2(new_n744), .A3(new_n725), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT53), .B1(new_n745), .B2(G106gat), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n543), .A2(G106gat), .A3(new_n676), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n729), .A2(KEYINPUT112), .A3(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT112), .B1(new_n729), .B2(new_n747), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n746), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(G106gat), .B1(new_n726), .B2(new_n658), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n747), .B(KEYINPUT111), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n729), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT53), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n751), .A2(new_n756), .ZN(G1339gat));
  NAND3_X1  g556(.A1(new_n356), .A2(KEYINPUT113), .A3(new_n617), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n669), .A2(new_n617), .A3(new_n672), .A4(new_n676), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT113), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT54), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n346), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n352), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n330), .B1(new_n338), .B2(new_n337), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n343), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n343), .A2(KEYINPUT114), .A3(new_n768), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT115), .ZN(new_n774));
  AOI22_X1  g573(.A1(new_n341), .A2(new_n342), .B1(KEYINPUT10), .B2(new_n344), .ZN(new_n775));
  OAI21_X1  g574(.A(KEYINPUT54), .B1(new_n775), .B2(new_n330), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n773), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT114), .B1(new_n343), .B2(new_n768), .ZN(new_n778));
  AOI211_X1 g577(.A(new_n770), .B(new_n767), .C1(new_n341), .C2(new_n342), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n346), .A2(new_n763), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT115), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n766), .B1(new_n777), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n353), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n774), .B1(new_n773), .B2(new_n776), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n780), .A2(new_n781), .A3(KEYINPUT115), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n765), .A2(new_n784), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n786), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n618), .A2(new_n785), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n615), .A2(new_n602), .A3(new_n610), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n605), .B1(new_n604), .B2(new_n606), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n611), .A2(new_n612), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n600), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(new_n676), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n273), .B1(new_n792), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n790), .B1(new_n777), .B2(new_n782), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n765), .B1(new_n787), .B2(new_n788), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n801), .B(new_n353), .C1(new_n802), .C2(KEYINPUT55), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n803), .A2(new_n797), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n273), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n328), .B1(new_n800), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n506), .B1(new_n762), .B2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n586), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n810), .A2(new_n633), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n617), .A2(G113gat), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT116), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n553), .B1(new_n762), .B2(new_n807), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n815), .A2(new_n630), .A3(new_n588), .A4(new_n653), .ZN(new_n816));
  OAI21_X1  g615(.A(G113gat), .B1(new_n816), .B2(new_n617), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n814), .A2(new_n817), .ZN(G1340gat));
  NOR3_X1   g617(.A1(new_n816), .A2(new_n470), .A3(new_n676), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n811), .A2(new_n355), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n820), .B2(new_n470), .ZN(G1341gat));
  INV_X1    g620(.A(new_n463), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n811), .A2(new_n822), .A3(new_n672), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n463), .B1(new_n816), .B2(new_n328), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(G1342gat));
  NAND2_X1  g624(.A1(new_n588), .A2(new_n273), .ZN(new_n826));
  OR3_X1    g625(.A1(new_n810), .A2(G134gat), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT56), .ZN(new_n828));
  XOR2_X1   g627(.A(new_n828), .B(KEYINPUT117), .Z(new_n829));
  OAI21_X1  g628(.A(G134gat), .B1(new_n816), .B2(new_n669), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n829), .B(new_n830), .C1(KEYINPUT56), .C2(new_n827), .ZN(G1343gat));
  NAND2_X1  g630(.A1(new_n588), .A2(new_n630), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n716), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n762), .A2(new_n807), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT57), .B1(new_n834), .B2(new_n744), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n617), .B1(new_n803), .B2(KEYINPUT119), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT119), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n785), .A2(new_n791), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n798), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n805), .B1(new_n840), .B2(new_n273), .ZN(new_n841));
  AOI22_X1  g640(.A1(new_n841), .A2(new_n328), .B1(new_n761), .B2(new_n758), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n553), .A2(KEYINPUT57), .ZN(new_n843));
  OAI22_X1  g642(.A1(new_n835), .A2(new_n836), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n835), .A2(new_n836), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n833), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(G141gat), .B1(new_n846), .B2(new_n617), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n808), .A2(new_n744), .A3(new_n651), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(new_n633), .ZN(new_n849));
  INV_X1    g648(.A(G141gat), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n849), .A2(new_n850), .A3(new_n618), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g652(.A(G148gat), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(KEYINPUT59), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n855), .B1(new_n846), .B2(new_n676), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n801), .A2(new_n353), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT55), .B1(new_n789), .B2(new_n766), .ZN(new_n859));
  OAI21_X1  g658(.A(KEYINPUT119), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n618), .A3(new_n839), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n273), .B1(new_n861), .B2(new_n799), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n857), .B1(new_n862), .B2(new_n806), .ZN(new_n863));
  OAI211_X1 g662(.A(KEYINPUT120), .B(new_n805), .C1(new_n840), .C2(new_n273), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(new_n328), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n658), .B1(new_n865), .B2(new_n759), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT121), .B1(new_n866), .B2(KEYINPUT57), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT121), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n869));
  INV_X1    g668(.A(new_n759), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n672), .B1(new_n841), .B2(new_n857), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n864), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n868), .B(new_n869), .C1(new_n872), .C2(new_n658), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n834), .A2(KEYINPUT57), .A3(new_n744), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n867), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n716), .A2(new_n832), .A3(new_n676), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n854), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n856), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n849), .A2(new_n854), .A3(new_n355), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT122), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n879), .A2(KEYINPUT122), .A3(new_n880), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(G1345gat));
  OAI21_X1  g684(.A(G155gat), .B1(new_n846), .B2(new_n328), .ZN(new_n886));
  INV_X1    g685(.A(G155gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n849), .A2(new_n887), .A3(new_n672), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n888), .ZN(G1346gat));
  OAI21_X1  g688(.A(G162gat), .B1(new_n846), .B2(new_n669), .ZN(new_n890));
  OR2_X1    g689(.A1(new_n826), .A2(G162gat), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n890), .B1(new_n848), .B2(new_n891), .ZN(G1347gat));
  NAND4_X1  g691(.A1(new_n815), .A2(new_n506), .A3(new_n633), .A4(new_n653), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT124), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n894), .A2(new_n371), .A3(new_n617), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n834), .A2(new_n506), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT123), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n897), .A2(new_n633), .A3(new_n809), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n618), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n895), .B1(new_n899), .B2(new_n371), .ZN(G1348gat));
  NAND3_X1  g699(.A1(new_n898), .A2(new_n372), .A3(new_n355), .ZN(new_n901));
  OAI21_X1  g700(.A(G176gat), .B1(new_n894), .B2(new_n676), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT125), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n903), .B(new_n904), .ZN(G1349gat));
  NAND3_X1  g704(.A1(new_n898), .A2(new_n377), .A3(new_n672), .ZN(new_n906));
  OAI21_X1  g705(.A(G183gat), .B1(new_n894), .B2(new_n328), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g708(.A1(new_n898), .A2(new_n378), .A3(new_n273), .ZN(new_n910));
  OAI21_X1  g709(.A(G190gat), .B1(new_n894), .B2(new_n669), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n911), .A2(KEYINPUT61), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n911), .A2(KEYINPUT61), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(G1351gat));
  AND4_X1   g713(.A1(new_n633), .A2(new_n897), .A3(new_n744), .A4(new_n651), .ZN(new_n915));
  INV_X1    g714(.A(G197gat), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n915), .A2(new_n916), .A3(new_n618), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n716), .A2(new_n630), .A3(new_n588), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n875), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(KEYINPUT126), .B1(new_n919), .B2(new_n617), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(G197gat), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n919), .A2(KEYINPUT126), .A3(new_n617), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n917), .B1(new_n921), .B2(new_n922), .ZN(G1352gat));
  INV_X1    g722(.A(G204gat), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n915), .A2(new_n924), .A3(new_n355), .ZN(new_n925));
  AND2_X1   g724(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n926));
  NOR2_X1   g725(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(G204gat), .B1(new_n919), .B2(new_n676), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n928), .B(new_n929), .C1(new_n926), .C2(new_n925), .ZN(G1353gat));
  NAND3_X1  g729(.A1(new_n915), .A2(new_n363), .A3(new_n672), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n875), .A2(new_n672), .A3(new_n918), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n932), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n933));
  AOI21_X1  g732(.A(KEYINPUT63), .B1(new_n932), .B2(G211gat), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(G1354gat));
  OAI21_X1  g734(.A(G218gat), .B1(new_n919), .B2(new_n669), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n915), .A2(new_n364), .A3(new_n273), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1355gat));
endmodule


