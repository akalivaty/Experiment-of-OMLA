

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581;

  AND2_X1 U321 ( .A1(n466), .A2(n444), .ZN(n445) );
  AND2_X1 U322 ( .A1(n565), .A2(n532), .ZN(n362) );
  XNOR2_X1 U323 ( .A(n450), .B(n449), .ZN(n526) );
  XOR2_X1 U324 ( .A(n321), .B(n435), .Z(n289) );
  AND2_X1 U325 ( .A1(G230GAT), .A2(G233GAT), .ZN(n290) );
  INV_X1 U326 ( .A(n573), .ZN(n400) );
  NAND2_X1 U327 ( .A1(n472), .A2(n400), .ZN(n401) );
  OR2_X1 U328 ( .A1(n402), .A2(n401), .ZN(n403) );
  XOR2_X1 U329 ( .A(G120GAT), .B(G71GAT), .Z(n345) );
  XNOR2_X1 U330 ( .A(n350), .B(n290), .ZN(n351) );
  INV_X1 U331 ( .A(n544), .ZN(n444) );
  XNOR2_X1 U332 ( .A(n352), .B(n351), .ZN(n355) );
  NAND2_X1 U333 ( .A1(n549), .A2(n546), .ZN(n458) );
  NOR2_X1 U334 ( .A1(n471), .A2(n470), .ZN(n485) );
  XOR2_X1 U335 ( .A(n569), .B(KEYINPUT41), .Z(n532) );
  INV_X1 U336 ( .A(n414), .ZN(n326) );
  INV_X1 U337 ( .A(G134GAT), .ZN(n451) );
  NOR2_X1 U338 ( .A1(n518), .A2(n497), .ZN(n498) );
  XNOR2_X1 U339 ( .A(n490), .B(n489), .ZN(n497) );
  XNOR2_X1 U340 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U341 ( .A(n454), .B(n453), .ZN(G1343GAT) );
  INV_X1 U342 ( .A(KEYINPUT117), .ZN(n450) );
  XOR2_X1 U343 ( .A(KEYINPUT21), .B(G218GAT), .Z(n292) );
  XNOR2_X1 U344 ( .A(KEYINPUT89), .B(G211GAT), .ZN(n291) );
  XNOR2_X1 U345 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U346 ( .A(G197GAT), .B(n293), .Z(n422) );
  XOR2_X1 U347 ( .A(G155GAT), .B(KEYINPUT2), .Z(n295) );
  XNOR2_X1 U348 ( .A(G162GAT), .B(KEYINPUT3), .ZN(n294) );
  XNOR2_X1 U349 ( .A(n295), .B(n294), .ZN(n438) );
  XOR2_X1 U350 ( .A(n438), .B(KEYINPUT23), .Z(n297) );
  NAND2_X1 U351 ( .A1(G228GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U352 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U353 ( .A(n422), .B(n298), .ZN(n310) );
  XOR2_X1 U354 ( .A(KEYINPUT92), .B(KEYINPUT90), .Z(n300) );
  XNOR2_X1 U355 ( .A(G204GAT), .B(KEYINPUT22), .ZN(n299) );
  XNOR2_X1 U356 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U357 ( .A(KEYINPUT24), .B(KEYINPUT87), .Z(n302) );
  XNOR2_X1 U358 ( .A(KEYINPUT88), .B(KEYINPUT91), .ZN(n301) );
  XNOR2_X1 U359 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U360 ( .A(n304), .B(n303), .Z(n308) );
  XNOR2_X1 U361 ( .A(G50GAT), .B(G22GAT), .ZN(n305) );
  XNOR2_X1 U362 ( .A(n305), .B(G141GAT), .ZN(n342) );
  XNOR2_X1 U363 ( .A(G106GAT), .B(G78GAT), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n306), .B(G148GAT), .ZN(n359) );
  XNOR2_X1 U365 ( .A(n342), .B(n359), .ZN(n307) );
  XNOR2_X1 U366 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U367 ( .A(n310), .B(n309), .ZN(n546) );
  XOR2_X1 U368 ( .A(n546), .B(KEYINPUT28), .Z(n518) );
  XOR2_X1 U369 ( .A(G176GAT), .B(KEYINPUT84), .Z(n312) );
  XNOR2_X1 U370 ( .A(KEYINPUT20), .B(KEYINPUT86), .ZN(n311) );
  XNOR2_X1 U371 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U372 ( .A(G99GAT), .B(n345), .Z(n314) );
  XOR2_X1 U373 ( .A(G190GAT), .B(G134GAT), .Z(n364) );
  XNOR2_X1 U374 ( .A(G43GAT), .B(n364), .ZN(n313) );
  XNOR2_X1 U375 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U376 ( .A(n316), .B(n315), .Z(n318) );
  NAND2_X1 U377 ( .A1(G227GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U378 ( .A(n318), .B(n317), .ZN(n321) );
  XOR2_X1 U379 ( .A(G127GAT), .B(KEYINPUT0), .Z(n320) );
  XNOR2_X1 U380 ( .A(G113GAT), .B(KEYINPUT83), .ZN(n319) );
  XNOR2_X1 U381 ( .A(n320), .B(n319), .ZN(n435) );
  XNOR2_X1 U382 ( .A(G169GAT), .B(G15GAT), .ZN(n322) );
  XNOR2_X1 U383 ( .A(n289), .B(n322), .ZN(n327) );
  XOR2_X1 U384 ( .A(KEYINPUT85), .B(KEYINPUT17), .Z(n324) );
  XNOR2_X1 U385 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n323) );
  XNOR2_X1 U386 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U387 ( .A(KEYINPUT19), .B(n325), .Z(n414) );
  XNOR2_X2 U388 ( .A(n327), .B(n326), .ZN(n549) );
  XOR2_X1 U389 ( .A(G197GAT), .B(G113GAT), .Z(n330) );
  XNOR2_X1 U390 ( .A(G169GAT), .B(G36GAT), .ZN(n328) );
  XNOR2_X1 U391 ( .A(n328), .B(G8GAT), .ZN(n416) );
  XNOR2_X1 U392 ( .A(KEYINPUT66), .B(n416), .ZN(n329) );
  XNOR2_X1 U393 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U394 ( .A(n331), .B(KEYINPUT65), .Z(n336) );
  XOR2_X1 U395 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n333) );
  NAND2_X1 U396 ( .A1(G229GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U397 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U398 ( .A(KEYINPUT69), .B(n334), .ZN(n335) );
  XNOR2_X1 U399 ( .A(n336), .B(n335), .ZN(n338) );
  XNOR2_X1 U400 ( .A(G15GAT), .B(G1GAT), .ZN(n337) );
  XNOR2_X1 U401 ( .A(n337), .B(KEYINPUT68), .ZN(n391) );
  XOR2_X1 U402 ( .A(n338), .B(n391), .Z(n344) );
  XOR2_X1 U403 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n340) );
  XNOR2_X1 U404 ( .A(G43GAT), .B(G29GAT), .ZN(n339) );
  XNOR2_X1 U405 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U406 ( .A(KEYINPUT67), .B(n341), .Z(n377) );
  XNOR2_X1 U407 ( .A(n377), .B(n342), .ZN(n343) );
  XNOR2_X1 U408 ( .A(n344), .B(n343), .ZN(n565) );
  XOR2_X1 U409 ( .A(KEYINPUT74), .B(KEYINPUT76), .Z(n347) );
  XOR2_X1 U410 ( .A(G99GAT), .B(G85GAT), .Z(n363) );
  XNOR2_X1 U411 ( .A(n345), .B(n363), .ZN(n346) );
  XNOR2_X1 U412 ( .A(n347), .B(n346), .ZN(n352) );
  XOR2_X1 U413 ( .A(KEYINPUT32), .B(KEYINPUT73), .Z(n349) );
  XNOR2_X1 U414 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n348) );
  XNOR2_X1 U415 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U416 ( .A(KEYINPUT13), .B(KEYINPUT71), .Z(n354) );
  XNOR2_X1 U417 ( .A(G57GAT), .B(KEYINPUT72), .ZN(n353) );
  XNOR2_X1 U418 ( .A(n354), .B(n353), .ZN(n395) );
  XOR2_X1 U419 ( .A(n355), .B(n395), .Z(n361) );
  XOR2_X1 U420 ( .A(G92GAT), .B(G64GAT), .Z(n357) );
  XNOR2_X1 U421 ( .A(G176GAT), .B(KEYINPUT75), .ZN(n356) );
  XNOR2_X1 U422 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U423 ( .A(G204GAT), .B(n358), .Z(n415) );
  XNOR2_X1 U424 ( .A(n359), .B(n415), .ZN(n360) );
  XNOR2_X1 U425 ( .A(n361), .B(n360), .ZN(n569) );
  XNOR2_X1 U426 ( .A(KEYINPUT46), .B(n362), .ZN(n402) );
  XOR2_X1 U427 ( .A(n363), .B(G106GAT), .Z(n366) );
  XNOR2_X1 U428 ( .A(n364), .B(G218GAT), .ZN(n365) );
  XNOR2_X1 U429 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U430 ( .A(KEYINPUT77), .B(KEYINPUT11), .Z(n368) );
  XNOR2_X1 U431 ( .A(G36GAT), .B(G162GAT), .ZN(n367) );
  XNOR2_X1 U432 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U433 ( .A(n370), .B(n369), .Z(n372) );
  XNOR2_X1 U434 ( .A(G50GAT), .B(G92GAT), .ZN(n371) );
  XNOR2_X1 U435 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U436 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n374) );
  NAND2_X1 U437 ( .A1(G232GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U438 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U439 ( .A(n376), .B(n375), .Z(n379) );
  XNOR2_X1 U440 ( .A(n377), .B(KEYINPUT78), .ZN(n378) );
  XOR2_X1 U441 ( .A(n379), .B(n378), .Z(n559) );
  INV_X1 U442 ( .A(n559), .ZN(n472) );
  XOR2_X1 U443 ( .A(KEYINPUT79), .B(KEYINPUT12), .Z(n381) );
  XNOR2_X1 U444 ( .A(KEYINPUT81), .B(KEYINPUT82), .ZN(n380) );
  XNOR2_X1 U445 ( .A(n381), .B(n380), .ZN(n399) );
  XOR2_X1 U446 ( .A(G155GAT), .B(G211GAT), .Z(n383) );
  XNOR2_X1 U447 ( .A(G22GAT), .B(G183GAT), .ZN(n382) );
  XNOR2_X1 U448 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U449 ( .A(KEYINPUT80), .B(G64GAT), .Z(n385) );
  XNOR2_X1 U450 ( .A(G8GAT), .B(G78GAT), .ZN(n384) );
  XNOR2_X1 U451 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U452 ( .A(n387), .B(n386), .Z(n393) );
  XOR2_X1 U453 ( .A(G71GAT), .B(G127GAT), .Z(n389) );
  NAND2_X1 U454 ( .A1(G231GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U455 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U456 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U457 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U458 ( .A(n394), .B(KEYINPUT15), .Z(n397) );
  XNOR2_X1 U459 ( .A(n395), .B(KEYINPUT14), .ZN(n396) );
  XNOR2_X1 U460 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U461 ( .A(n399), .B(n398), .Z(n573) );
  XNOR2_X1 U462 ( .A(KEYINPUT47), .B(n403), .ZN(n409) );
  XOR2_X1 U463 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n405) );
  XNOR2_X1 U464 ( .A(KEYINPUT36), .B(n559), .ZN(n576) );
  NAND2_X1 U465 ( .A1(n573), .A2(n576), .ZN(n404) );
  XNOR2_X1 U466 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U467 ( .A(n565), .B(KEYINPUT70), .ZN(n550) );
  INV_X1 U468 ( .A(n550), .ZN(n457) );
  NAND2_X1 U469 ( .A1(n406), .A2(n457), .ZN(n407) );
  NOR2_X1 U470 ( .A1(n569), .A2(n407), .ZN(n408) );
  NOR2_X1 U471 ( .A1(n409), .A2(n408), .ZN(n410) );
  XNOR2_X1 U472 ( .A(KEYINPUT48), .B(n410), .ZN(n542) );
  INV_X1 U473 ( .A(n542), .ZN(n446) );
  XOR2_X1 U474 ( .A(G190GAT), .B(KEYINPUT97), .Z(n412) );
  NAND2_X1 U475 ( .A1(G226GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U476 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U477 ( .A(n414), .B(n413), .ZN(n420) );
  XOR2_X1 U478 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n418) );
  XNOR2_X1 U479 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U481 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U482 ( .A(n422), .B(n421), .ZN(n541) );
  XOR2_X1 U483 ( .A(KEYINPUT27), .B(KEYINPUT100), .Z(n423) );
  XNOR2_X1 U484 ( .A(n541), .B(n423), .ZN(n466) );
  XOR2_X1 U485 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n425) );
  XNOR2_X1 U486 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n424) );
  XNOR2_X1 U487 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U488 ( .A(KEYINPUT95), .B(KEYINPUT5), .Z(n427) );
  XNOR2_X1 U489 ( .A(G57GAT), .B(KEYINPUT96), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U492 ( .A(G148GAT), .B(G120GAT), .Z(n431) );
  XNOR2_X1 U493 ( .A(G29GAT), .B(G141GAT), .ZN(n430) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U495 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U496 ( .A(n434), .B(KEYINPUT93), .Z(n437) );
  XNOR2_X1 U497 ( .A(n435), .B(KEYINPUT94), .ZN(n436) );
  XNOR2_X1 U498 ( .A(n437), .B(n436), .ZN(n443) );
  XOR2_X1 U499 ( .A(G85GAT), .B(n438), .Z(n440) );
  NAND2_X1 U500 ( .A1(G225GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U501 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U502 ( .A(G134GAT), .B(n441), .Z(n442) );
  XNOR2_X1 U503 ( .A(n443), .B(n442), .ZN(n544) );
  NAND2_X1 U504 ( .A1(n446), .A2(n445), .ZN(n447) );
  XNOR2_X1 U505 ( .A(KEYINPUT116), .B(n447), .ZN(n530) );
  NOR2_X1 U506 ( .A1(n549), .A2(n530), .ZN(n448) );
  AND2_X1 U507 ( .A1(n518), .A2(n448), .ZN(n449) );
  NAND2_X1 U508 ( .A1(n526), .A2(n559), .ZN(n454) );
  XOR2_X1 U509 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n452) );
  XOR2_X1 U510 ( .A(KEYINPUT104), .B(KEYINPUT103), .Z(n456) );
  XNOR2_X1 U511 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n455) );
  XNOR2_X1 U512 ( .A(n456), .B(n455), .ZN(n476) );
  NOR2_X1 U513 ( .A1(n457), .A2(n569), .ZN(n488) );
  XOR2_X1 U514 ( .A(KEYINPUT101), .B(KEYINPUT26), .Z(n459) );
  XOR2_X1 U515 ( .A(n459), .B(n458), .Z(n529) );
  NAND2_X1 U516 ( .A1(n529), .A2(n466), .ZN(n460) );
  XNOR2_X1 U517 ( .A(n460), .B(KEYINPUT102), .ZN(n461) );
  NAND2_X1 U518 ( .A1(n461), .A2(n544), .ZN(n465) );
  NOR2_X1 U519 ( .A1(n549), .A2(n541), .ZN(n462) );
  NOR2_X1 U520 ( .A1(n546), .A2(n462), .ZN(n463) );
  XOR2_X1 U521 ( .A(KEYINPUT25), .B(n463), .Z(n464) );
  NOR2_X1 U522 ( .A1(n465), .A2(n464), .ZN(n471) );
  NAND2_X1 U523 ( .A1(n466), .A2(n518), .ZN(n468) );
  INV_X1 U524 ( .A(n549), .ZN(n467) );
  NOR2_X1 U525 ( .A1(n468), .A2(n467), .ZN(n469) );
  NOR2_X1 U526 ( .A1(n544), .A2(n469), .ZN(n470) );
  NAND2_X1 U527 ( .A1(n472), .A2(n573), .ZN(n473) );
  XOR2_X1 U528 ( .A(KEYINPUT16), .B(n473), .Z(n474) );
  AND2_X1 U529 ( .A1(n485), .A2(n474), .ZN(n500) );
  NAND2_X1 U530 ( .A1(n488), .A2(n500), .ZN(n482) );
  NOR2_X1 U531 ( .A1(n544), .A2(n482), .ZN(n475) );
  XOR2_X1 U532 ( .A(n476), .B(n475), .Z(G1324GAT) );
  NOR2_X1 U533 ( .A1(n541), .A2(n482), .ZN(n477) );
  XOR2_X1 U534 ( .A(G8GAT), .B(n477), .Z(G1325GAT) );
  NOR2_X1 U535 ( .A1(n482), .A2(n549), .ZN(n481) );
  XOR2_X1 U536 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n479) );
  XNOR2_X1 U537 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n481), .B(n480), .ZN(G1326GAT) );
  NOR2_X1 U540 ( .A1(n518), .A2(n482), .ZN(n484) );
  XNOR2_X1 U541 ( .A(G22GAT), .B(KEYINPUT107), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n484), .B(n483), .ZN(G1327GAT) );
  XNOR2_X1 U543 ( .A(KEYINPUT108), .B(KEYINPUT38), .ZN(n490) );
  NAND2_X1 U544 ( .A1(n576), .A2(n485), .ZN(n486) );
  NOR2_X1 U545 ( .A1(n573), .A2(n486), .ZN(n487) );
  XOR2_X1 U546 ( .A(KEYINPUT37), .B(n487), .Z(n511) );
  NAND2_X1 U547 ( .A1(n511), .A2(n488), .ZN(n489) );
  NOR2_X1 U548 ( .A1(n544), .A2(n497), .ZN(n492) );
  XNOR2_X1 U549 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n492), .B(n491), .ZN(G1328GAT) );
  NOR2_X1 U551 ( .A1(n541), .A2(n497), .ZN(n493) );
  XOR2_X1 U552 ( .A(G36GAT), .B(n493), .Z(G1329GAT) );
  NOR2_X1 U553 ( .A1(n549), .A2(n497), .ZN(n495) );
  XNOR2_X1 U554 ( .A(KEYINPUT40), .B(KEYINPUT109), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(n496), .ZN(G1330GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT110), .B(n498), .Z(n499) );
  XNOR2_X1 U558 ( .A(G50GAT), .B(n499), .ZN(G1331GAT) );
  XNOR2_X1 U559 ( .A(n532), .B(KEYINPUT111), .ZN(n523) );
  NOR2_X1 U560 ( .A1(n523), .A2(n565), .ZN(n510) );
  AND2_X1 U561 ( .A1(n510), .A2(n500), .ZN(n501) );
  XOR2_X1 U562 ( .A(KEYINPUT112), .B(n501), .Z(n506) );
  NOR2_X1 U563 ( .A1(n506), .A2(n544), .ZN(n502) );
  XOR2_X1 U564 ( .A(n502), .B(KEYINPUT42), .Z(n503) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(n503), .ZN(G1332GAT) );
  NOR2_X1 U566 ( .A1(n506), .A2(n541), .ZN(n504) );
  XOR2_X1 U567 ( .A(G64GAT), .B(n504), .Z(G1333GAT) );
  NOR2_X1 U568 ( .A1(n549), .A2(n506), .ZN(n505) );
  XOR2_X1 U569 ( .A(G71GAT), .B(n505), .Z(G1334GAT) );
  XNOR2_X1 U570 ( .A(KEYINPUT113), .B(KEYINPUT43), .ZN(n508) );
  NOR2_X1 U571 ( .A1(n518), .A2(n506), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U573 ( .A(G78GAT), .B(n509), .Z(G1335GAT) );
  NAND2_X1 U574 ( .A1(n511), .A2(n510), .ZN(n517) );
  NOR2_X1 U575 ( .A1(n544), .A2(n517), .ZN(n512) );
  XOR2_X1 U576 ( .A(n512), .B(KEYINPUT114), .Z(n513) );
  XNOR2_X1 U577 ( .A(G85GAT), .B(n513), .ZN(G1336GAT) );
  NOR2_X1 U578 ( .A1(n541), .A2(n517), .ZN(n515) );
  XNOR2_X1 U579 ( .A(G92GAT), .B(KEYINPUT115), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(G1337GAT) );
  NOR2_X1 U581 ( .A1(n549), .A2(n517), .ZN(n516) );
  XOR2_X1 U582 ( .A(G99GAT), .B(n516), .Z(G1338GAT) );
  NOR2_X1 U583 ( .A1(n518), .A2(n517), .ZN(n519) );
  XOR2_X1 U584 ( .A(KEYINPUT44), .B(n519), .Z(n520) );
  XNOR2_X1 U585 ( .A(G106GAT), .B(n520), .ZN(G1339GAT) );
  NAND2_X1 U586 ( .A1(n550), .A2(n526), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n521), .B(KEYINPUT118), .ZN(n522) );
  XNOR2_X1 U588 ( .A(G113GAT), .B(n522), .ZN(G1340GAT) );
  XOR2_X1 U589 ( .A(G120GAT), .B(KEYINPUT49), .Z(n525) );
  INV_X1 U590 ( .A(n523), .ZN(n553) );
  NAND2_X1 U591 ( .A1(n526), .A2(n553), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(G1341GAT) );
  NAND2_X1 U593 ( .A1(n526), .A2(n573), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n527), .B(KEYINPUT50), .ZN(n528) );
  XNOR2_X1 U595 ( .A(G127GAT), .B(n528), .ZN(G1342GAT) );
  INV_X1 U596 ( .A(n529), .ZN(n564) );
  NOR2_X1 U597 ( .A1(n530), .A2(n564), .ZN(n538) );
  NAND2_X1 U598 ( .A1(n565), .A2(n538), .ZN(n531) );
  XNOR2_X1 U599 ( .A(G141GAT), .B(n531), .ZN(G1344GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n534) );
  NAND2_X1 U601 ( .A1(n538), .A2(n532), .ZN(n533) );
  XNOR2_X1 U602 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U603 ( .A(G148GAT), .B(n535), .ZN(G1345GAT) );
  NAND2_X1 U604 ( .A1(n538), .A2(n573), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n536), .B(KEYINPUT120), .ZN(n537) );
  XNOR2_X1 U606 ( .A(G155GAT), .B(n537), .ZN(G1346GAT) );
  XOR2_X1 U607 ( .A(G162GAT), .B(KEYINPUT121), .Z(n540) );
  NAND2_X1 U608 ( .A1(n538), .A2(n559), .ZN(n539) );
  XNOR2_X1 U609 ( .A(n540), .B(n539), .ZN(G1347GAT) );
  NOR2_X1 U610 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n543), .B(KEYINPUT54), .ZN(n545) );
  NAND2_X1 U612 ( .A1(n545), .A2(n544), .ZN(n563) );
  NOR2_X1 U613 ( .A1(n546), .A2(n563), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n547), .B(KEYINPUT55), .ZN(n548) );
  NOR2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n560) );
  NAND2_X1 U616 ( .A1(n550), .A2(n560), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n551), .B(KEYINPUT122), .ZN(n552) );
  XNOR2_X1 U618 ( .A(G169GAT), .B(n552), .ZN(G1348GAT) );
  XOR2_X1 U619 ( .A(G176GAT), .B(KEYINPUT123), .Z(n555) );
  NAND2_X1 U620 ( .A1(n553), .A2(n560), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(n557) );
  XOR2_X1 U622 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1349GAT) );
  NAND2_X1 U624 ( .A1(n560), .A2(n573), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U626 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n562) );
  NAND2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1351GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n567) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n577) );
  NAND2_X1 U631 ( .A1(n577), .A2(n565), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n571) );
  NAND2_X1 U635 ( .A1(n577), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G204GAT), .B(n572), .ZN(G1353GAT) );
  XOR2_X1 U638 ( .A(G211GAT), .B(KEYINPUT125), .Z(n575) );
  NAND2_X1 U639 ( .A1(n577), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1354GAT) );
  XNOR2_X1 U641 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n581) );
  XOR2_X1 U642 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n579) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(G1355GAT) );
endmodule

