//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 0 0 1 1 0 1 0 0 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000;
  XNOR2_X1  g000(.A(G116), .B(G119), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT2), .B(G113), .ZN(new_n188));
  XOR2_X1   g002(.A(new_n187), .B(new_n188), .Z(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(G128), .A3(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n192), .A2(G146), .ZN(new_n198));
  OAI21_X1  g012(.A(G128), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT68), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n191), .A2(KEYINPUT65), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(new_n190), .A3(G143), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(new_n193), .A3(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n199), .A2(new_n200), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n200), .B1(new_n199), .B2(new_n204), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n197), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT11), .ZN(new_n209));
  INV_X1    g023(.A(G134), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(G137), .ZN(new_n211));
  AOI21_X1  g025(.A(G131), .B1(new_n210), .B2(G137), .ZN(new_n212));
  INV_X1    g026(.A(G137), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(KEYINPUT11), .A3(G134), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n211), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT66), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n211), .A2(new_n212), .A3(new_n217), .A4(new_n214), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n210), .A2(G137), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n213), .A2(G134), .ZN(new_n221));
  OAI21_X1  g035(.A(G131), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n189), .B1(new_n208), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n211), .A2(new_n214), .ZN(new_n225));
  OAI21_X1  g039(.A(G131), .B1(new_n225), .B2(new_n221), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n219), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n204), .A2(new_n232), .B1(new_n195), .B2(new_n230), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n219), .A2(KEYINPUT69), .A3(new_n226), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n229), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT28), .B1(new_n224), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(KEYINPUT70), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n229), .A2(new_n238), .A3(new_n233), .A4(new_n234), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n237), .A2(new_n239), .A3(new_n224), .ZN(new_n240));
  INV_X1    g054(.A(new_n189), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n208), .A2(new_n223), .B1(new_n227), .B2(new_n233), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n236), .B1(new_n243), .B2(KEYINPUT28), .ZN(new_n244));
  NOR2_X1   g058(.A1(G237), .A2(G953), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G210), .ZN(new_n246));
  XOR2_X1   g060(.A(new_n246), .B(KEYINPUT27), .Z(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT26), .B(G101), .ZN(new_n248));
  XOR2_X1   g062(.A(new_n247), .B(new_n248), .Z(new_n249));
  NOR2_X1   g063(.A1(new_n244), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n240), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT30), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n253), .B1(new_n208), .B2(new_n223), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n237), .A2(new_n239), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT71), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n237), .A2(new_n257), .A3(new_n239), .A4(new_n254), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n189), .B1(new_n242), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n252), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(KEYINPUT31), .B1(new_n263), .B2(new_n249), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n261), .B1(new_n256), .B2(new_n258), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT31), .ZN(new_n266));
  INV_X1    g080(.A(new_n249), .ZN(new_n267));
  NOR4_X1   g081(.A1(new_n265), .A2(new_n266), .A3(new_n252), .A4(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n251), .B1(new_n264), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT32), .ZN(new_n270));
  NOR2_X1   g084(.A1(G472), .A2(G902), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n270), .B1(new_n269), .B2(new_n271), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G472), .ZN(new_n275));
  INV_X1    g089(.A(G902), .ZN(new_n276));
  INV_X1    g090(.A(new_n236), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n240), .A2(KEYINPUT74), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT74), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n237), .A2(new_n279), .A3(new_n239), .A4(new_n224), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n208), .A2(new_n223), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n237), .A2(new_n281), .A3(new_n239), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n278), .A2(new_n280), .B1(new_n189), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT28), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n277), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n249), .A2(KEYINPUT29), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n276), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n288), .B1(new_n263), .B2(new_n249), .ZN(new_n289));
  OAI211_X1 g103(.A(KEYINPUT72), .B(new_n267), .C1(new_n265), .C2(new_n252), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT29), .B1(new_n244), .B2(new_n249), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n287), .B1(new_n292), .B2(KEYINPUT73), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT73), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n289), .A2(new_n294), .A3(new_n290), .A4(new_n291), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n275), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT75), .B1(new_n274), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n292), .A2(KEYINPUT73), .ZN(new_n298));
  INV_X1    g112(.A(new_n287), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n295), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G472), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n259), .A2(new_n262), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n240), .A3(new_n249), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n266), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n263), .A2(KEYINPUT31), .A3(new_n249), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n250), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n271), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT32), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n301), .A2(new_n302), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G469), .ZN(new_n313));
  INV_X1    g127(.A(G104), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G107), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n314), .A2(G107), .ZN(new_n317));
  OAI21_X1  g131(.A(G101), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT3), .B1(new_n314), .B2(G107), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT3), .ZN(new_n320));
  INV_X1    g134(.A(G107), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(G104), .ZN(new_n322));
  INV_X1    g136(.A(G101), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n319), .A2(new_n322), .A3(new_n323), .A4(new_n315), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n318), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT10), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT82), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n328), .B1(new_n191), .B2(KEYINPUT1), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n191), .A2(new_n328), .A3(KEYINPUT1), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G128), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n194), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n197), .ZN(new_n333));
  INV_X1    g147(.A(new_n325), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n208), .A2(new_n327), .B1(new_n335), .B2(new_n326), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n229), .A2(new_n234), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n319), .A2(new_n322), .A3(new_n315), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G101), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(KEYINPUT4), .A3(new_n324), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT4), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n338), .A2(new_n341), .A3(G101), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n233), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT81), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT81), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n340), .A2(new_n233), .A3(new_n345), .A4(new_n342), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n336), .A2(new_n337), .A3(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(G110), .B(G140), .ZN(new_n349));
  INV_X1    g163(.A(G953), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G227), .ZN(new_n351));
  XOR2_X1   g165(.A(new_n349), .B(new_n351), .Z(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  XOR2_X1   g168(.A(KEYINPUT83), .B(KEYINPUT12), .Z(new_n355));
  NAND2_X1  g169(.A1(new_n227), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n197), .B(new_n325), .C1(new_n206), .C2(new_n207), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n356), .B1(new_n357), .B2(new_n335), .ZN(new_n358));
  INV_X1    g172(.A(new_n337), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n335), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT12), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n358), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n354), .A2(new_n363), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n344), .A2(new_n346), .ZN(new_n365));
  INV_X1    g179(.A(new_n197), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n199), .A2(new_n204), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT68), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n366), .B1(new_n368), .B2(new_n205), .ZN(new_n369));
  INV_X1    g183(.A(new_n327), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n325), .B1(new_n332), .B2(new_n197), .ZN(new_n371));
  OAI22_X1  g185(.A1(new_n369), .A2(new_n370), .B1(KEYINPUT10), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n359), .B1(new_n365), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n353), .B1(new_n373), .B2(new_n348), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n313), .B(new_n276), .C1(new_n364), .C2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(KEYINPUT12), .B1(new_n359), .B2(new_n360), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n348), .B1(new_n376), .B2(new_n358), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n352), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n373), .A2(new_n348), .A3(new_n353), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(G469), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(G469), .A2(G902), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n375), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G221), .ZN(new_n383));
  XNOR2_X1  g197(.A(KEYINPUT9), .B(G234), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n383), .B1(new_n385), .B2(new_n276), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n382), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(G214), .B1(G237), .B2(G902), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(G210), .B1(G237), .B2(G902), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G224), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n393), .A2(G953), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NOR3_X1   g209(.A1(new_n208), .A2(KEYINPUT87), .A3(G125), .ZN(new_n396));
  INV_X1    g210(.A(G125), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT87), .B1(new_n233), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n398), .B1(new_n369), .B2(new_n397), .ZN(new_n399));
  OAI211_X1 g213(.A(KEYINPUT7), .B(new_n395), .C1(new_n396), .C2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n398), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n401), .B1(new_n208), .B2(G125), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT7), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT87), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n369), .A2(new_n404), .A3(new_n397), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n402), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n402), .A2(new_n394), .A3(new_n405), .ZN(new_n407));
  INV_X1    g221(.A(new_n187), .ZN(new_n408));
  OR2_X1    g222(.A1(new_n408), .A2(new_n188), .ZN(new_n409));
  XOR2_X1   g223(.A(KEYINPUT84), .B(KEYINPUT5), .Z(new_n410));
  INV_X1    g224(.A(G116), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(G119), .ZN(new_n412));
  AOI21_X1  g226(.A(KEYINPUT85), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  OR2_X1    g227(.A1(KEYINPUT84), .A2(KEYINPUT5), .ZN(new_n414));
  NAND2_X1  g228(.A1(KEYINPUT84), .A2(KEYINPUT5), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n412), .A2(new_n414), .A3(KEYINPUT85), .A4(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G113), .ZN(new_n417));
  OR2_X1    g231(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  OR2_X1    g232(.A1(new_n408), .A2(new_n410), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n409), .B(new_n334), .C1(new_n418), .C2(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(G110), .B(G122), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n189), .A2(new_n340), .A3(new_n342), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n400), .A2(new_n406), .A3(new_n407), .A4(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT90), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n416), .A2(G113), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n410), .A2(new_n412), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n427), .B(KEYINPUT88), .C1(new_n428), .C2(KEYINPUT85), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n187), .A2(KEYINPUT5), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT88), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n431), .B1(new_n413), .B2(new_n417), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n429), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n409), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT89), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT89), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n433), .A2(new_n436), .A3(new_n409), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n435), .A2(new_n437), .A3(new_n334), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n422), .B(KEYINPUT8), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n409), .B1(new_n418), .B2(new_n420), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n439), .B1(new_n440), .B2(new_n334), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n426), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n325), .B1(new_n434), .B2(KEYINPUT89), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n437), .ZN(new_n444));
  INV_X1    g258(.A(new_n441), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n445), .A3(KEYINPUT90), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n425), .B1(new_n442), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n395), .B1(new_n396), .B2(new_n399), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n407), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n421), .A2(new_n423), .ZN(new_n450));
  INV_X1    g264(.A(new_n422), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT6), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n450), .B(new_n451), .C1(KEYINPUT86), .C2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n450), .A2(new_n451), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n452), .A2(KEYINPUT86), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n424), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n449), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n276), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n392), .B1(new_n447), .B2(new_n458), .ZN(new_n459));
  AND4_X1   g273(.A1(new_n400), .A2(new_n406), .A3(new_n407), .A4(new_n424), .ZN(new_n460));
  AOI21_X1  g274(.A(KEYINPUT90), .B1(new_n444), .B2(new_n445), .ZN(new_n461));
  AOI211_X1 g275(.A(new_n426), .B(new_n441), .C1(new_n443), .C2(new_n437), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n463), .A2(new_n276), .A3(new_n391), .A4(new_n457), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n390), .B1(new_n459), .B2(new_n464), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n388), .A2(new_n465), .ZN(new_n466));
  XOR2_X1   g280(.A(G113), .B(G122), .Z(new_n467));
  XOR2_X1   g281(.A(KEYINPUT93), .B(G104), .Z(new_n468));
  XOR2_X1   g282(.A(new_n467), .B(new_n468), .Z(new_n469));
  NAND2_X1  g283(.A1(new_n245), .A2(G214), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(G143), .ZN(new_n471));
  INV_X1    g285(.A(G131), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n471), .B(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(KEYINPUT77), .A2(G125), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(G140), .ZN(new_n475));
  XOR2_X1   g289(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n476));
  XNOR2_X1  g290(.A(G125), .B(G140), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n475), .A2(KEYINPUT19), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n190), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n475), .A2(KEYINPUT16), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT16), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n481), .B1(new_n397), .B2(G140), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G146), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n473), .A2(new_n479), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT91), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT18), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n487), .A2(new_n472), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n486), .B1(new_n471), .B2(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n470), .B(new_n192), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(KEYINPUT91), .A3(new_n488), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n471), .A2(new_n489), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n475), .A2(G146), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n477), .A2(new_n190), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n493), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n469), .B1(new_n485), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n494), .A2(new_n497), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n500), .B1(new_n490), .B2(new_n492), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT17), .ZN(new_n502));
  NOR3_X1   g316(.A1(new_n471), .A2(new_n502), .A3(new_n472), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n471), .B(G131), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n503), .B1(new_n504), .B2(new_n502), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT78), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n480), .A2(new_n190), .A3(new_n482), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n484), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n483), .A2(KEYINPUT78), .A3(G146), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n501), .B1(new_n505), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n499), .B1(new_n511), .B2(new_n469), .ZN(new_n512));
  NOR2_X1   g326(.A1(G475), .A2(G902), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT20), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT20), .ZN(new_n516));
  INV_X1    g330(.A(new_n469), .ZN(new_n517));
  AOI211_X1 g331(.A(new_n517), .B(new_n501), .C1(new_n510), .C2(new_n505), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n516), .B(new_n513), .C1(new_n518), .C2(new_n499), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n511), .A2(new_n469), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n276), .B1(new_n521), .B2(new_n518), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(G475), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(G116), .B(G122), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n321), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT94), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(G128), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n529), .A2(G143), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n192), .A2(G128), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n532), .B(new_n210), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n411), .A2(KEYINPUT14), .A3(G122), .ZN(new_n534));
  INV_X1    g348(.A(new_n525), .ZN(new_n535));
  OAI211_X1 g349(.A(G107), .B(new_n534), .C1(new_n535), .C2(KEYINPUT14), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n528), .A2(new_n533), .A3(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n525), .B(new_n321), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n532), .A2(new_n210), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n530), .A2(KEYINPUT13), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n530), .A2(KEYINPUT13), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n540), .A2(new_n541), .A3(new_n531), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n538), .B(new_n539), .C1(new_n542), .C2(new_n210), .ZN(new_n543));
  INV_X1    g357(.A(G217), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n384), .A2(new_n544), .A3(G953), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n537), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n545), .B1(new_n537), .B2(new_n543), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(G478), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n549), .A2(KEYINPUT15), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n548), .A2(new_n276), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n551), .B1(new_n548), .B2(new_n276), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n524), .A2(new_n556), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n350), .A2(G952), .ZN(new_n558));
  INV_X1    g372(.A(G234), .ZN(new_n559));
  INV_X1    g373(.A(G237), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT21), .B(G898), .ZN(new_n563));
  XOR2_X1   g377(.A(new_n563), .B(KEYINPUT95), .Z(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  AOI211_X1 g379(.A(new_n276), .B(new_n350), .C1(G234), .C2(G237), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n562), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(G119), .B(G128), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT76), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n569), .B(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT24), .B(G110), .ZN(new_n572));
  OR2_X1    g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT23), .ZN(new_n574));
  INV_X1    g388(.A(G119), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n574), .B1(new_n575), .B2(G128), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n529), .A2(KEYINPUT23), .A3(G119), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n576), .B(new_n577), .C1(G119), .C2(new_n529), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(G110), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n508), .A2(new_n509), .A3(new_n573), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n571), .A2(new_n572), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT79), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n582), .B1(new_n578), .B2(G110), .ZN(new_n583));
  OR3_X1    g397(.A1(new_n578), .A2(new_n582), .A3(G110), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(new_n496), .A3(new_n484), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n580), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(KEYINPUT22), .B(G137), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n383), .A2(new_n559), .A3(G953), .ZN(new_n589));
  XOR2_X1   g403(.A(new_n588), .B(new_n589), .Z(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n580), .A2(new_n586), .A3(new_n590), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n544), .B1(G234), .B2(new_n276), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(G902), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT80), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n599), .A2(KEYINPUT25), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n600), .B1(new_n594), .B2(G902), .ZN(new_n601));
  INV_X1    g415(.A(new_n600), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n592), .A2(new_n276), .A3(new_n593), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n598), .B1(new_n604), .B2(new_n595), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n557), .A2(new_n568), .A3(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n297), .A2(new_n312), .A3(new_n466), .A4(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT96), .B(G101), .Z(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G3));
  NAND3_X1  g423(.A1(new_n548), .A2(new_n549), .A3(new_n276), .ZN(new_n610));
  NAND2_X1  g424(.A1(G478), .A2(G902), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT33), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n548), .B(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n612), .B1(new_n614), .B2(G478), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n524), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n465), .A2(new_n568), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT97), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT97), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n465), .A2(new_n619), .A3(new_n568), .A4(new_n616), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n269), .A2(new_n276), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(G472), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n269), .A2(new_n271), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n623), .A2(new_n624), .A3(new_n388), .A4(new_n605), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT34), .B(G104), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  NOR2_X1   g442(.A1(new_n524), .A2(new_n555), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n465), .A2(new_n568), .A3(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT98), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n465), .A2(new_n629), .A3(KEYINPUT98), .A4(new_n568), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n634), .A2(new_n625), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT35), .B(G107), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G9));
  NAND2_X1  g451(.A1(new_n459), .A2(new_n464), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n389), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n587), .A2(KEYINPUT99), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT99), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n580), .A2(new_n586), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n591), .A2(KEYINPUT36), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n596), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n604), .A2(new_n595), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(new_n557), .A3(new_n568), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n639), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n650), .A2(new_n623), .A3(new_n624), .A4(new_n388), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT37), .B(G110), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G12));
  NAND2_X1  g467(.A1(new_n388), .A2(new_n648), .ZN(new_n654));
  INV_X1    g468(.A(G900), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n562), .B1(new_n566), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n629), .A2(new_n657), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n654), .A2(new_n639), .A3(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n297), .A2(new_n312), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G128), .ZN(G30));
  INV_X1    g475(.A(KEYINPUT38), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n638), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n524), .A2(new_n556), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n663), .A2(new_n390), .A3(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n283), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n276), .B1(new_n666), .B2(new_n249), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n263), .A2(new_n267), .ZN(new_n668));
  OAI21_X1  g482(.A(G472), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n311), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n648), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n665), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(KEYINPUT100), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n656), .B(KEYINPUT39), .Z(new_n674));
  NAND2_X1  g488(.A1(new_n388), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT101), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(KEYINPUT40), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n675), .B(KEYINPUT101), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT40), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT100), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n665), .A2(new_n670), .A3(new_n683), .A4(new_n671), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n673), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT102), .B(G143), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G45));
  NAND3_X1  g501(.A1(new_n524), .A2(new_n615), .A3(new_n657), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n671), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n297), .A2(new_n312), .A3(new_n466), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G146), .ZN(G48));
  NAND2_X1  g505(.A1(new_n373), .A2(new_n348), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n352), .ZN(new_n693));
  OAI211_X1 g507(.A(new_n348), .B(new_n353), .C1(new_n376), .C2(new_n358), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n313), .B1(new_n695), .B2(new_n276), .ZN(new_n696));
  AOI211_X1 g510(.A(G469), .B(G902), .C1(new_n693), .C2(new_n694), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n387), .ZN(new_n699));
  INV_X1    g513(.A(new_n605), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n618), .A2(new_n620), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n297), .A2(new_n312), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT41), .B(G113), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G15));
  NAND2_X1  g519(.A1(new_n297), .A2(new_n312), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n632), .A2(new_n633), .A3(new_n701), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G116), .ZN(G18));
  NOR2_X1   g524(.A1(new_n639), .A2(new_n699), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n649), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n707), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G119), .ZN(G21));
  NAND2_X1  g529(.A1(new_n285), .A2(new_n267), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n716), .B1(new_n264), .B2(new_n268), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n622), .A2(G472), .B1(new_n271), .B2(new_n717), .ZN(new_n718));
  XOR2_X1   g532(.A(new_n605), .B(KEYINPUT103), .Z(new_n719));
  AND2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n664), .A2(new_n567), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n720), .A2(new_n711), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G122), .ZN(G24));
  NOR3_X1   g537(.A1(new_n639), .A2(new_n699), .A3(new_n688), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n718), .A2(new_n724), .A3(new_n648), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT104), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT104), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n718), .A2(new_n724), .A3(new_n727), .A4(new_n648), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G125), .ZN(G27));
  INV_X1    g544(.A(KEYINPUT42), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n382), .A2(KEYINPUT105), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT105), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n375), .A2(new_n733), .A3(new_n380), .A4(new_n381), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n732), .A2(new_n387), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n459), .A2(new_n464), .A3(new_n389), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n688), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n297), .A2(new_n312), .A3(new_n605), .A4(new_n738), .ZN(new_n739));
  NOR4_X1   g553(.A1(new_n735), .A2(new_n731), .A3(new_n736), .A4(new_n688), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n719), .B(new_n740), .C1(new_n274), .C2(new_n296), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT106), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n301), .A2(new_n311), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n744), .A2(KEYINPUT106), .A3(new_n719), .A4(new_n740), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n731), .A2(new_n739), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n472), .ZN(G33));
  NOR2_X1   g561(.A1(new_n737), .A2(new_n658), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n297), .A2(new_n312), .A3(new_n605), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G134), .ZN(G36));
  NAND2_X1  g564(.A1(new_n378), .A2(new_n379), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n378), .A2(KEYINPUT45), .A3(new_n379), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(G469), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n381), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT46), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n755), .A2(KEYINPUT46), .A3(new_n381), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(new_n375), .A3(new_n759), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n760), .A2(new_n387), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n761), .A2(new_n674), .ZN(new_n762));
  INV_X1    g576(.A(new_n736), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n623), .A2(new_n624), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n615), .A2(new_n523), .A3(new_n520), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT43), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n671), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n764), .A2(KEYINPUT44), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n764), .A2(new_n767), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n762), .A2(new_n763), .A3(new_n768), .A4(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G137), .ZN(G39));
  XNOR2_X1  g587(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n760), .A2(new_n387), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n774), .B1(new_n760), .B2(new_n387), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n736), .A2(new_n605), .A3(new_n688), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n706), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G140), .ZN(G42));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n617), .A2(new_n630), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n651), .B1(new_n625), .B2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n607), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT109), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n607), .A2(KEYINPUT109), .A3(new_n784), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n739), .A2(new_n731), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n743), .A2(new_n745), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n297), .B(new_n312), .C1(new_n708), .C2(new_n713), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(new_n703), .A3(new_n722), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n557), .A2(new_n657), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n654), .A2(new_n736), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n297), .A2(new_n312), .A3(new_n796), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n718), .A2(new_n648), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n738), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n749), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n794), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n789), .A2(new_n792), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n465), .A2(new_n556), .A3(new_n524), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n803), .A2(new_n656), .A3(new_n735), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n670), .A2(new_n671), .A3(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n690), .A2(new_n729), .A3(new_n660), .A4(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT52), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n781), .B1(new_n802), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT110), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n806), .B(new_n810), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n746), .A2(new_n794), .A3(new_n800), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n811), .A2(new_n812), .A3(KEYINPUT53), .A4(new_n789), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n808), .A2(new_n809), .A3(new_n813), .ZN(new_n814));
  OAI211_X1 g628(.A(KEYINPUT110), .B(new_n781), .C1(new_n802), .C2(new_n807), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(KEYINPUT54), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n794), .B(KEYINPUT111), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n749), .A2(new_n797), .A3(KEYINPUT53), .A4(new_n799), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n746), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n811), .A2(new_n817), .A3(new_n789), .A4(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n808), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n816), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n766), .A2(new_n561), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n720), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n558), .B1(new_n825), .B2(new_n712), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n744), .A2(new_n719), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n699), .A2(new_n736), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n829), .A2(new_n766), .A3(new_n561), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  XOR2_X1   g645(.A(new_n831), .B(KEYINPUT48), .Z(new_n832));
  NOR4_X1   g646(.A1(new_n670), .A2(new_n561), .A3(new_n700), .A4(new_n829), .ZN(new_n833));
  AOI211_X1 g647(.A(new_n826), .B(new_n832), .C1(new_n616), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n798), .A2(new_n830), .ZN(new_n835));
  XOR2_X1   g649(.A(new_n835), .B(KEYINPUT113), .Z(new_n836));
  NOR2_X1   g650(.A1(new_n524), .A2(new_n615), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n836), .B1(new_n833), .B2(new_n837), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n698), .B(KEYINPUT108), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n840), .A2(KEYINPUT112), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(KEYINPUT112), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n841), .A2(new_n386), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n843), .B1(new_n775), .B2(new_n776), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n825), .A2(new_n736), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n844), .A2(new_n845), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n663), .ZN(new_n850));
  NOR4_X1   g664(.A1(new_n825), .A2(new_n389), .A3(new_n850), .A4(new_n699), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT50), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n838), .A2(new_n849), .A3(new_n852), .A4(KEYINPUT51), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n838), .A2(new_n852), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n844), .A2(new_n847), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n834), .B(new_n853), .C1(KEYINPUT51), .C2(new_n856), .ZN(new_n857));
  OAI22_X1  g671(.A1(new_n823), .A2(new_n857), .B1(G952), .B2(G953), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n839), .A2(KEYINPUT49), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n765), .A2(new_n390), .A3(new_n386), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n719), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n862), .B(new_n663), .C1(KEYINPUT49), .C2(new_n839), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n858), .B1(new_n670), .B2(new_n863), .ZN(G75));
  INV_X1    g678(.A(KEYINPUT116), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n456), .A2(new_n453), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n866), .A2(new_n448), .A3(new_n407), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n457), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(KEYINPUT55), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(G210), .A2(G902), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n793), .A2(new_n703), .A3(new_n722), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n749), .A2(new_n797), .A3(new_n799), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n792), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n607), .A2(KEYINPUT109), .A3(new_n784), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT109), .B1(new_n607), .B2(new_n784), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT53), .B1(new_n879), .B2(new_n811), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT111), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n703), .A2(new_n722), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n881), .B1(new_n882), .B2(new_n793), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n794), .A2(KEYINPUT111), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n819), .B(new_n789), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n885), .A2(new_n807), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n872), .B1(new_n880), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT56), .B1(new_n887), .B2(KEYINPUT115), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n871), .B1(new_n808), .B2(new_n820), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT115), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n870), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT56), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n887), .A2(new_n893), .A3(new_n870), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n350), .A2(G952), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n865), .B1(new_n892), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n893), .B1(new_n889), .B2(new_n890), .ZN(new_n899));
  AOI211_X1 g713(.A(KEYINPUT115), .B(new_n871), .C1(new_n808), .C2(new_n820), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n869), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n901), .A2(KEYINPUT116), .A3(new_n896), .A4(new_n894), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n898), .A2(new_n902), .ZN(G51));
  XOR2_X1   g717(.A(new_n381), .B(KEYINPUT57), .Z(new_n904));
  AND3_X1   g718(.A1(new_n808), .A2(new_n821), .A3(new_n820), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n821), .B1(new_n808), .B2(new_n820), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n695), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n880), .A2(new_n886), .ZN(new_n909));
  OR3_X1    g723(.A1(new_n909), .A2(new_n276), .A3(new_n755), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n895), .B1(new_n908), .B2(new_n910), .ZN(G54));
  NAND2_X1  g725(.A1(KEYINPUT58), .A2(G475), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n909), .A2(new_n276), .A3(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n512), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n896), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n915), .B1(new_n914), .B2(new_n913), .ZN(G60));
  INV_X1    g730(.A(new_n614), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n611), .B(KEYINPUT118), .ZN(new_n918));
  XNOR2_X1  g732(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n917), .B(new_n920), .C1(new_n905), .C2(new_n906), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT119), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n921), .A2(new_n922), .A3(new_n896), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n922), .B1(new_n921), .B2(new_n896), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n917), .B1(new_n823), .B2(new_n920), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(G63));
  OAI21_X1  g740(.A(new_n896), .B1(KEYINPUT120), .B2(KEYINPUT61), .ZN(new_n927));
  NAND2_X1  g741(.A1(G217), .A2(G902), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT60), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n909), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n927), .B1(new_n930), .B2(new_n645), .ZN(new_n931));
  NAND2_X1  g745(.A1(KEYINPUT120), .A2(KEYINPUT61), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n594), .B1(new_n909), .B2(new_n929), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n932), .B1(new_n931), .B2(new_n933), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n934), .A2(new_n935), .ZN(G66));
  AOI21_X1  g750(.A(new_n350), .B1(new_n564), .B2(G224), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n789), .A2(new_n873), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n937), .B1(new_n938), .B2(new_n350), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n866), .B1(G898), .B2(new_n350), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n939), .B(new_n940), .Z(G69));
  OAI21_X1  g755(.A(new_n259), .B1(new_n242), .B2(new_n260), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(new_n478), .Z(new_n943));
  NAND2_X1  g757(.A1(new_n707), .A2(new_n605), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n677), .B(new_n763), .C1(new_n616), .C2(new_n629), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n772), .B(new_n779), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n690), .A2(new_n729), .A3(new_n660), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n685), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n946), .B1(new_n948), .B2(KEYINPUT62), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n947), .A2(new_n685), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT121), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT121), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n948), .A2(new_n953), .A3(KEYINPUT62), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n949), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n943), .B1(new_n955), .B2(new_n350), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n761), .A2(new_n674), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n957), .A2(new_n803), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n827), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(KEYINPUT122), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT122), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n958), .A2(new_n961), .A3(new_n827), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n772), .A2(new_n779), .A3(new_n749), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n963), .A2(new_n964), .A3(new_n792), .A4(new_n947), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n965), .A2(G953), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n943), .B1(new_n655), .B2(new_n350), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OR3_X1    g782(.A1(new_n956), .A2(KEYINPUT123), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n350), .B1(G227), .B2(G900), .ZN(new_n970));
  OAI21_X1  g784(.A(KEYINPUT123), .B1(new_n956), .B2(new_n968), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n970), .B1(new_n969), .B2(new_n971), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n972), .A2(new_n973), .ZN(G72));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n975));
  INV_X1    g789(.A(new_n938), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n976), .B(new_n949), .C1(new_n952), .C2(new_n954), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT125), .ZN(new_n978));
  XNOR2_X1  g792(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n275), .A2(new_n276), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n979), .B(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n977), .A2(new_n978), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n668), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n978), .B1(new_n977), .B2(new_n981), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n289), .A2(new_n304), .A3(new_n290), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n814), .A2(new_n815), .A3(new_n981), .A4(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT126), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n981), .B1(new_n965), .B2(new_n938), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n263), .A2(new_n267), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n988), .B1(new_n992), .B2(new_n896), .ZN(new_n993));
  AOI211_X1 g807(.A(KEYINPUT126), .B(new_n895), .C1(new_n989), .C2(new_n991), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n987), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n975), .B1(new_n985), .B2(new_n995), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n993), .A2(new_n994), .ZN(new_n997));
  INV_X1    g811(.A(new_n984), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n998), .A2(new_n668), .A3(new_n982), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n997), .A2(new_n999), .A3(KEYINPUT127), .A4(new_n987), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n996), .A2(new_n1000), .ZN(G57));
endmodule


