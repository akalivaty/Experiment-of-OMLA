//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 0 1 1 0 1 0 0 1 0 0 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962;
  INV_X1    g000(.A(KEYINPUT25), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT77), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT16), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(G125), .ZN(new_n192));
  INV_X1    g006(.A(G125), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G140), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n191), .B1(new_n195), .B2(new_n189), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  OR2_X1    g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n197), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT70), .B(G128), .ZN(new_n201));
  INV_X1    g015(.A(G119), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n203), .B1(new_n202), .B2(G128), .ZN(new_n204));
  XOR2_X1   g018(.A(KEYINPUT24), .B(G110), .Z(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT75), .B(KEYINPUT23), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n207), .B1(new_n202), .B2(G128), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(G119), .B2(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n210), .B1(KEYINPUT23), .B2(new_n203), .ZN(new_n211));
  INV_X1    g025(.A(G110), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n200), .B(new_n206), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n204), .A2(new_n205), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT76), .B(G110), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n214), .B1(new_n211), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(G125), .B(G140), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(new_n197), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n198), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n213), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT22), .B(G137), .ZN(new_n221));
  INV_X1    g035(.A(G221), .ZN(new_n222));
  INV_X1    g036(.A(G234), .ZN(new_n223));
  NOR3_X1   g037(.A1(new_n222), .A2(new_n223), .A3(G953), .ZN(new_n224));
  XOR2_X1   g038(.A(new_n221), .B(new_n224), .Z(new_n225));
  XNOR2_X1  g039(.A(new_n220), .B(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n188), .B1(new_n227), .B2(G902), .ZN(new_n228));
  INV_X1    g042(.A(G902), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G234), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n226), .A2(KEYINPUT77), .A3(new_n187), .A4(new_n229), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n228), .A2(G217), .A3(new_n230), .A4(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(G902), .B1(new_n223), .B2(G217), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n226), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT82), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT81), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT11), .ZN(new_n238));
  INV_X1    g052(.A(G134), .ZN(new_n239));
  NOR3_X1   g053(.A1(new_n238), .A2(new_n239), .A3(G137), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT65), .B(G134), .ZN(new_n241));
  INV_X1    g055(.A(G137), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT67), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT67), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT65), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n245), .A2(G134), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n239), .A2(KEYINPUT65), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n244), .B(G137), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n240), .B1(new_n243), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G131), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n239), .A2(KEYINPUT65), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n245), .A2(G134), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(new_n242), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n251), .B1(new_n254), .B2(new_n238), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n254), .A2(new_n251), .A3(new_n238), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n249), .A2(new_n250), .A3(new_n256), .A4(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n257), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(new_n255), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n262), .A2(KEYINPUT68), .A3(new_n250), .A4(new_n249), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n249), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G131), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT10), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n197), .A2(G143), .ZN(new_n269));
  INV_X1    g083(.A(G143), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G146), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n269), .A2(new_n271), .A3(G128), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT1), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT1), .B1(new_n270), .B2(G146), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G128), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n269), .A2(new_n271), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n272), .A2(new_n273), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n278));
  INV_X1    g092(.A(G107), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n278), .A2(G104), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G104), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n281), .A2(G107), .B1(KEYINPUT79), .B2(KEYINPUT3), .ZN(new_n282));
  OAI22_X1  g096(.A1(new_n281), .A2(G107), .B1(KEYINPUT79), .B2(KEYINPUT3), .ZN(new_n283));
  INV_X1    g097(.A(G101), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n280), .A2(new_n282), .A3(new_n283), .A4(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n281), .A2(G107), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n279), .A2(G104), .ZN(new_n287));
  OAI21_X1  g101(.A(G101), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n268), .B1(new_n277), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT80), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n201), .B1(KEYINPUT69), .B2(new_n274), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n274), .A2(KEYINPUT69), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n276), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n276), .A2(KEYINPUT1), .A3(new_n209), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n289), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(KEYINPUT10), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n280), .A2(new_n282), .A3(new_n283), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G101), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(KEYINPUT4), .A3(new_n285), .ZN(new_n302));
  NAND2_X1  g116(.A1(KEYINPUT0), .A2(G128), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT0), .B(G128), .ZN(new_n304));
  MUX2_X1   g118(.A(new_n303), .B(new_n304), .S(new_n276), .Z(new_n305));
  INV_X1    g119(.A(KEYINPUT4), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n300), .A2(new_n306), .A3(G101), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n302), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n274), .A2(G128), .B1(new_n269), .B2(new_n271), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n288), .B(new_n285), .C1(new_n295), .C2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT80), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(new_n311), .A3(new_n268), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n291), .A2(new_n299), .A3(new_n308), .A4(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n237), .B1(new_n267), .B2(new_n313), .ZN(new_n314));
  AND4_X1   g128(.A1(new_n308), .A2(new_n291), .A3(new_n299), .A4(new_n312), .ZN(new_n315));
  AOI22_X1  g129(.A1(new_n260), .A2(new_n263), .B1(G131), .B2(new_n265), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(KEYINPUT81), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G953), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G227), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(new_n190), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT78), .B(G110), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n321), .B(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n267), .A2(new_n313), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n318), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT12), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n310), .B1(new_n297), .B2(new_n298), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n327), .B1(new_n267), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n328), .ZN(new_n330));
  NOR3_X1   g144(.A1(new_n316), .A2(KEYINPUT12), .A3(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n323), .B1(new_n332), .B2(new_n318), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n326), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n236), .B(G469), .C1(new_n334), .C2(G902), .ZN(new_n335));
  INV_X1    g149(.A(new_n323), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n267), .A2(new_n237), .A3(new_n313), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT81), .B1(new_n315), .B2(new_n316), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n267), .A2(new_n327), .A3(new_n328), .ZN(new_n340));
  OAI21_X1  g154(.A(KEYINPUT12), .B1(new_n316), .B2(new_n330), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n336), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(G902), .B1(new_n343), .B2(new_n325), .ZN(new_n344));
  INV_X1    g158(.A(G469), .ZN(new_n345));
  OAI21_X1  g159(.A(KEYINPUT82), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n324), .B1(new_n337), .B2(new_n338), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n336), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n332), .A2(new_n318), .A3(new_n323), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(new_n345), .A3(new_n229), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n335), .A2(new_n346), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G475), .ZN(new_n353));
  NOR2_X1   g167(.A1(G237), .A2(G953), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(G143), .A3(G214), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(G143), .B1(new_n354), .B2(G214), .ZN(new_n357));
  OAI21_X1  g171(.A(G131), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT17), .ZN(new_n359));
  INV_X1    g173(.A(G237), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(new_n319), .A3(G214), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n270), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(new_n250), .A3(new_n355), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n358), .A2(new_n359), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT91), .ZN(new_n365));
  OR2_X1    g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n200), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n250), .B1(new_n362), .B2(new_n355), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT17), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n364), .A2(new_n365), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n366), .A2(new_n367), .A3(new_n369), .A4(new_n370), .ZN(new_n371));
  AND2_X1   g185(.A1(KEYINPUT87), .A2(KEYINPUT18), .ZN(new_n372));
  OAI211_X1 g186(.A(G131), .B(new_n372), .C1(new_n356), .C2(new_n357), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n195), .A2(G146), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n218), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n372), .A2(G131), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n362), .A2(new_n355), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n373), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT88), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT88), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n373), .A2(new_n375), .A3(new_n377), .A4(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n371), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(G113), .B(G122), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(new_n281), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n371), .A2(new_n385), .A3(new_n382), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n353), .B1(new_n389), .B2(new_n229), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT89), .ZN(new_n391));
  INV_X1    g205(.A(new_n363), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n391), .B1(new_n392), .B2(new_n368), .ZN(new_n393));
  OR2_X1    g207(.A1(new_n195), .A2(KEYINPUT19), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n195), .A2(KEYINPUT19), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n197), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n358), .A2(KEYINPUT89), .A3(new_n363), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n393), .A2(new_n198), .A3(new_n396), .A4(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n382), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT90), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n382), .A2(new_n398), .A3(KEYINPUT90), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n386), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n388), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(new_n353), .A3(new_n229), .ZN(new_n405));
  XNOR2_X1  g219(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT20), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n404), .A2(new_n408), .A3(new_n353), .A4(new_n229), .ZN(new_n409));
  AOI211_X1 g223(.A(KEYINPUT92), .B(new_n390), .C1(new_n407), .C2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT92), .ZN(new_n411));
  AOI211_X1 g225(.A(G475), .B(G902), .C1(new_n403), .C2(new_n388), .ZN(new_n412));
  INV_X1    g226(.A(new_n406), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n409), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n390), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n411), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n270), .A2(G128), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n417), .B1(new_n201), .B2(new_n270), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n418), .A2(new_n241), .ZN(new_n419));
  OR2_X1    g233(.A1(new_n419), .A2(KEYINPUT93), .ZN(new_n420));
  XOR2_X1   g234(.A(G116), .B(G122), .Z(new_n421));
  OR2_X1    g235(.A1(new_n421), .A2(G107), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(G107), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT13), .ZN(new_n425));
  OAI22_X1  g239(.A1(new_n201), .A2(new_n270), .B1(new_n425), .B2(new_n417), .ZN(new_n426));
  AOI21_X1  g240(.A(KEYINPUT13), .B1(new_n270), .B2(G128), .ZN(new_n427));
  OAI21_X1  g241(.A(G134), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n419), .A2(KEYINPUT93), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n420), .A2(new_n424), .A3(new_n428), .A4(new_n429), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n418), .A2(new_n241), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n422), .B1(new_n431), .B2(new_n419), .ZN(new_n432));
  INV_X1    g246(.A(G116), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(KEYINPUT14), .A3(G122), .ZN(new_n434));
  OAI211_X1 g248(.A(G107), .B(new_n434), .C1(new_n421), .C2(KEYINPUT14), .ZN(new_n435));
  XOR2_X1   g249(.A(new_n435), .B(KEYINPUT94), .Z(new_n436));
  OAI21_X1  g250(.A(new_n430), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  XOR2_X1   g251(.A(KEYINPUT9), .B(G234), .Z(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(G217), .A3(new_n319), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n437), .A2(new_n439), .ZN(new_n442));
  OAI211_X1 g256(.A(KEYINPUT95), .B(new_n229), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G478), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(KEYINPUT15), .ZN(new_n445));
  OR2_X1    g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n229), .B1(new_n441), .B2(new_n442), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT95), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n445), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n443), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n446), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n410), .A2(new_n416), .A3(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(G214), .B1(G237), .B2(G902), .ZN(new_n453));
  XOR2_X1   g267(.A(new_n453), .B(KEYINPUT83), .Z(new_n454));
  XOR2_X1   g268(.A(new_n454), .B(KEYINPUT84), .Z(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n319), .A2(G952), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n457), .B1(G234), .B2(G237), .ZN(new_n458));
  XOR2_X1   g272(.A(KEYINPUT21), .B(G898), .Z(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  OAI211_X1 g274(.A(G902), .B(G953), .C1(new_n223), .C2(new_n360), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n458), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n297), .A2(new_n193), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n305), .A2(G125), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(G224), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n467), .A2(G953), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n468), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n464), .A2(new_n470), .A3(new_n465), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n469), .B(new_n471), .C1(KEYINPUT7), .C2(new_n468), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT5), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(new_n202), .A3(G116), .ZN(new_n474));
  XOR2_X1   g288(.A(G116), .B(G119), .Z(new_n475));
  OAI211_X1 g289(.A(G113), .B(new_n474), .C1(new_n475), .C2(new_n473), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT2), .B(G113), .ZN(new_n477));
  OR2_X1    g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n298), .ZN(new_n480));
  XOR2_X1   g294(.A(G110), .B(G122), .Z(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n302), .A2(new_n307), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n475), .B(new_n477), .Z(new_n484));
  OAI211_X1 g298(.A(new_n480), .B(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n298), .A2(KEYINPUT85), .ZN(new_n486));
  OR2_X1    g300(.A1(new_n486), .A2(new_n479), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n479), .ZN(new_n488));
  XOR2_X1   g302(.A(new_n481), .B(KEYINPUT8), .Z(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  OR3_X1    g304(.A1(new_n466), .A2(KEYINPUT7), .A3(new_n468), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n472), .A2(new_n485), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n480), .B1(new_n483), .B2(new_n484), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n481), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(KEYINPUT6), .A3(new_n485), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n469), .A2(new_n471), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT6), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n493), .A2(new_n497), .A3(new_n481), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n495), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n492), .A2(new_n499), .A3(new_n229), .ZN(new_n500));
  OAI21_X1  g314(.A(G210), .B1(G237), .B2(G902), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n492), .A2(new_n499), .A3(new_n229), .A4(new_n501), .ZN(new_n504));
  AOI211_X1 g318(.A(new_n456), .B(new_n463), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n222), .B1(new_n438), .B2(new_n229), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n352), .A2(new_n452), .A3(new_n505), .A4(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(G472), .A2(G902), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n354), .A2(G210), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(new_n284), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n512));
  XOR2_X1   g326(.A(new_n511), .B(new_n512), .Z(new_n513));
  INV_X1    g327(.A(new_n484), .ZN(new_n514));
  INV_X1    g328(.A(new_n305), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n515), .B1(new_n264), .B2(new_n266), .ZN(new_n516));
  INV_X1    g330(.A(new_n297), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n239), .A2(G137), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n250), .B1(new_n254), .B2(new_n518), .ZN(new_n519));
  AOI211_X1 g333(.A(new_n517), .B(new_n519), .C1(new_n260), .C2(new_n263), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n514), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n519), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n264), .A2(new_n297), .A3(new_n522), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n523), .B(new_n484), .C1(new_n316), .C2(new_n515), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  XOR2_X1   g339(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(KEYINPUT72), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT72), .ZN(new_n529));
  AOI211_X1 g343(.A(new_n529), .B(new_n526), .C1(new_n521), .C2(new_n524), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT73), .B1(new_n516), .B2(new_n520), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT73), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n523), .B(new_n533), .C1(new_n316), .C2(new_n515), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n532), .A2(new_n534), .A3(new_n484), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT28), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n513), .B1(new_n531), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n539), .B1(new_n516), .B2(new_n520), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n523), .B(KEYINPUT30), .C1(new_n316), .C2(new_n515), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n541), .A3(new_n514), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n542), .A2(new_n513), .A3(new_n524), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT31), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT31), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n542), .A2(new_n545), .A3(new_n513), .A4(new_n524), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  OAI211_X1 g361(.A(KEYINPUT32), .B(new_n509), .C1(new_n538), .C2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT74), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n525), .A2(new_n527), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n529), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n525), .A2(KEYINPUT72), .A3(new_n527), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n537), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n513), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n544), .A2(new_n546), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n558), .A2(KEYINPUT74), .A3(KEYINPUT32), .A4(new_n509), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n550), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n525), .A2(KEYINPUT28), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n537), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n513), .A2(KEYINPUT29), .ZN(new_n563));
  AOI21_X1  g377(.A(G902), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n542), .A2(new_n524), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n565), .A2(new_n513), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n566), .B1(new_n554), .B2(new_n513), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n564), .B1(new_n567), .B2(KEYINPUT29), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n509), .B1(new_n538), .B2(new_n547), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT32), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n568), .A2(G472), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AOI211_X1 g385(.A(new_n235), .B(new_n508), .C1(new_n560), .C2(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(new_n284), .ZN(G3));
  AOI211_X1 g387(.A(G469), .B(G902), .C1(new_n348), .C2(new_n349), .ZN(new_n574));
  OAI21_X1  g388(.A(G469), .B1(new_n334), .B2(G902), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n574), .B1(new_n575), .B2(KEYINPUT82), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n506), .B1(new_n576), .B2(new_n335), .ZN(new_n577));
  INV_X1    g391(.A(new_n235), .ZN(new_n578));
  AOI21_X1  g392(.A(G902), .B1(new_n556), .B2(new_n557), .ZN(new_n579));
  INV_X1    g393(.A(G472), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(KEYINPUT96), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n547), .B1(new_n555), .B2(new_n554), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n581), .B1(new_n584), .B2(G902), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n577), .A2(new_n578), .A3(new_n583), .A4(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n410), .A2(new_n416), .ZN(new_n588));
  INV_X1    g402(.A(new_n442), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n589), .A2(KEYINPUT33), .A3(new_n440), .ZN(new_n590));
  AOI21_X1  g404(.A(KEYINPUT33), .B1(new_n589), .B2(new_n440), .ZN(new_n591));
  OAI21_X1  g405(.A(G478), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OR2_X1    g406(.A1(new_n447), .A2(G478), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n444), .A2(new_n229), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n588), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n454), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n463), .B1(new_n503), .B2(new_n504), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n587), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT34), .B(G104), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G6));
  MUX2_X1   g417(.A(new_n445), .B(new_n449), .S(new_n443), .Z(new_n604));
  NOR2_X1   g418(.A1(new_n604), .A2(new_n454), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n412), .A2(new_n413), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n390), .B1(new_n606), .B2(new_n407), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n605), .A2(new_n599), .A3(new_n607), .ZN(new_n608));
  XOR2_X1   g422(.A(new_n608), .B(KEYINPUT97), .Z(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n587), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(KEYINPUT98), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT35), .B(G107), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G9));
  INV_X1    g427(.A(new_n585), .ZN(new_n614));
  INV_X1    g428(.A(new_n583), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n352), .A2(new_n452), .A3(new_n507), .ZN(new_n617));
  INV_X1    g431(.A(new_n225), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(KEYINPUT36), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n220), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n233), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n232), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n616), .A2(new_n505), .A3(new_n617), .A4(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT37), .B(G110), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G12));
  INV_X1    g439(.A(new_n622), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n626), .B1(new_n560), .B2(new_n571), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT100), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n458), .B(KEYINPUT99), .ZN(new_n629));
  INV_X1    g443(.A(G900), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n629), .B1(new_n630), .B2(new_n462), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n607), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n628), .B1(new_n633), .B2(new_n604), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n451), .A2(new_n607), .A3(KEYINPUT100), .A4(new_n632), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n454), .B1(new_n503), .B2(new_n504), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n627), .A2(new_n577), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G128), .ZN(G30));
  XNOR2_X1  g453(.A(new_n631), .B(KEYINPUT39), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n577), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT40), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n569), .A2(new_n570), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n565), .A2(new_n513), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n229), .B1(new_n525), .B2(new_n513), .ZN(new_n647));
  OAI21_X1  g461(.A(G472), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n560), .A2(new_n644), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n414), .A2(new_n415), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT92), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n414), .A2(new_n411), .A3(new_n415), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n653), .A2(new_n605), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n503), .A2(new_n504), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT38), .ZN(new_n656));
  AND4_X1   g470(.A1(new_n643), .A2(new_n649), .A3(new_n654), .A4(new_n656), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n657), .B(new_n626), .C1(KEYINPUT40), .C2(new_n642), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G143), .ZN(G45));
  AOI211_X1 g473(.A(new_n631), .B(new_n596), .C1(new_n651), .C2(new_n652), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n627), .A2(new_n577), .A3(new_n637), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G146), .ZN(G48));
  AOI21_X1  g476(.A(new_n235), .B1(new_n560), .B2(new_n571), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n345), .B1(new_n350), .B2(new_n229), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n574), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n507), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n663), .A2(new_n600), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT41), .B(G113), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G15));
  NAND3_X1  g484(.A1(new_n663), .A2(new_n609), .A3(new_n667), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G116), .ZN(G18));
  NAND2_X1  g486(.A1(new_n560), .A2(new_n571), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n651), .A2(new_n652), .A3(new_n604), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n350), .A2(new_n229), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(G469), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n676), .A2(new_n507), .A3(new_n351), .A4(new_n637), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(KEYINPUT101), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT101), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n665), .A2(new_n679), .A3(new_n507), .A4(new_n637), .ZN(new_n680));
  AOI211_X1 g494(.A(new_n463), .B(new_n674), .C1(new_n678), .C2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n673), .A2(new_n681), .A3(new_n622), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n627), .A2(KEYINPUT102), .A3(new_n681), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G119), .ZN(G21));
  XNOR2_X1  g501(.A(new_n509), .B(KEYINPUT103), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n562), .A2(new_n513), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n688), .B1(new_n689), .B2(new_n547), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n578), .B(new_n690), .C1(new_n579), .C2(new_n580), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(KEYINPUT104), .ZN(new_n692));
  OAI21_X1  g506(.A(G472), .B1(new_n584), .B2(G902), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n693), .A2(new_n694), .A3(new_n578), .A4(new_n690), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n463), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n654), .A2(new_n655), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n696), .A2(new_n697), .A3(new_n667), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G122), .ZN(G24));
  NAND4_X1  g515(.A1(new_n693), .A2(new_n660), .A3(new_n622), .A4(new_n690), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n678), .A2(new_n680), .ZN(new_n703));
  OAI21_X1  g517(.A(KEYINPUT105), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n622), .B(new_n690), .C1(new_n579), .C2(new_n580), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n678), .A2(new_n680), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n706), .A2(new_n707), .A3(new_n660), .A4(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n704), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G125), .ZN(G27));
  INV_X1    g525(.A(KEYINPUT106), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n325), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n318), .A2(KEYINPUT106), .A3(new_n323), .A4(new_n324), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n713), .A2(G469), .A3(new_n343), .A4(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(G469), .A2(G902), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n351), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n503), .A2(new_n598), .A3(new_n504), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n506), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n718), .B1(new_n717), .B2(new_n720), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n673), .A2(new_n578), .A3(new_n660), .A4(new_n724), .ZN(new_n725));
  XOR2_X1   g539(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n235), .B1(new_n571), .B2(new_n548), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n728), .A2(KEYINPUT42), .A3(new_n660), .A4(new_n724), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G131), .ZN(G33));
  AOI211_X1 g545(.A(new_n235), .B(new_n723), .C1(new_n560), .C2(new_n571), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n636), .B(KEYINPUT109), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G134), .ZN(G36));
  INV_X1    g549(.A(new_n596), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n588), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(KEYINPUT43), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n616), .A2(new_n738), .A3(new_n626), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(KEYINPUT44), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n719), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(KEYINPUT44), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT110), .ZN(new_n743));
  OR2_X1    g557(.A1(new_n334), .A2(KEYINPUT45), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n713), .A2(KEYINPUT45), .A3(new_n343), .A4(new_n714), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n744), .A2(G469), .A3(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(KEYINPUT46), .A3(new_n716), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n351), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT46), .B1(new_n746), .B2(new_n716), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n507), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n743), .B1(new_n751), .B2(new_n640), .ZN(new_n752));
  INV_X1    g566(.A(new_n751), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(KEYINPUT110), .A3(new_n641), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n741), .A2(new_n742), .A3(new_n752), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(KEYINPUT111), .B(G137), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(G39));
  NAND2_X1  g571(.A1(new_n753), .A2(KEYINPUT47), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT47), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n751), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n673), .A2(new_n578), .A3(new_n719), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n660), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G140), .ZN(G42));
  INV_X1    g578(.A(new_n665), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n737), .B1(KEYINPUT49), .B2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n766), .A2(new_n578), .A3(new_n455), .A4(new_n507), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(KEYINPUT112), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n656), .ZN(new_n769));
  INV_X1    g583(.A(new_n649), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n767), .A2(KEYINPUT112), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n765), .A2(KEYINPUT49), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n769), .A2(new_n770), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT119), .ZN(new_n774));
  INV_X1    g588(.A(new_n719), .ZN(new_n775));
  INV_X1    g589(.A(new_n629), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n738), .A2(new_n776), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n777), .A2(new_n696), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n765), .A2(new_n507), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n775), .B(new_n778), .C1(new_n761), .C2(new_n779), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n777), .A2(new_n665), .A3(new_n720), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n706), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n665), .A2(new_n458), .A3(new_n720), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n770), .A2(new_n578), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT120), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n786), .A2(new_n588), .A3(new_n596), .A4(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n780), .A2(new_n782), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n656), .A2(new_n598), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n777), .A2(new_n667), .A3(new_n696), .A4(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT50), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n774), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n774), .B(KEYINPUT51), .C1(new_n789), .C2(new_n792), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n457), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n786), .A2(new_n597), .A3(new_n787), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n781), .A2(new_n728), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT48), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n778), .A2(new_n708), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n797), .A2(new_n798), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n724), .A2(new_n706), .A3(new_n660), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n803), .B1(new_n732), .B2(new_n733), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n604), .A2(new_n607), .A3(new_n632), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n805), .A2(KEYINPUT114), .A3(new_n719), .ZN(new_n806));
  AOI211_X1 g620(.A(new_n626), .B(new_n806), .C1(new_n560), .C2(new_n571), .ZN(new_n807));
  OAI21_X1  g621(.A(KEYINPUT114), .B1(new_n805), .B2(new_n719), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n577), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT115), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n806), .ZN(new_n811));
  AND4_X1   g625(.A1(KEYINPUT115), .A2(new_n627), .A3(new_n811), .A4(new_n809), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n804), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(KEYINPUT116), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n673), .A2(new_n622), .A3(new_n811), .A4(new_n809), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n627), .A2(KEYINPUT115), .A3(new_n811), .A4(new_n809), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n819), .A2(new_n820), .A3(new_n804), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n814), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n698), .A2(new_n631), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n626), .A2(new_n717), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n649), .A2(new_n507), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n638), .A2(new_n661), .A3(new_n710), .A4(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n654), .A2(new_n655), .A3(new_n697), .ZN(new_n829));
  AOI211_X1 g643(.A(new_n666), .B(new_n829), .C1(new_n692), .C2(new_n695), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n617), .A2(new_n505), .A3(new_n583), .A4(new_n585), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n736), .B(new_n505), .C1(new_n410), .C2(new_n416), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT113), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT113), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n653), .A2(new_n834), .A3(new_n505), .A4(new_n736), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n588), .A2(new_n505), .A3(new_n451), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n833), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  OAI22_X1  g651(.A1(new_n831), .A2(new_n626), .B1(new_n586), .B2(new_n837), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n830), .A2(new_n838), .A3(new_n572), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n671), .A2(new_n668), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n839), .A2(new_n730), .A3(new_n840), .A4(new_n686), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n822), .A2(new_n828), .A3(KEYINPUT53), .A4(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  INV_X1    g661(.A(new_n685), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT102), .B1(new_n627), .B2(new_n681), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n663), .A2(new_n505), .A3(new_n617), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n586), .A2(new_n837), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n700), .A2(new_n851), .A3(new_n623), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n671), .A2(new_n668), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n850), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n819), .A2(new_n820), .A3(new_n804), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n820), .B1(new_n819), .B2(new_n804), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n855), .B(new_n730), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n826), .B(KEYINPUT52), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n847), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n841), .B1(new_n814), .B2(new_n821), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(KEYINPUT117), .A3(KEYINPUT53), .A4(new_n828), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n845), .A2(new_n846), .A3(new_n860), .A4(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n864));
  INV_X1    g678(.A(new_n843), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT53), .B1(new_n861), .B2(new_n828), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT54), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n863), .A2(new_n864), .A3(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n864), .B1(new_n863), .B2(new_n867), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n802), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(G952), .A2(G953), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n773), .B1(new_n872), .B2(new_n873), .ZN(G75));
  NOR2_X1   g688(.A1(new_n319), .A2(G952), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT122), .Z(new_n876));
  NAND3_X1  g690(.A1(new_n845), .A2(new_n860), .A3(new_n862), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(G210), .A3(G902), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT56), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n495), .A2(new_n498), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT121), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT55), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(new_n496), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n880), .A2(new_n884), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n876), .B1(new_n885), .B2(new_n886), .ZN(G51));
  NAND2_X1  g701(.A1(new_n877), .A2(KEYINPUT54), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n863), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n716), .A2(KEYINPUT57), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n716), .A2(KEYINPUT57), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n350), .ZN(new_n893));
  INV_X1    g707(.A(new_n746), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n877), .A2(G902), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n875), .B1(new_n893), .B2(new_n895), .ZN(G54));
  NAND4_X1  g710(.A1(new_n877), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n897));
  INV_X1    g711(.A(new_n404), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n897), .A2(new_n898), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n899), .A2(new_n900), .A3(new_n875), .ZN(G60));
  NOR2_X1   g715(.A1(new_n590), .A2(new_n591), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n868), .A2(new_n870), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n594), .B(KEYINPUT59), .Z(new_n904));
  AOI21_X1  g718(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n889), .A2(new_n902), .A3(new_n904), .ZN(new_n906));
  INV_X1    g720(.A(new_n876), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n905), .A2(new_n908), .ZN(G63));
  NAND2_X1  g723(.A1(G217), .A2(G902), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT60), .Z(new_n911));
  NAND3_X1  g725(.A1(new_n877), .A2(new_n620), .A3(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n877), .A2(new_n911), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n907), .B(new_n912), .C1(new_n913), .C2(new_n226), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT61), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n914), .B(new_n915), .ZN(G66));
  INV_X1    g730(.A(new_n855), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n319), .B1(new_n459), .B2(G224), .ZN(new_n919));
  AOI22_X1  g733(.A1(new_n917), .A2(new_n319), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n920), .B1(new_n918), .B2(new_n919), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n882), .B1(G898), .B2(new_n319), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n921), .B(new_n922), .ZN(G69));
  NAND2_X1  g737(.A1(new_n540), .A2(new_n541), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n394), .A2(new_n395), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n924), .B(new_n925), .Z(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n630), .A2(new_n319), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n755), .A2(new_n763), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n638), .A2(new_n661), .A3(new_n710), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n754), .A2(new_n699), .A3(new_n728), .A4(new_n752), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n931), .A2(new_n932), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n930), .A2(new_n936), .A3(new_n730), .A4(new_n734), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n927), .B(new_n929), .C1(new_n937), .C2(G953), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n933), .A2(new_n658), .A3(new_n935), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT62), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n653), .A2(new_n604), .ZN(new_n943));
  OAI21_X1  g757(.A(KEYINPUT125), .B1(new_n943), .B2(new_n597), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n663), .A2(new_n944), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n943), .A2(new_n597), .A3(KEYINPUT125), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n946), .A2(new_n642), .A3(new_n719), .ZN(new_n947));
  AOI22_X1  g761(.A1(new_n941), .A2(new_n942), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(G953), .B1(new_n948), .B2(new_n930), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n938), .B1(new_n949), .B2(new_n927), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n319), .B1(G227), .B2(G900), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n938), .B2(KEYINPUT126), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n950), .B(new_n952), .Z(G72));
  NAND3_X1  g767(.A1(new_n948), .A2(new_n855), .A3(new_n930), .ZN(new_n954));
  NAND2_X1  g768(.A1(G472), .A2(G902), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT63), .Z(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT127), .Z(new_n957));
  AOI21_X1  g771(.A(new_n645), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n957), .B1(new_n937), .B2(new_n917), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n566), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(G952), .B2(new_n319), .ZN(new_n961));
  AOI211_X1 g775(.A(new_n566), .B(new_n646), .C1(new_n860), .C2(new_n843), .ZN(new_n962));
  AOI211_X1 g776(.A(new_n958), .B(new_n961), .C1(new_n956), .C2(new_n962), .ZN(G57));
endmodule


