//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 1 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 0 1 1 1 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n577, new_n578, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n595, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n642, new_n643, new_n646,
    new_n648, new_n649, new_n650, new_n652, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT66), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  AOI22_X1  g033(.A1(new_n457), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  INV_X1    g034(.A(G137), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(KEYINPUT67), .A3(new_n461), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n470), .B1(G2104), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NOR3_X1   g048(.A1(new_n473), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n474));
  OAI21_X1  g049(.A(G101), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT69), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(G101), .C1(new_n472), .C2(new_n474), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n469), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(KEYINPUT70), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT70), .ZN(new_n481));
  NAND4_X1  g056(.A1(new_n469), .A2(new_n476), .A3(new_n481), .A4(new_n478), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(G113), .A2(G2104), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n462), .A2(new_n463), .ZN(new_n485));
  INV_X1    g060(.A(G125), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G160));
  AND2_X1   g065(.A1(new_n467), .A2(KEYINPUT71), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n467), .A2(KEYINPUT71), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n471), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G136), .ZN(new_n495));
  OAI21_X1  g070(.A(G2105), .B1(new_n491), .B2(new_n492), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G124), .ZN(new_n498));
  OR2_X1    g073(.A1(G100), .A2(G2105), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n500));
  AND3_X1   g075(.A1(new_n495), .A2(new_n498), .A3(new_n500), .ZN(G162));
  AND2_X1   g076(.A1(G126), .A2(G2105), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n502), .B1(new_n462), .B2(new_n463), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT72), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n505), .B(new_n502), .C1(new_n462), .C2(new_n463), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT73), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n471), .A2(G114), .ZN(new_n509));
  OAI21_X1  g084(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OR2_X1    g086(.A1(G102), .A2(G2105), .ZN(new_n512));
  INV_X1    g087(.A(G114), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G2105), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n512), .A2(new_n514), .A3(KEYINPUT73), .A4(G2104), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT74), .A2(KEYINPUT4), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT74), .A2(KEYINPUT4), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(G138), .A3(new_n471), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n517), .B1(new_n485), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n519), .ZN(new_n521));
  INV_X1    g096(.A(new_n517), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(new_n467), .A3(new_n522), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n507), .A2(new_n516), .A3(new_n520), .A4(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(G164));
  INV_X1    g100(.A(G543), .ZN(new_n526));
  AND2_X1   g101(.A1(KEYINPUT75), .A2(G651), .ZN(new_n527));
  NOR2_X1   g102(.A1(KEYINPUT75), .A2(G651), .ZN(new_n528));
  OAI21_X1  g103(.A(KEYINPUT6), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n526), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G50), .ZN(new_n533));
  INV_X1    g108(.A(G88), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n529), .A2(new_n531), .ZN(new_n535));
  XNOR2_X1  g110(.A(KEYINPUT5), .B(G543), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n533), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g113(.A(KEYINPUT75), .B(G651), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n536), .A2(G62), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n541), .A2(KEYINPUT76), .B1(G75), .B2(G543), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT76), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n536), .A2(new_n543), .A3(G62), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n540), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n538), .A2(new_n545), .ZN(G303));
  INV_X1    g121(.A(G303), .ZN(G166));
  NAND3_X1  g122(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT7), .ZN(new_n549));
  INV_X1    g124(.A(G89), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n537), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(KEYINPUT77), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT77), .ZN(new_n553));
  OAI211_X1 g128(.A(new_n553), .B(new_n549), .C1(new_n537), .C2(new_n550), .ZN(new_n554));
  AND2_X1   g129(.A1(G63), .A2(G651), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n532), .A2(G51), .B1(new_n536), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n552), .A2(new_n554), .A3(new_n556), .ZN(G286));
  INV_X1    g132(.A(G286), .ZN(G168));
  AOI22_X1  g133(.A1(new_n536), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n559), .A2(new_n540), .ZN(new_n560));
  AND2_X1   g135(.A1(KEYINPUT5), .A2(G543), .ZN(new_n561));
  NOR2_X1   g136(.A1(KEYINPUT5), .A2(G543), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n563), .B1(new_n529), .B2(new_n531), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G90), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n532), .A2(G52), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n560), .A2(new_n565), .A3(new_n566), .ZN(G301));
  INV_X1    g142(.A(G301), .ZN(G171));
  AOI22_X1  g143(.A1(new_n536), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n569), .A2(new_n540), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n564), .A2(G81), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n532), .A2(G43), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G860), .ZN(G153));
  NAND4_X1  g150(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g151(.A1(G1), .A2(G3), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT8), .ZN(new_n578));
  NAND4_X1  g153(.A1(G319), .A2(G483), .A3(G661), .A4(new_n578), .ZN(G188));
  NAND2_X1  g154(.A1(new_n532), .A2(G53), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT9), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT78), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g158(.A(KEYINPUT79), .B1(new_n580), .B2(KEYINPUT9), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT9), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n532), .A2(new_n585), .A3(new_n586), .A4(G53), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n580), .A2(KEYINPUT78), .A3(KEYINPUT9), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n583), .A2(new_n584), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n536), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT80), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(G651), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(new_n590), .B2(new_n591), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n592), .A2(new_n594), .B1(G91), .B2(new_n564), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n589), .A2(new_n595), .ZN(G299));
  INV_X1    g171(.A(KEYINPUT82), .ZN(new_n597));
  NAND2_X1  g172(.A1(G49), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(KEYINPUT81), .B1(new_n535), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT81), .ZN(new_n601));
  AOI211_X1 g176(.A(new_n601), .B(new_n598), .C1(new_n529), .C2(new_n531), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(G74), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n593), .B1(new_n563), .B2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G87), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n537), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n597), .B1(new_n603), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n605), .B1(new_n564), .B2(G87), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n610), .B(KEYINPUT82), .C1(new_n600), .C2(new_n602), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(G288));
  NAND2_X1  g188(.A1(G73), .A2(G543), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT83), .ZN(new_n615));
  INV_X1    g190(.A(G61), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(new_n563), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n617), .A2(new_n539), .B1(new_n564), .B2(G86), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n619));
  AND2_X1   g194(.A1(G48), .A2(G543), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n535), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n619), .B1(new_n535), .B2(new_n620), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n618), .B1(new_n622), .B2(new_n623), .ZN(G305));
  AOI22_X1  g199(.A1(G47), .A2(new_n532), .B1(new_n564), .B2(G85), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT85), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n536), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n627), .A2(new_n540), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n628), .ZN(G290));
  NAND2_X1  g204(.A1(G301), .A2(G868), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n564), .A2(G92), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT10), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(G79), .A2(G543), .ZN(new_n634));
  INV_X1    g209(.A(G66), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n563), .B2(new_n635), .ZN(new_n636));
  AOI22_X1  g211(.A1(new_n532), .A2(G54), .B1(new_n636), .B2(G651), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n630), .B1(new_n639), .B2(G868), .ZN(G284));
  OAI21_X1  g215(.A(new_n630), .B1(new_n639), .B2(G868), .ZN(G321));
  NAND2_X1  g216(.A1(G286), .A2(G868), .ZN(new_n642));
  INV_X1    g217(.A(G299), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n642), .B1(new_n643), .B2(G868), .ZN(G297));
  OAI21_X1  g219(.A(new_n642), .B1(new_n643), .B2(G868), .ZN(G280));
  INV_X1    g220(.A(G559), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n639), .B1(new_n646), .B2(G860), .ZN(G148));
  NOR2_X1   g222(.A1(new_n574), .A2(G868), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n639), .A2(new_n646), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n648), .B1(new_n649), .B2(G868), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT86), .ZN(G323));
  XNOR2_X1  g226(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n652));
  XNOR2_X1  g227(.A(G323), .B(new_n652), .ZN(G282));
  OR2_X1    g228(.A1(new_n472), .A2(new_n474), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(new_n467), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT12), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT13), .ZN(new_n657));
  INV_X1    g232(.A(G2100), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT88), .Z(new_n660));
  OAI21_X1  g235(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n661));
  INV_X1    g236(.A(G111), .ZN(new_n662));
  AOI22_X1  g237(.A1(new_n661), .A2(KEYINPUT89), .B1(new_n662), .B2(G2105), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n663), .B1(KEYINPUT89), .B2(new_n661), .ZN(new_n664));
  INV_X1    g239(.A(G135), .ZN(new_n665));
  INV_X1    g240(.A(G123), .ZN(new_n666));
  OAI221_X1 g241(.A(new_n664), .B1(new_n493), .B2(new_n665), .C1(new_n666), .C2(new_n496), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(G2096), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n667), .A2(G2096), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n657), .A2(new_n658), .ZN(new_n670));
  NAND4_X1  g245(.A1(new_n660), .A2(new_n668), .A3(new_n669), .A4(new_n670), .ZN(G156));
  XNOR2_X1  g246(.A(G2451), .B(G2454), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT16), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1341), .B(G1348), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n673), .B(new_n674), .Z(new_n675));
  INV_X1    g250(.A(KEYINPUT14), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2427), .B(G2438), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2430), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT15), .B(G2435), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n676), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(new_n679), .B2(new_n678), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n675), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2443), .B(G2446), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g260(.A(G14), .B1(new_n682), .B2(new_n684), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(G401));
  XNOR2_X1  g262(.A(G2072), .B(G2078), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT90), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT91), .B(KEYINPUT17), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G2067), .B(G2678), .ZN(new_n692));
  XOR2_X1   g267(.A(G2084), .B(G2090), .Z(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  NOR3_X1   g269(.A1(new_n691), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT92), .Z(new_n696));
  NAND3_X1  g271(.A1(new_n689), .A2(new_n692), .A3(new_n693), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT18), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n691), .A2(new_n692), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n689), .A2(new_n692), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n700), .A2(new_n693), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n698), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n696), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G2096), .B(G2100), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT93), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n703), .B(new_n705), .ZN(G227));
  XNOR2_X1  g281(.A(G1971), .B(G1976), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT19), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XOR2_X1   g284(.A(G1956), .B(G2474), .Z(new_n710));
  XOR2_X1   g285(.A(G1961), .B(G1966), .Z(new_n711));
  AND2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT20), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n710), .A2(new_n711), .ZN(new_n715));
  NOR3_X1   g290(.A1(new_n709), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n709), .B2(new_n715), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT94), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT94), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n718), .B(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n720), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g301(.A(G1991), .B(G1996), .Z(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(G1981), .B(G1986), .ZN(new_n729));
  INV_X1    g304(.A(new_n727), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n721), .A2(new_n725), .A3(new_n730), .ZN(new_n731));
  AND3_X1   g306(.A1(new_n728), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n729), .B1(new_n728), .B2(new_n731), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(new_n733), .ZN(G229));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G35), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G162), .B2(new_n735), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT29), .B(G2090), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(KEYINPUT103), .B1(new_n667), .B2(new_n735), .ZN(new_n740));
  NOR3_X1   g315(.A1(new_n667), .A2(KEYINPUT103), .A3(new_n735), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n735), .A2(G27), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G164), .B2(new_n735), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n741), .B1(G2078), .B2(new_n743), .ZN(new_n744));
  AND3_X1   g319(.A1(new_n739), .A2(new_n740), .A3(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G16), .ZN(new_n746));
  NOR2_X1   g321(.A1(G171), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G5), .B2(new_n746), .ZN(new_n748));
  INV_X1    g323(.A(G1961), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(KEYINPUT105), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n735), .A2(G32), .ZN(new_n752));
  NAND3_X1  g327(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT26), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n654), .A2(G105), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(G141), .ZN(new_n758));
  INV_X1    g333(.A(G129), .ZN(new_n759));
  OAI221_X1 g334(.A(new_n757), .B1(new_n493), .B2(new_n758), .C1(new_n759), .C2(new_n496), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n752), .B1(new_n761), .B2(new_n735), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT27), .B(G1996), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n751), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n735), .A2(G26), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT28), .Z(new_n768));
  OR2_X1    g343(.A1(new_n471), .A2(G116), .ZN(new_n769));
  OAI21_X1  g344(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n497), .A2(G128), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n494), .A2(G140), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n768), .B1(new_n774), .B2(G29), .ZN(new_n775));
  INV_X1    g350(.A(G2067), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(KEYINPUT105), .B2(new_n750), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n574), .A2(G16), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G16), .B2(G19), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT100), .B(G1341), .Z(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n748), .A2(new_n749), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n780), .A2(new_n782), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT30), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n785), .A2(G28), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n735), .B1(new_n785), .B2(G28), .ZN(new_n787));
  AND2_X1   g362(.A1(KEYINPUT31), .A2(G11), .ZN(new_n788));
  NOR2_X1   g363(.A1(KEYINPUT31), .A2(G11), .ZN(new_n789));
  OAI22_X1  g364(.A1(new_n786), .A2(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n743), .ZN(new_n791));
  INV_X1    g366(.A(G2078), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AND3_X1   g368(.A1(new_n783), .A2(new_n784), .A3(new_n793), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n745), .A2(new_n766), .A3(new_n778), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n746), .A2(G4), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n639), .B2(new_n746), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT99), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT98), .B(G1348), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(new_n471), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT25), .Z(new_n805));
  INV_X1    g380(.A(G139), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n493), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n807), .A2(KEYINPUT101), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n807), .A2(KEYINPUT101), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n803), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT102), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI211_X1 g387(.A(KEYINPUT102), .B(new_n803), .C1(new_n808), .C2(new_n809), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n735), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n735), .A2(G33), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(G2072), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n746), .A2(G20), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT23), .Z(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(G299), .B2(G16), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G1956), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n817), .A2(new_n821), .ZN(new_n822));
  NOR3_X1   g397(.A1(new_n814), .A2(G2072), .A3(new_n816), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n746), .A2(G21), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(G168), .B2(new_n746), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n826), .A2(G1966), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT104), .Z(new_n828));
  INV_X1    g403(.A(KEYINPUT24), .ZN(new_n829));
  INV_X1    g404(.A(G34), .ZN(new_n830));
  AOI21_X1  g405(.A(G29), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(new_n829), .B2(new_n830), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(G160), .B2(new_n735), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n833), .A2(G2084), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n833), .A2(G2084), .B1(new_n826), .B2(G1966), .ZN(new_n835));
  AND3_X1   g410(.A1(new_n828), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n801), .A2(new_n824), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(G16), .A2(G23), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT96), .Z(new_n839));
  OR2_X1    g414(.A1(new_n600), .A2(new_n602), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(new_n610), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n839), .B1(new_n841), .B2(new_n746), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT97), .Z(new_n843));
  XOR2_X1   g418(.A(KEYINPUT33), .B(G1976), .Z(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n746), .A2(G22), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(G166), .B2(new_n746), .ZN(new_n848));
  INV_X1    g423(.A(G1971), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  MUX2_X1   g425(.A(G6), .B(G305), .S(G16), .Z(new_n851));
  XOR2_X1   g426(.A(KEYINPUT32), .B(G1981), .Z(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  AND3_X1   g428(.A1(new_n846), .A2(new_n850), .A3(new_n853), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n843), .A2(new_n845), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(KEYINPUT34), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n735), .A2(G25), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n497), .A2(G119), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT95), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n863));
  INV_X1    g438(.A(G107), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n863), .B1(new_n864), .B2(G2105), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n865), .B1(new_n494), .B2(G131), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n859), .B1(new_n867), .B2(G29), .ZN(new_n868));
  XOR2_X1   g443(.A(KEYINPUT35), .B(G1991), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n746), .A2(G24), .ZN(new_n871));
  INV_X1    g446(.A(G290), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n871), .B1(new_n872), .B2(new_n746), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n873), .A2(G1986), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n873), .A2(G1986), .ZN(new_n875));
  NOR3_X1   g450(.A1(new_n870), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(new_n856), .B2(KEYINPUT34), .ZN(new_n877));
  OAI21_X1  g452(.A(KEYINPUT36), .B1(new_n858), .B2(new_n877), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n856), .A2(KEYINPUT34), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT36), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n879), .A2(new_n880), .A3(new_n857), .A4(new_n876), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n837), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT106), .ZN(G311));
  INV_X1    g458(.A(new_n882), .ZN(G150));
  NAND2_X1  g459(.A1(new_n639), .A2(G559), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(KEYINPUT38), .Z(new_n886));
  NAND2_X1  g461(.A1(G80), .A2(G543), .ZN(new_n887));
  INV_X1    g462(.A(G67), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n887), .B1(new_n563), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT107), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n539), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n891), .B1(new_n890), .B2(new_n889), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n532), .A2(G55), .ZN(new_n893));
  INV_X1    g468(.A(G93), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n893), .B1(new_n894), .B2(new_n537), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(new_n574), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n573), .B1(new_n892), .B2(new_n895), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n886), .B(new_n899), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n900), .A2(KEYINPUT39), .ZN(new_n901));
  INV_X1    g476(.A(G860), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(KEYINPUT39), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n896), .A2(new_n902), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT37), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n906), .ZN(G145));
  XOR2_X1   g482(.A(new_n489), .B(new_n667), .Z(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(G162), .ZN(new_n909));
  INV_X1    g484(.A(new_n656), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n867), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n862), .A2(new_n656), .A3(new_n866), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n812), .A2(new_n813), .A3(new_n761), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n761), .B1(new_n812), .B2(new_n813), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n911), .B(new_n912), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n774), .B(G164), .ZN(new_n917));
  OAI21_X1  g492(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n918));
  INV_X1    g493(.A(G118), .ZN(new_n919));
  AOI22_X1  g494(.A1(new_n918), .A2(KEYINPUT108), .B1(new_n919), .B2(G2105), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(KEYINPUT108), .B2(new_n918), .ZN(new_n921));
  INV_X1    g496(.A(G142), .ZN(new_n922));
  INV_X1    g497(.A(G130), .ZN(new_n923));
  OAI221_X1 g498(.A(new_n921), .B1(new_n493), .B2(new_n922), .C1(new_n923), .C2(new_n496), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n917), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n917), .A2(new_n924), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n915), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n911), .A2(new_n912), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(new_n929), .A3(new_n913), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n916), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n927), .B1(new_n916), .B2(new_n930), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n909), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n916), .A2(new_n930), .ZN(new_n935));
  INV_X1    g510(.A(new_n927), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n909), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n937), .A2(new_n938), .A3(new_n931), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n934), .A2(new_n939), .ZN(new_n940));
  XOR2_X1   g515(.A(KEYINPUT109), .B(G37), .Z(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g518(.A1(new_n872), .A2(G303), .ZN(new_n944));
  NAND2_X1  g519(.A1(G290), .A2(G166), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n841), .B(G305), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n944), .A2(new_n947), .A3(new_n945), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(KEYINPUT42), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n643), .A2(KEYINPUT110), .A3(new_n638), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT110), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(G299), .B2(new_n639), .ZN(new_n955));
  NAND2_X1  g530(.A1(G299), .A2(new_n639), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  XOR2_X1   g533(.A(new_n649), .B(new_n899), .Z(new_n959));
  OR2_X1    g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n957), .A2(KEYINPUT41), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT41), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n953), .A2(new_n955), .A3(new_n962), .A4(new_n956), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n959), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n952), .A2(new_n960), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n952), .B1(new_n960), .B2(new_n964), .ZN(new_n966));
  OAI21_X1  g541(.A(G868), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT111), .ZN(new_n968));
  OR2_X1    g543(.A1(new_n896), .A2(G868), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n968), .B1(new_n967), .B2(new_n969), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(G295));
  NAND2_X1  g547(.A1(new_n967), .A2(new_n969), .ZN(G331));
  NAND2_X1  g548(.A1(G168), .A2(G171), .ZN(new_n974));
  NAND2_X1  g549(.A1(G286), .A2(G301), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n899), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n974), .A2(new_n898), .A3(new_n897), .A4(new_n975), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(new_n978), .A3(KEYINPUT112), .ZN(new_n979));
  INV_X1    g554(.A(new_n899), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n980), .A2(new_n981), .A3(new_n975), .A4(new_n974), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n957), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n977), .A2(new_n978), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n961), .A2(new_n963), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n984), .A2(new_n986), .A3(new_n951), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n987), .A2(new_n941), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT43), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n961), .A2(new_n963), .A3(new_n979), .A4(new_n982), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n957), .A2(new_n977), .A3(new_n978), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n951), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n992), .A2(KEYINPUT113), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n994));
  AOI211_X1 g569(.A(new_n994), .B(new_n951), .C1(new_n990), .C2(new_n991), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n988), .B(new_n989), .C1(new_n993), .C2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G37), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n987), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n951), .B1(new_n984), .B2(new_n986), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT43), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1001), .A2(KEYINPUT44), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n993), .A2(new_n995), .ZN(new_n1003));
  INV_X1    g578(.A(new_n988), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT43), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n998), .ZN(new_n1006));
  INV_X1    g581(.A(new_n999), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1006), .A2(new_n989), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT114), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1006), .A2(new_n1007), .A3(KEYINPUT114), .A4(new_n989), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1005), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1002), .B1(KEYINPUT44), .B2(new_n1012), .ZN(G397));
  AND2_X1   g588(.A1(new_n488), .A2(G40), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n480), .A2(new_n482), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT115), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1384), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n516), .A2(new_n523), .A3(new_n520), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n505), .B1(new_n467), .B2(new_n502), .ZN(new_n1020));
  INV_X1    g595(.A(new_n506), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1018), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n480), .A2(KEYINPUT115), .A3(new_n482), .A4(new_n1014), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1017), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n840), .A2(G1976), .A3(new_n610), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1026), .A2(G8), .A3(new_n1027), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n1028), .A2(KEYINPUT52), .ZN(new_n1029));
  INV_X1    g604(.A(G1976), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n609), .A2(new_n1030), .A3(new_n611), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1033), .A2(new_n1026), .A3(G8), .A4(new_n1027), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT49), .ZN(new_n1035));
  NOR2_X1   g610(.A1(G305), .A2(G1981), .ZN(new_n1036));
  INV_X1    g611(.A(G1981), .ZN(new_n1037));
  INV_X1    g612(.A(new_n623), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n621), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1037), .B1(new_n1039), .B2(new_n618), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1035), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(G305), .A2(G1981), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1039), .A2(new_n1037), .A3(new_n618), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1042), .A2(KEYINPUT49), .A3(new_n1043), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1026), .A2(G8), .A3(new_n1041), .A4(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1034), .A2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT119), .B1(new_n1029), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1028), .A2(KEYINPUT52), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT119), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1048), .A2(new_n1049), .A3(new_n1034), .A4(new_n1045), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1047), .A2(new_n1050), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n1017), .A2(new_n1025), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT50), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1053), .B(new_n1018), .C1(new_n1019), .C2(new_n1022), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT117), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1023), .A2(KEYINPUT50), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1023), .A2(KEYINPUT117), .A3(KEYINPUT50), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G2084), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1052), .A2(new_n1059), .A3(KEYINPUT121), .A4(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT121), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1017), .A2(new_n1057), .A3(new_n1025), .A4(new_n1058), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1062), .B1(new_n1063), .B2(G2084), .ZN(new_n1064));
  OAI211_X1 g639(.A(KEYINPUT45), .B(new_n1018), .C1(new_n1019), .C2(new_n1022), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT45), .B1(new_n524), .B2(new_n1018), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1017), .A2(new_n1025), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G1966), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1061), .A2(new_n1064), .A3(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1072), .A2(G8), .A3(G168), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(G303), .A2(G8), .ZN(new_n1075));
  XNOR2_X1  g650(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1017), .A2(new_n1025), .A3(new_n1068), .ZN(new_n1078));
  OAI22_X1  g653(.A1(new_n1078), .A2(G1971), .B1(new_n1063), .B2(G2090), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G8), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1077), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  XOR2_X1   g657(.A(new_n1075), .B(new_n1076), .Z(new_n1083));
  NAND3_X1  g658(.A1(new_n1079), .A2(new_n1083), .A3(G8), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1084), .A2(KEYINPUT63), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1051), .A2(new_n1074), .A3(new_n1082), .A4(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT63), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1054), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1053), .B1(new_n524), .B2(new_n1018), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1017), .A2(new_n1025), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G2090), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1091), .A2(new_n1092), .B1(new_n1069), .B2(new_n849), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1077), .B1(new_n1093), .B2(new_n1081), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n1034), .A2(new_n1045), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1094), .A2(new_n1084), .A3(new_n1048), .A4(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1087), .B1(new_n1096), .B2(new_n1073), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1086), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1084), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1026), .A2(G8), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n612), .A2(new_n1030), .ZN(new_n1101));
  XOR2_X1   g676(.A(new_n1101), .B(KEYINPUT120), .Z(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n1045), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1100), .B1(new_n1103), .B2(new_n1043), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1099), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1098), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1072), .A2(G8), .ZN(new_n1109));
  NOR2_X1   g684(.A1(G168), .A2(new_n1081), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT51), .B1(new_n1111), .B2(KEYINPUT125), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1109), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1114));
  OAI211_X1 g689(.A(G8), .B(new_n1112), .C1(new_n1072), .C2(G286), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1072), .A2(new_n1110), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT62), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT62), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1114), .A2(new_n1119), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT53), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1121), .A2(G2078), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1078), .A2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1017), .A2(new_n1068), .A3(new_n792), .A4(new_n1025), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n1121), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1063), .A2(new_n749), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1123), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(G171), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1096), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1118), .A2(new_n1120), .A3(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1068), .A2(new_n483), .A3(new_n1014), .A4(new_n1122), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1125), .A2(new_n1126), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(G171), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1121), .A2(new_n1124), .B1(new_n1063), .B2(new_n749), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1134), .A2(G301), .A3(new_n1123), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1133), .A2(new_n1135), .A3(KEYINPUT54), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1136), .A2(new_n1096), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT126), .B1(new_n1132), .B2(G171), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1134), .A2(new_n1139), .A3(G301), .A4(new_n1131), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1138), .A2(new_n1128), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT54), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1137), .A2(new_n1117), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT57), .ZN(new_n1145));
  AOI211_X1 g720(.A(KEYINPUT123), .B(new_n1145), .C1(new_n589), .C2(new_n595), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(KEYINPUT123), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT123), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT57), .ZN(new_n1149));
  AND4_X1   g724(.A1(new_n589), .A2(new_n595), .A3(new_n1147), .A4(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1146), .A2(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(KEYINPUT56), .B(G2072), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1078), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(G1956), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1017), .A2(new_n1025), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1090), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1154), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1151), .B1(new_n1153), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(G1348), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1063), .A2(new_n1159), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1017), .A2(new_n776), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n638), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1151), .A2(new_n1153), .A3(new_n1157), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1158), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(KEYINPUT60), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1160), .A2(KEYINPUT60), .A3(new_n1161), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(KEYINPUT124), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(new_n639), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1166), .A2(KEYINPUT124), .A3(new_n638), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OR2_X1    g745(.A1(new_n1166), .A2(KEYINPUT124), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1165), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1163), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1173), .B1(new_n1174), .B2(new_n1158), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1153), .A2(new_n1157), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1151), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1178), .A2(KEYINPUT61), .A3(new_n1163), .ZN(new_n1179));
  INV_X1    g754(.A(G1996), .ZN(new_n1180));
  XOR2_X1   g755(.A(KEYINPUT58), .B(G1341), .Z(new_n1181));
  AOI22_X1  g756(.A1(new_n1078), .A2(new_n1180), .B1(new_n1026), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT59), .ZN(new_n1183));
  OR3_X1    g758(.A1(new_n1182), .A2(new_n1183), .A3(new_n573), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1183), .B1(new_n1182), .B2(new_n573), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1175), .A2(new_n1179), .A3(new_n1184), .A4(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1164), .B1(new_n1172), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1144), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1098), .A2(KEYINPUT122), .A3(new_n1105), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1108), .A2(new_n1130), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  NOR3_X1   g765(.A1(new_n1155), .A2(KEYINPUT45), .A3(new_n1024), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n867), .B(new_n869), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n774), .A2(G2067), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n772), .A2(new_n776), .A3(new_n773), .ZN(new_n1194));
  AND2_X1   g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n760), .B(new_n1180), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(G1986), .ZN(new_n1199));
  OAI211_X1 g774(.A(new_n1192), .B(new_n1198), .C1(new_n1199), .C2(new_n872), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n872), .A2(new_n1199), .ZN(new_n1201));
  XOR2_X1   g776(.A(new_n1201), .B(KEYINPUT116), .Z(new_n1202));
  OAI21_X1  g777(.A(new_n1191), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1190), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g779(.A(new_n1195), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1191), .B1(new_n1205), .B2(new_n760), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1191), .A2(new_n1180), .ZN(new_n1207));
  AND2_X1   g782(.A1(new_n1207), .A2(KEYINPUT46), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n1207), .A2(KEYINPUT46), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1206), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  XOR2_X1   g785(.A(new_n1210), .B(KEYINPUT47), .Z(new_n1211));
  AND2_X1   g786(.A1(new_n1202), .A2(new_n1191), .ZN(new_n1212));
  OR2_X1    g787(.A1(new_n1212), .A2(KEYINPUT48), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1192), .A2(new_n1198), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1214), .A2(new_n1191), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1212), .A2(KEYINPUT48), .ZN(new_n1216));
  AND3_X1   g791(.A1(new_n1213), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n862), .A2(new_n869), .A3(new_n866), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1194), .B1(new_n1197), .B2(new_n1218), .ZN(new_n1219));
  AOI211_X1 g794(.A(new_n1211), .B(new_n1217), .C1(new_n1191), .C2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1204), .A2(new_n1220), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g796(.A(G319), .B1(new_n685), .B2(new_n686), .ZN(new_n1223));
  NOR2_X1   g797(.A1(G227), .A2(new_n1223), .ZN(new_n1224));
  OAI21_X1  g798(.A(new_n1224), .B1(new_n732), .B2(new_n733), .ZN(new_n1225));
  AOI21_X1  g799(.A(new_n1225), .B1(new_n940), .B2(new_n941), .ZN(new_n1226));
  INV_X1    g800(.A(KEYINPUT127), .ZN(new_n1227));
  AND3_X1   g801(.A1(new_n1001), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  AOI21_X1  g802(.A(new_n1227), .B1(new_n1001), .B2(new_n1226), .ZN(new_n1229));
  NOR2_X1   g803(.A1(new_n1228), .A2(new_n1229), .ZN(G308));
  NAND2_X1  g804(.A1(new_n1001), .A2(new_n1226), .ZN(G225));
endmodule


