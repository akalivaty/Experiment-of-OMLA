//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 1 0 0 1 1 1 0 0 1 1 1 1 0 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 1 0 1 0 1 0 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981;
  XOR2_X1   g000(.A(G116), .B(G119), .Z(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT2), .B(G113), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT3), .B1(new_n190), .B2(G107), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G104), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n190), .A2(G107), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT4), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(G101), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n197), .B1(new_n196), .B2(G101), .ZN(new_n199));
  INV_X1    g013(.A(G101), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT80), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT80), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G101), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n204), .A2(new_n194), .A3(new_n195), .A4(new_n191), .ZN(new_n205));
  AND3_X1   g019(.A1(new_n199), .A2(KEYINPUT81), .A3(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(KEYINPUT81), .B1(new_n199), .B2(new_n205), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n189), .B(new_n198), .C1(new_n206), .C2(new_n207), .ZN(new_n208));
  XOR2_X1   g022(.A(G110), .B(G122), .Z(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT5), .ZN(new_n211));
  INV_X1    g025(.A(G119), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(G116), .ZN(new_n213));
  OAI211_X1 g027(.A(G113), .B(new_n213), .C1(new_n187), .C2(new_n211), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n214), .B1(new_n188), .B2(new_n187), .ZN(new_n215));
  INV_X1    g029(.A(new_n195), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n190), .A2(G107), .ZN(new_n217));
  OAI21_X1  g031(.A(G101), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n205), .A2(new_n218), .ZN(new_n219));
  OR2_X1    g033(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n208), .A2(new_n210), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT87), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n208), .A2(KEYINPUT87), .A3(new_n210), .A4(new_n220), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n210), .B1(new_n208), .B2(new_n220), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT86), .ZN(new_n227));
  OR2_X1    g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT6), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n229), .B1(new_n226), .B2(new_n227), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n225), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n226), .A2(new_n229), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT88), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT88), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n226), .A2(new_n234), .A3(new_n229), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G143), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT65), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G143), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G146), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n237), .A2(G146), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n242), .A2(G128), .A3(new_n244), .A4(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(G128), .B1(new_n245), .B2(new_n243), .ZN(new_n247));
  INV_X1    g061(.A(G146), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n238), .A2(new_n240), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n237), .A2(G146), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n246), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT90), .B1(new_n253), .B2(G125), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT90), .ZN(new_n255));
  INV_X1    g069(.A(G125), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n246), .A2(new_n252), .A3(new_n255), .A4(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT0), .ZN(new_n259));
  INV_X1    g073(.A(G128), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(KEYINPUT0), .A2(G128), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT64), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n262), .B(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n251), .A2(new_n261), .A3(new_n264), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n242), .A2(KEYINPUT0), .A3(G128), .A4(new_n244), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G125), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT89), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n267), .A2(KEYINPUT89), .A3(G125), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n258), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G224), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(G953), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n272), .B(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n231), .A2(new_n236), .A3(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G902), .ZN(new_n277));
  INV_X1    g091(.A(new_n274), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT91), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n258), .A2(new_n270), .A3(new_n271), .A4(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT7), .B1(new_n278), .B2(KEYINPUT91), .ZN(new_n281));
  OR3_X1    g095(.A1(new_n280), .A2(KEYINPUT92), .A3(new_n281), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n258), .A2(new_n268), .B1(KEYINPUT7), .B2(new_n278), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n283), .B1(new_n223), .B2(new_n224), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n215), .B(new_n219), .ZN(new_n285));
  XOR2_X1   g099(.A(new_n209), .B(KEYINPUT8), .Z(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT92), .B1(new_n280), .B2(new_n281), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n282), .A2(new_n284), .A3(new_n287), .A4(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n276), .A2(new_n277), .A3(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(G210), .B1(G237), .B2(G902), .ZN(new_n291));
  XOR2_X1   g105(.A(new_n291), .B(KEYINPUT93), .Z(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(G214), .B1(G237), .B2(G902), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n276), .A2(new_n277), .A3(new_n292), .A4(new_n289), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  XOR2_X1   g111(.A(KEYINPUT9), .B(G234), .Z(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G217), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n299), .A2(new_n300), .A3(G953), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n241), .A2(G128), .ZN(new_n302));
  INV_X1    g116(.A(G134), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n302), .B(new_n303), .C1(G128), .C2(new_n237), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT65), .B(G143), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n305), .A2(new_n260), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n237), .A2(G128), .ZN(new_n307));
  OAI21_X1  g121(.A(G134), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G122), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n309), .A2(G116), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT102), .B(G122), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n310), .B1(new_n311), .B2(G116), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n304), .A2(new_n308), .B1(new_n312), .B2(new_n193), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(G116), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT14), .B1(new_n309), .B2(G116), .ZN(new_n315));
  OR3_X1    g129(.A1(new_n309), .A2(KEYINPUT14), .A3(G116), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G107), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT103), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT103), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n317), .A2(new_n320), .A3(G107), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n313), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT13), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n306), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n302), .B1(G128), .B2(new_n237), .ZN(new_n325));
  OAI211_X1 g139(.A(G134), .B(new_n324), .C1(new_n325), .C2(new_n323), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n312), .B(new_n193), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(new_n304), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n301), .B1(new_n322), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n322), .A2(new_n328), .A3(new_n301), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n277), .ZN(new_n333));
  INV_X1    g147(.A(G478), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(KEYINPUT15), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n333), .B(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(G234), .A2(G237), .ZN(new_n338));
  INV_X1    g152(.A(G953), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n338), .A2(G952), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(G902), .A3(G953), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(KEYINPUT104), .ZN(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT21), .B(G898), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n340), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n337), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT20), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT100), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n347), .A2(KEYINPUT100), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT94), .ZN(new_n351));
  INV_X1    g165(.A(G214), .ZN(new_n352));
  NOR3_X1   g166(.A1(new_n352), .A2(G237), .A3(G953), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n351), .B1(new_n305), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G237), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(new_n339), .A3(G214), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n241), .A2(KEYINPUT94), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n353), .A2(G143), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n354), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G131), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT17), .ZN(new_n361));
  INV_X1    g175(.A(G131), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n354), .A2(new_n357), .A3(new_n362), .A4(new_n358), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n360), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT99), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(G125), .B(G140), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT16), .ZN(new_n368));
  OR3_X1    g182(.A1(new_n256), .A2(KEYINPUT16), .A3(G140), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n248), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(G146), .A3(new_n369), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n359), .A2(KEYINPUT17), .A3(G131), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n360), .A2(KEYINPUT99), .A3(new_n361), .A4(new_n363), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n366), .A2(new_n374), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(G113), .B(G122), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n378), .B(new_n190), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n359), .A2(KEYINPUT18), .A3(G131), .ZN(new_n380));
  NAND2_X1  g194(.A1(KEYINPUT18), .A2(G131), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n354), .A2(new_n357), .A3(new_n381), .A4(new_n358), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n367), .B(new_n248), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT95), .B1(new_n380), .B2(new_n384), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n382), .A2(new_n383), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT95), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n359), .A2(KEYINPUT18), .A3(G131), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n377), .A2(new_n379), .A3(new_n390), .ZN(new_n391));
  XOR2_X1   g205(.A(KEYINPUT96), .B(KEYINPUT19), .Z(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n367), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT97), .ZN(new_n394));
  INV_X1    g208(.A(new_n367), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT19), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT97), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n392), .A2(new_n397), .A3(new_n367), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n394), .A2(new_n248), .A3(new_n396), .A4(new_n398), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n399), .A2(new_n372), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n360), .A2(new_n363), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n385), .A2(new_n389), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT98), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n400), .A2(new_n401), .ZN(new_n405));
  NOR3_X1   g219(.A1(new_n380), .A2(KEYINPUT95), .A3(new_n384), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n387), .B1(new_n386), .B2(new_n388), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n379), .B1(new_n408), .B2(KEYINPUT98), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n391), .B1(new_n404), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(G475), .A2(G902), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n348), .B(new_n350), .C1(new_n410), .C2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n377), .A2(new_n390), .ZN(new_n414));
  INV_X1    g228(.A(new_n379), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(KEYINPUT101), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n377), .A2(new_n379), .A3(new_n390), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT101), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n379), .B1(new_n377), .B2(new_n390), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n277), .B(new_n416), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G475), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n415), .B1(new_n402), .B2(new_n403), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n408), .A2(KEYINPUT98), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n417), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(new_n349), .A3(new_n411), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n413), .A2(new_n422), .A3(new_n426), .ZN(new_n427));
  NOR3_X1   g241(.A1(new_n297), .A2(new_n346), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n300), .B1(G234), .B2(new_n277), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n367), .A2(new_n248), .ZN(new_n431));
  OAI21_X1  g245(.A(KEYINPUT73), .B1(new_n212), .B2(G128), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT23), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n212), .A2(G128), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT23), .ZN(new_n435));
  OAI211_X1 g249(.A(KEYINPUT73), .B(new_n435), .C1(new_n212), .C2(G128), .ZN(new_n436));
  XNOR2_X1  g250(.A(KEYINPUT74), .B(G110), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n433), .A2(new_n434), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT75), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n438), .B(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n212), .A2(G128), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT72), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n441), .B1(new_n442), .B2(new_n434), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n443), .B1(new_n442), .B2(new_n434), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT24), .B(G110), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n372), .B(new_n431), .C1(new_n440), .C2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n433), .A2(new_n434), .A3(new_n436), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G110), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n373), .B(new_n449), .C1(new_n445), .C2(new_n444), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n339), .A2(G221), .A3(G234), .ZN(new_n452));
  INV_X1    g266(.A(G137), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n452), .B(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(KEYINPUT76), .B(KEYINPUT22), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n452), .B(G137), .ZN(new_n457));
  INV_X1    g271(.A(new_n455), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n456), .A2(new_n459), .A3(KEYINPUT77), .ZN(new_n460));
  AOI21_X1  g274(.A(KEYINPUT77), .B1(new_n456), .B2(new_n459), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n451), .A2(new_n463), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n456), .A2(new_n459), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n447), .A2(new_n450), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n464), .A2(new_n277), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT25), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n464), .A2(KEYINPUT25), .A3(new_n277), .A4(new_n466), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n430), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n429), .A2(G902), .ZN(new_n472));
  XOR2_X1   g286(.A(new_n472), .B(KEYINPUT78), .Z(new_n473));
  AND3_X1   g287(.A1(new_n447), .A2(new_n450), .A3(new_n465), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n462), .B1(new_n447), .B2(new_n450), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n471), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(G472), .A2(G902), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT66), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n480), .B1(new_n303), .B2(G137), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT11), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n453), .A2(G134), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT11), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n480), .B(new_n485), .C1(new_n303), .C2(G137), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n482), .A2(new_n362), .A3(new_n484), .A4(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n303), .A2(G137), .ZN(new_n488));
  OAI21_X1  g302(.A(G131), .B1(new_n483), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT67), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n487), .A2(KEYINPUT67), .A3(new_n489), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n253), .A3(new_n493), .ZN(new_n494));
  AOI211_X1 g308(.A(new_n260), .B(new_n243), .C1(new_n241), .C2(G146), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n249), .A2(new_n250), .B1(new_n259), .B2(new_n260), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n495), .A2(KEYINPUT0), .B1(new_n496), .B2(new_n264), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G131), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n487), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT30), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n494), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n487), .A2(new_n489), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n253), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n502), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n189), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT31), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n501), .A2(new_n505), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(new_n189), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT26), .B(G101), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n355), .A2(new_n339), .A3(G210), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n507), .A2(new_n508), .A3(new_n511), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n494), .A2(new_n501), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n189), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT28), .ZN(new_n521));
  INV_X1    g335(.A(new_n189), .ZN(new_n522));
  AND4_X1   g336(.A1(new_n521), .A2(new_n501), .A3(new_n522), .A4(new_n505), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n497), .A2(new_n500), .B1(new_n253), .B2(new_n504), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n521), .B1(new_n524), .B2(new_n522), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n520), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT70), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n516), .B(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n518), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n494), .A2(new_n501), .A3(new_n502), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n532), .B1(new_n502), .B2(new_n524), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n510), .B1(new_n533), .B2(new_n189), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n508), .B1(new_n534), .B2(new_n517), .ZN(new_n535));
  OAI211_X1 g349(.A(KEYINPUT32), .B(new_n479), .C1(new_n531), .C2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n507), .A2(new_n511), .A3(new_n517), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT31), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(new_n518), .A3(new_n530), .ZN(new_n540));
  AOI21_X1  g354(.A(KEYINPUT32), .B1(new_n540), .B2(new_n479), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n534), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n516), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT71), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT29), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n528), .B(new_n520), .C1(new_n525), .C2(new_n523), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n544), .A2(new_n545), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n547), .B(new_n546), .C1(new_n534), .C2(new_n517), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT71), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n509), .A2(new_n189), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n551), .B1(new_n523), .B2(new_n525), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(new_n516), .ZN(new_n553));
  AOI21_X1  g367(.A(G902), .B1(new_n553), .B2(KEYINPUT29), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n548), .A2(new_n550), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(G472), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n478), .B1(new_n542), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(G221), .B1(new_n299), .B2(G902), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n500), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n196), .A2(G101), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(new_n205), .A3(KEYINPUT4), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT81), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n199), .A2(KEYINPUT81), .A3(new_n205), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n265), .A2(new_n266), .A3(new_n198), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n219), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT10), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n570), .B1(new_n246), .B2(new_n252), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n566), .A2(new_n568), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  OAI211_X1 g386(.A(G128), .B(new_n244), .C1(new_n305), .C2(new_n248), .ZN(new_n573));
  INV_X1    g387(.A(new_n245), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT82), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n243), .B1(new_n241), .B2(G146), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT82), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n576), .A2(new_n577), .A3(G128), .A4(new_n245), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n244), .B1(new_n305), .B2(new_n248), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT1), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n580), .B1(new_n305), .B2(new_n248), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n579), .B1(new_n581), .B2(new_n260), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n575), .A2(new_n578), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n569), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n570), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n560), .B1(new_n572), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(KEYINPUT10), .B1(new_n583), .B2(new_n569), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n567), .B1(new_n564), .B2(new_n565), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n253), .A2(KEYINPUT10), .A3(new_n569), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(KEYINPUT83), .B1(new_n591), .B2(new_n560), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n572), .A2(new_n585), .A3(KEYINPUT83), .A4(new_n560), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n587), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(G110), .B(G140), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n339), .A2(G227), .ZN(new_n597));
  XOR2_X1   g411(.A(new_n596), .B(new_n597), .Z(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n595), .A2(KEYINPUT85), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT85), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n572), .A2(new_n585), .A3(new_n560), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT83), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n586), .B1(new_n604), .B2(new_n593), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n601), .B1(new_n605), .B2(new_n598), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n599), .B1(new_n604), .B2(new_n593), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n246), .A2(new_n219), .A3(new_n252), .ZN(new_n608));
  OR2_X1    g422(.A1(new_n608), .A2(KEYINPUT84), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(KEYINPUT84), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(new_n584), .A3(new_n610), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n611), .A2(KEYINPUT12), .A3(new_n500), .ZN(new_n612));
  AOI21_X1  g426(.A(KEYINPUT12), .B1(new_n611), .B2(new_n500), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n607), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n600), .A2(new_n606), .A3(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(G469), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n616), .A3(new_n277), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n277), .ZN(new_n618));
  OAI22_X1  g432(.A1(new_n592), .A2(new_n594), .B1(new_n612), .B2(new_n613), .ZN(new_n619));
  XOR2_X1   g433(.A(new_n598), .B(KEYINPUT79), .Z(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  AOI22_X1  g435(.A1(new_n619), .A2(new_n621), .B1(new_n607), .B2(new_n587), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n618), .B1(new_n622), .B2(G469), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n559), .B1(new_n617), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n428), .A2(new_n557), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(new_n625), .B(new_n204), .Z(G3));
  NAND2_X1  g440(.A1(new_n540), .A2(new_n277), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(G472), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n540), .A2(new_n479), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(new_n478), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n631), .A2(new_n624), .ZN(new_n632));
  INV_X1    g446(.A(new_n297), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT105), .ZN(new_n634));
  OAI21_X1  g448(.A(KEYINPUT33), .B1(new_n301), .B2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n331), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n635), .B1(new_n636), .B2(new_n329), .ZN(new_n637));
  INV_X1    g451(.A(new_n635), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n330), .A2(new_n331), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n637), .A2(new_n639), .A3(new_n277), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(G478), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n332), .A2(new_n334), .A3(new_n277), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(KEYINPUT106), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT106), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n641), .A2(new_n645), .A3(new_n642), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n427), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n648), .A2(new_n344), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n632), .A2(new_n633), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  NAND2_X1  g466(.A1(new_n408), .A2(KEYINPUT98), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(new_n404), .A3(new_n415), .ZN(new_n654));
  AOI211_X1 g468(.A(new_n350), .B(new_n412), .C1(new_n654), .C2(new_n417), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n350), .A2(new_n348), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n656), .B1(new_n425), .B2(new_n411), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT107), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n422), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n421), .A2(KEYINPUT107), .A3(G475), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n658), .A2(new_n660), .A3(new_n336), .A4(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n344), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n632), .A2(new_n633), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G107), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT108), .B(KEYINPUT35), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G9));
  INV_X1    g481(.A(new_n630), .ZN(new_n668));
  AOI21_X1  g482(.A(KEYINPUT25), .B1(new_n476), .B2(new_n277), .ZN(new_n669));
  INV_X1    g483(.A(new_n470), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n429), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT36), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n462), .A2(new_n672), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n451), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n451), .A2(new_n673), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n674), .A2(new_n473), .A3(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n671), .A2(new_n676), .A3(KEYINPUT109), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT109), .ZN(new_n678));
  INV_X1    g492(.A(new_n676), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n678), .B1(new_n471), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n428), .A2(new_n624), .A3(new_n668), .A4(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT37), .B(G110), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G12));
  INV_X1    g499(.A(G900), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n340), .B1(new_n342), .B2(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n662), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n681), .B1(new_n542), .B2(new_n556), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n688), .A2(new_n689), .A3(new_n624), .A4(new_n633), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G128), .ZN(G30));
  NAND2_X1  g505(.A1(new_n294), .A2(new_n296), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT38), .ZN(new_n693));
  INV_X1    g507(.A(new_n538), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n528), .B1(new_n511), .B2(new_n551), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n277), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n696), .A2(G472), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n537), .A2(new_n697), .A3(new_n541), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n427), .A2(new_n295), .A3(new_n336), .ZN(new_n699));
  NOR4_X1   g513(.A1(new_n693), .A2(new_n682), .A3(new_n698), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n687), .B(KEYINPUT39), .ZN(new_n701));
  AOI211_X1 g515(.A(new_n559), .B(new_n701), .C1(new_n617), .C2(new_n623), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n702), .A2(KEYINPUT40), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(KEYINPUT40), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n700), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n241), .B(KEYINPUT110), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G45));
  INV_X1    g521(.A(new_n687), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n647), .A2(new_n427), .A3(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n709), .A2(new_n689), .A3(new_n624), .A4(new_n633), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G146), .ZN(G48));
  AND3_X1   g525(.A1(new_n615), .A2(new_n616), .A3(new_n277), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n616), .B1(new_n615), .B2(new_n277), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n712), .A2(new_n713), .A3(new_n559), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n649), .A2(new_n714), .A3(new_n557), .A4(new_n633), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT41), .B(G113), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G15));
  NAND4_X1  g531(.A1(new_n714), .A2(new_n557), .A3(new_n663), .A4(new_n633), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G116), .ZN(G18));
  NOR2_X1   g533(.A1(new_n346), .A2(new_n427), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n714), .A2(new_n633), .A3(new_n720), .A4(new_n689), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G119), .ZN(G21));
  NAND2_X1  g536(.A1(new_n552), .A2(new_n529), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n518), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n479), .B1(new_n724), .B2(new_n535), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT111), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT111), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n727), .B(new_n479), .C1(new_n724), .C2(new_n535), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  AND4_X1   g543(.A1(new_n477), .A2(new_n729), .A3(new_n345), .A4(new_n628), .ZN(new_n730));
  INV_X1    g544(.A(new_n427), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n337), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n714), .A2(new_n730), .A3(new_n633), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G122), .ZN(G24));
  NAND3_X1  g548(.A1(new_n539), .A2(new_n518), .A3(new_n723), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n727), .B1(new_n735), .B2(new_n479), .ZN(new_n736));
  INV_X1    g550(.A(new_n728), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n628), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n738), .A2(new_n681), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n714), .A2(new_n739), .A3(new_n709), .A4(new_n633), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G125), .ZN(G27));
  NAND2_X1  g555(.A1(new_n617), .A2(new_n623), .ZN(new_n742));
  INV_X1    g556(.A(new_n295), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n743), .B1(new_n294), .B2(new_n296), .ZN(new_n744));
  AND4_X1   g558(.A1(KEYINPUT112), .A2(new_n742), .A3(new_n744), .A4(new_n558), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT112), .B1(new_n624), .B2(new_n744), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(KEYINPUT113), .A2(KEYINPUT42), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n747), .A2(new_n557), .A3(new_n709), .A4(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n742), .A2(new_n744), .A3(new_n558), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT112), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n624), .A2(KEYINPUT112), .A3(new_n744), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n753), .A2(new_n557), .A3(new_n709), .A4(new_n754), .ZN(new_n755));
  XOR2_X1   g569(.A(KEYINPUT113), .B(KEYINPUT42), .Z(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n750), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G131), .ZN(G33));
  AND4_X1   g574(.A1(new_n557), .A2(new_n753), .A3(new_n688), .A4(new_n754), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(new_n303), .ZN(G36));
  OR2_X1    g576(.A1(new_n622), .A2(KEYINPUT45), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n622), .A2(KEYINPUT45), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(G469), .A3(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n618), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(KEYINPUT46), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n617), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT46), .B1(new_n765), .B2(new_n766), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n558), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n770), .A2(new_n701), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT114), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n731), .A2(new_n647), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT43), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(new_n630), .A3(new_n682), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(KEYINPUT44), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n744), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n772), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(new_n453), .ZN(G39));
  XOR2_X1   g594(.A(new_n770), .B(KEYINPUT47), .Z(new_n781));
  INV_X1    g595(.A(new_n744), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n647), .A2(new_n427), .A3(new_n708), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n782), .A2(new_n783), .A3(new_n477), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n781), .A2(new_n542), .A3(new_n556), .A4(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G140), .ZN(G42));
  AOI22_X1  g600(.A1(new_n726), .A2(new_n728), .B1(new_n627), .B2(G472), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n477), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n775), .A2(new_n340), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT117), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n775), .A2(new_n791), .A3(new_n340), .ZN(new_n792));
  AOI211_X1 g606(.A(new_n295), .B(new_n788), .C1(new_n790), .C2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(new_n693), .A3(new_n714), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n793), .A2(KEYINPUT50), .A3(new_n693), .A4(new_n714), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n714), .A2(new_n744), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n799), .B1(new_n790), .B2(new_n792), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n739), .ZN(new_n801));
  INV_X1    g615(.A(new_n799), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(new_n477), .A3(new_n340), .A4(new_n698), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n803), .A2(new_n427), .A3(new_n647), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n798), .A2(new_n801), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n788), .B1(new_n790), .B2(new_n792), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n712), .A2(new_n713), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n558), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n744), .B(new_n807), .C1(new_n781), .C2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT118), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n806), .B(new_n810), .C1(new_n811), .C2(KEYINPUT51), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n798), .A2(new_n811), .A3(new_n801), .A4(new_n805), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n798), .A2(new_n801), .A3(new_n805), .A4(new_n810), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n800), .A2(new_n557), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT48), .ZN(new_n819));
  OAI211_X1 g633(.A(G952), .B(new_n339), .C1(new_n803), .C2(new_n648), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n714), .A2(new_n633), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n820), .B1(new_n807), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT119), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n715), .A2(new_n733), .A3(new_n718), .A4(new_n721), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n542), .A2(new_n556), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n828), .A2(new_n658), .A3(new_n660), .A4(new_n661), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n624), .A2(new_n682), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n337), .A2(new_n708), .ZN(new_n831));
  NOR4_X1   g645(.A1(new_n829), .A2(new_n830), .A3(new_n782), .A4(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n827), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n761), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n658), .A2(new_n422), .A3(new_n336), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n344), .B1(new_n648), .B2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n836), .A2(new_n624), .A3(new_n633), .A4(new_n631), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n683), .A3(new_n625), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n783), .A2(new_n738), .A3(new_n681), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n753), .A2(new_n839), .A3(new_n754), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n759), .A2(new_n833), .A3(new_n834), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n671), .A2(new_n676), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n698), .A2(new_n699), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n692), .ZN(new_n845));
  AOI211_X1 g659(.A(new_n559), .B(new_n687), .C1(new_n617), .C2(new_n623), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n847), .A2(new_n690), .A3(new_n740), .A4(new_n710), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(KEYINPUT52), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n826), .B1(new_n842), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n740), .A2(new_n690), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT116), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT52), .ZN(new_n853));
  NOR4_X1   g667(.A1(new_n698), .A2(new_n699), .A3(new_n692), .A4(new_n843), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n853), .B1(new_n854), .B2(new_n846), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n740), .A2(new_n690), .A3(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n852), .A2(new_n710), .A3(new_n855), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n848), .A2(new_n853), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n753), .A2(new_n839), .A3(new_n754), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(new_n625), .A3(new_n683), .A4(new_n837), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n862), .B1(new_n758), .B2(new_n750), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n827), .A2(new_n761), .A3(new_n832), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n860), .A2(KEYINPUT53), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n850), .A2(new_n865), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n866), .A2(KEYINPUT54), .ZN(new_n867));
  INV_X1    g681(.A(new_n842), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT53), .B1(new_n868), .B2(new_n860), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n842), .A2(new_n849), .A3(new_n826), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT54), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n819), .A2(KEYINPUT119), .A3(new_n822), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n825), .A2(new_n867), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  OAI22_X1  g687(.A1(new_n817), .A2(new_n873), .B1(G952), .B2(G953), .ZN(new_n874));
  OR2_X1    g688(.A1(new_n808), .A2(KEYINPUT49), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n808), .A2(KEYINPUT49), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n875), .A2(new_n558), .A3(new_n295), .A4(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n693), .A2(new_n731), .A3(new_n647), .ZN(new_n878));
  INV_X1    g692(.A(new_n698), .ZN(new_n879));
  NOR4_X1   g693(.A1(new_n877), .A2(new_n878), .A3(new_n478), .A4(new_n879), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT115), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n874), .A2(new_n881), .ZN(G75));
  AOI21_X1  g696(.A(new_n277), .B1(new_n850), .B2(new_n865), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT56), .B1(new_n883), .B2(new_n292), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n231), .A2(new_n236), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(new_n275), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT55), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n884), .B(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n339), .A2(G952), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(G51));
  XNOR2_X1  g704(.A(new_n866), .B(KEYINPUT54), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n766), .A2(KEYINPUT57), .ZN(new_n892));
  OR2_X1    g706(.A1(new_n766), .A2(KEYINPUT57), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n615), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n883), .A2(G469), .A3(new_n763), .A4(new_n764), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n889), .B1(new_n895), .B2(new_n896), .ZN(G54));
  AND3_X1   g711(.A1(new_n883), .A2(KEYINPUT58), .A3(G475), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n898), .A2(new_n425), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n899), .A2(KEYINPUT120), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n899), .A2(KEYINPUT120), .ZN(new_n901));
  INV_X1    g715(.A(new_n889), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n902), .B1(new_n898), .B2(new_n425), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n900), .A2(new_n901), .A3(new_n903), .ZN(G60));
  NAND2_X1  g718(.A1(G478), .A2(G902), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT59), .Z(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n637), .A2(new_n639), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT121), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n891), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n906), .B1(new_n867), .B2(new_n871), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n910), .B(new_n902), .C1(new_n911), .C2(new_n909), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(G63));
  NAND2_X1  g727(.A1(G217), .A2(G902), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT60), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n866), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(KEYINPUT122), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n866), .A2(new_n919), .A3(new_n916), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n674), .A2(new_n675), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT123), .Z(new_n923));
  AOI21_X1  g737(.A(new_n889), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n925));
  INV_X1    g739(.A(new_n476), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n918), .A2(new_n926), .A3(new_n920), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n924), .A2(KEYINPUT124), .A3(new_n925), .A4(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n919), .B1(new_n866), .B2(new_n916), .ZN(new_n929));
  AOI211_X1 g743(.A(KEYINPUT122), .B(new_n915), .C1(new_n850), .C2(new_n865), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n923), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n927), .A2(new_n931), .A3(new_n902), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n925), .A2(KEYINPUT124), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n925), .A2(KEYINPUT124), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n928), .A2(new_n935), .ZN(G66));
  OAI21_X1  g750(.A(G953), .B1(new_n343), .B2(new_n273), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n827), .A2(new_n838), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n937), .B1(new_n938), .B2(G953), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n885), .B1(G898), .B2(new_n339), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(G69));
  AND3_X1   g755(.A1(new_n852), .A2(new_n710), .A3(new_n857), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n705), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT62), .ZN(new_n944));
  INV_X1    g758(.A(new_n785), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n648), .A2(new_n835), .ZN(new_n946));
  INV_X1    g760(.A(new_n557), .ZN(new_n947));
  NOR4_X1   g761(.A1(new_n946), .A2(new_n947), .A3(new_n751), .A4(new_n701), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT125), .Z(new_n949));
  NOR4_X1   g763(.A1(new_n944), .A2(new_n779), .A3(new_n945), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n339), .ZN(new_n951));
  NAND3_X1  g765(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n394), .A2(new_n396), .A3(new_n398), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n533), .B(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n951), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n954), .ZN(new_n956));
  INV_X1    g770(.A(new_n772), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n557), .A2(new_n295), .A3(new_n845), .A4(new_n732), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n778), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n834), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n785), .A2(new_n759), .A3(new_n942), .ZN(new_n962));
  OAI21_X1  g776(.A(KEYINPUT126), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n962), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT126), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n964), .A2(new_n965), .A3(new_n834), .A4(new_n960), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n956), .B1(new_n967), .B2(G953), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n686), .A2(new_n339), .A3(G227), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n955), .B1(new_n968), .B2(new_n969), .ZN(G72));
  XNOR2_X1  g784(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n971));
  NAND2_X1  g785(.A1(G472), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n544), .A2(new_n538), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n973), .B(new_n974), .C1(new_n869), .C2(new_n870), .ZN(new_n975));
  INV_X1    g789(.A(new_n973), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n950), .B2(new_n938), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n543), .A2(new_n517), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n902), .B(new_n975), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n963), .A2(new_n938), .A3(new_n966), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n543), .B1(new_n980), .B2(new_n973), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n979), .B1(new_n516), .B2(new_n981), .ZN(G57));
endmodule


