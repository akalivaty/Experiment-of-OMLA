//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 1 1 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n207));
  INV_X1    g0007(.A(G87), .ZN(new_n208));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(G226), .ZN(new_n214));
  INV_X1    g0014(.A(G77), .ZN(new_n215));
  INV_X1    g0015(.A(G244), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n213), .B1(new_n202), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n206), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  OAI21_X1  g0019(.A(G50), .B1(G58), .B2(G68), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT64), .Z(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  OR3_X1    g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n206), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT0), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n219), .A2(new_n224), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n218), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G226), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT65), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n234), .B(new_n238), .Z(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NOR2_X1   g0046(.A1(G20), .A2(G33), .ZN(new_n247));
  AOI22_X1  g0047(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT8), .B(G58), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n222), .A2(G33), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n223), .B1(new_n206), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G13), .ZN(new_n255));
  NOR3_X1   g0055(.A1(new_n255), .A2(new_n222), .A3(G1), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(new_n253), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n202), .B1(new_n258), .B2(G20), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n257), .A2(new_n259), .B1(new_n202), .B2(new_n256), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT9), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT67), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n263), .B(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G190), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT3), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(G223), .A3(G1698), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G222), .ZN(new_n274));
  OAI221_X1 g0074(.A(new_n271), .B1(new_n215), .B2(new_n270), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n258), .B1(G41), .B2(G45), .ZN(new_n278));
  INV_X1    g0078(.A(G274), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n276), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n278), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n280), .B1(new_n283), .B2(G226), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n277), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n265), .B1(new_n266), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(G200), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n287), .B1(new_n262), .B2(new_n261), .ZN(new_n288));
  OR3_X1    g0088(.A1(new_n286), .A2(KEYINPUT10), .A3(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(KEYINPUT10), .B1(new_n286), .B2(new_n288), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G179), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n285), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n293), .B1(G169), .B2(new_n285), .ZN(new_n294));
  INV_X1    g0094(.A(new_n261), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n256), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT66), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT66), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n256), .A2(new_n301), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  AOI211_X1 g0103(.A(new_n253), .B(new_n303), .C1(new_n258), .C2(G20), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G68), .ZN(new_n305));
  INV_X1    g0105(.A(new_n247), .ZN(new_n306));
  OAI22_X1  g0106(.A1(new_n306), .A2(new_n202), .B1(new_n222), .B2(G68), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n250), .A2(new_n215), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n253), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT11), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  NOR3_X1   g0111(.A1(new_n299), .A2(KEYINPUT12), .A3(G68), .ZN(new_n312));
  INV_X1    g0112(.A(G68), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n303), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n312), .B1(new_n314), .B2(KEYINPUT12), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT13), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n270), .A2(G232), .A3(G1698), .ZN(new_n319));
  NAND2_X1  g0119(.A1(G33), .A2(G97), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n319), .B(new_n320), .C1(new_n273), .C2(new_n214), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n276), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n280), .B1(new_n283), .B2(G238), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n318), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n322), .A2(new_n318), .A3(new_n323), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G169), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n328), .A2(KEYINPUT68), .A3(KEYINPUT14), .ZN(new_n329));
  INV_X1    g0129(.A(new_n326), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(new_n324), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G179), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(KEYINPUT68), .A2(KEYINPUT14), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(KEYINPUT68), .A2(KEYINPUT14), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n335), .B1(new_n328), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n317), .B1(new_n333), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n331), .A2(new_n266), .ZN(new_n340));
  INV_X1    g0140(.A(G200), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n327), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n316), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n304), .A2(G77), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n303), .A2(new_n215), .ZN(new_n347));
  INV_X1    g0147(.A(new_n253), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G20), .A2(G77), .ZN(new_n349));
  XNOR2_X1  g0149(.A(KEYINPUT15), .B(G87), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n349), .B1(new_n350), .B2(new_n250), .ZN(new_n351));
  INV_X1    g0151(.A(new_n249), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n351), .B1(new_n247), .B2(new_n352), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n346), .B(new_n347), .C1(new_n348), .C2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n270), .A2(G238), .A3(G1698), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n270), .A2(G232), .A3(new_n272), .ZN(new_n356));
  INV_X1    g0156(.A(G107), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n355), .B(new_n356), .C1(new_n357), .C2(new_n270), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n276), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n280), .B1(new_n283), .B2(G244), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n361), .A2(G190), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n362), .B1(new_n341), .B2(new_n361), .ZN(new_n363));
  OR2_X1    g0163(.A1(new_n354), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n361), .A2(G169), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n292), .B2(new_n361), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n354), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NOR3_X1   g0168(.A1(new_n298), .A2(new_n345), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT16), .ZN(new_n370));
  INV_X1    g0170(.A(G58), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n371), .A2(new_n313), .ZN(new_n372));
  OAI21_X1  g0172(.A(G20), .B1(new_n372), .B2(new_n201), .ZN(new_n373));
  INV_X1    g0173(.A(G159), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n373), .B1(new_n374), .B2(new_n306), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n375), .B(KEYINPUT72), .ZN(new_n376));
  INV_X1    g0176(.A(new_n270), .ZN(new_n377));
  NOR2_X1   g0177(.A1(KEYINPUT7), .A2(G20), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT69), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n252), .ZN(new_n381));
  NAND2_X1  g0181(.A1(KEYINPUT69), .A2(G33), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n267), .ZN(new_n384));
  AOI21_X1  g0184(.A(G20), .B1(new_n384), .B2(new_n269), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  OAI211_X1 g0186(.A(G68), .B(new_n379), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT73), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n376), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AND2_X1   g0189(.A1(KEYINPUT69), .A2(G33), .ZN(new_n390));
  NOR2_X1   g0190(.A1(KEYINPUT69), .A2(G33), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n269), .B1(new_n392), .B2(KEYINPUT3), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n222), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n394), .A2(KEYINPUT7), .B1(new_n378), .B2(new_n377), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT73), .B1(new_n395), .B2(G68), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n370), .B1(new_n389), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n381), .A2(KEYINPUT3), .A3(new_n382), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n398), .A2(KEYINPUT70), .A3(new_n268), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT70), .B1(new_n398), .B2(new_n268), .ZN(new_n400));
  INV_X1    g0200(.A(new_n378), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(G20), .B1(new_n398), .B2(new_n268), .ZN(new_n403));
  OAI21_X1  g0203(.A(G68), .B1(new_n403), .B2(new_n386), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT71), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT70), .ZN(new_n406));
  NOR3_X1   g0206(.A1(new_n390), .A2(new_n391), .A3(new_n267), .ZN(new_n407));
  INV_X1    g0207(.A(new_n268), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n398), .A2(KEYINPUT70), .A3(new_n268), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(new_n378), .A3(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT71), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n408), .B1(new_n392), .B2(KEYINPUT3), .ZN(new_n413));
  OAI21_X1  g0213(.A(KEYINPUT7), .B1(new_n413), .B2(G20), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n411), .A2(new_n412), .A3(G68), .A4(new_n414), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n405), .A2(KEYINPUT16), .A3(new_n376), .A4(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n397), .A2(new_n416), .A3(new_n253), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n282), .A2(new_n233), .B1(new_n279), .B2(new_n278), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n272), .A2(G223), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n214), .B2(new_n272), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n398), .A2(new_n421), .A3(new_n268), .ZN(new_n422));
  NAND2_X1  g0222(.A1(G33), .A2(G87), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n281), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n341), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(G190), .B2(new_n426), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n249), .B1(new_n258), .B2(G20), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n429), .A2(new_n257), .B1(new_n256), .B2(new_n249), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n417), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  XNOR2_X1  g0231(.A(new_n431), .B(KEYINPUT17), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT18), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n417), .A2(new_n430), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT74), .ZN(new_n435));
  OAI21_X1  g0235(.A(G169), .B1(new_n418), .B2(new_n424), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n418), .A2(new_n424), .A3(new_n292), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n435), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n436), .B(KEYINPUT74), .C1(new_n426), .C2(new_n292), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n433), .B1(new_n434), .B2(new_n442), .ZN(new_n443));
  AOI211_X1 g0243(.A(KEYINPUT18), .B(new_n441), .C1(new_n417), .C2(new_n430), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n432), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n369), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n413), .A2(new_n222), .A3(G87), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT22), .ZN(new_n450));
  NOR3_X1   g0250(.A1(new_n208), .A2(KEYINPUT22), .A3(G20), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n270), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT80), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n270), .A2(KEYINPUT80), .A3(new_n451), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n450), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n383), .A2(new_n222), .A3(G116), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n357), .A2(G20), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT23), .ZN(new_n460));
  XNOR2_X1  g0260(.A(new_n459), .B(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n457), .A2(KEYINPUT24), .A3(new_n458), .A4(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT24), .ZN(new_n463));
  AOI22_X1  g0263(.A1(KEYINPUT22), .A2(new_n449), .B1(new_n454), .B2(new_n455), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n461), .A2(new_n458), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n462), .A2(new_n466), .A3(new_n253), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n257), .B1(G1), .B2(new_n252), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G107), .ZN(new_n470));
  INV_X1    g0270(.A(new_n459), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n255), .A2(G1), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n471), .A2(KEYINPUT25), .A3(new_n472), .ZN(new_n473));
  OR2_X1    g0273(.A1(new_n473), .A2(KEYINPUT81), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT25), .B1(new_n471), .B2(new_n472), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n473), .B1(new_n475), .B2(KEYINPUT81), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  AND2_X1   g0277(.A1(new_n470), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n467), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(G45), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(G1), .ZN(new_n481));
  AND2_X1   g0281(.A1(KEYINPUT5), .A2(G41), .ZN(new_n482));
  NOR2_X1   g0282(.A1(KEYINPUT5), .A2(G41), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n281), .A2(new_n484), .A3(G264), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G257), .A2(G1698), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(new_n209), .B2(G1698), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n413), .A2(new_n487), .B1(G294), .B2(new_n383), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n485), .B1(new_n488), .B2(new_n281), .ZN(new_n489));
  OR2_X1    g0289(.A1(new_n484), .A2(new_n279), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NOR3_X1   g0291(.A1(new_n489), .A2(G190), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT82), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n485), .B(KEYINPUT82), .C1(new_n488), .C2(new_n281), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n494), .A2(new_n490), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n492), .B1(new_n496), .B2(new_n341), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n479), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n494), .A2(G179), .A3(new_n490), .A4(new_n495), .ZN(new_n499));
  OAI21_X1  g0299(.A(G169), .B1(new_n489), .B2(new_n491), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT83), .ZN(new_n502));
  XNOR2_X1  g0302(.A(new_n501), .B(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n498), .B1(new_n503), .B2(new_n479), .ZN(new_n504));
  OR2_X1    g0304(.A1(new_n210), .A2(KEYINPUT6), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n210), .A2(new_n357), .A3(KEYINPUT6), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OR2_X1    g0307(.A1(KEYINPUT75), .A2(G107), .ZN(new_n508));
  NAND2_X1  g0308(.A1(KEYINPUT75), .A2(G107), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n505), .A2(new_n506), .A3(new_n508), .A4(new_n509), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n511), .A2(G20), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n247), .A2(G77), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g0315(.A(G107), .B(new_n379), .C1(new_n385), .C2(new_n386), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n348), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n256), .A2(G97), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n518), .B1(new_n468), .B2(G97), .ZN(new_n519));
  OAI21_X1  g0319(.A(KEYINPUT76), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT76), .ZN(new_n521));
  INV_X1    g0321(.A(new_n519), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n513), .A2(new_n514), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n523), .B1(new_n395), .B2(G107), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n521), .B(new_n522), .C1(new_n524), .C2(new_n348), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n398), .A2(G244), .A3(new_n272), .A4(new_n268), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT4), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n527), .A2(new_n216), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n529), .A2(new_n272), .A3(new_n268), .A4(new_n269), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n268), .A2(new_n269), .A3(G250), .A4(G1698), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G33), .A2(G283), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n281), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n281), .A2(new_n484), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n490), .B1(new_n211), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n341), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n536), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n528), .A2(new_n533), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n538), .B1(new_n539), .B2(new_n281), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n537), .B1(new_n540), .B2(G190), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n520), .A2(new_n525), .A3(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n398), .A2(G244), .A3(G1698), .A4(new_n268), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n398), .A2(G238), .A3(new_n272), .A4(new_n268), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n383), .A2(G116), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT78), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT78), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n543), .A2(new_n544), .A3(new_n548), .A4(new_n545), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n276), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n481), .A2(G274), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n209), .B2(new_n481), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n281), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT77), .ZN(new_n554));
  XNOR2_X1  g0354(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n550), .A2(new_n292), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n413), .A2(new_n222), .A3(G68), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT19), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n222), .B1(new_n320), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n208), .A2(new_n210), .A3(new_n357), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n222), .A2(G33), .A3(G97), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n559), .A2(new_n560), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n253), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n303), .A2(new_n350), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n564), .B(new_n565), .C1(new_n350), .C2(new_n468), .ZN(new_n566));
  XNOR2_X1  g0366(.A(new_n553), .B(KEYINPUT77), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n549), .A2(new_n276), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n567), .B1(new_n547), .B2(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n556), .B(new_n566), .C1(new_n569), .C2(G169), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n550), .A2(G190), .A3(new_n555), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n469), .A2(G87), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n564), .A2(new_n572), .A3(new_n565), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n571), .B(new_n573), .C1(new_n569), .C2(new_n341), .ZN(new_n574));
  INV_X1    g0374(.A(G169), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n540), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n538), .B(new_n292), .C1(new_n539), .C2(new_n281), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n576), .B(new_n577), .C1(new_n517), .C2(new_n519), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n542), .A2(new_n570), .A3(new_n574), .A4(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(G264), .A2(G1698), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n211), .B2(G1698), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n413), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n377), .A2(G303), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n281), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(G270), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n490), .B1(new_n586), .B2(new_n535), .ZN(new_n587));
  OR2_X1    g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n588), .A2(G190), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(new_n341), .B2(new_n588), .ZN(new_n590));
  INV_X1    g0390(.A(G116), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n253), .B1(new_n300), .B2(new_n302), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n591), .B1(new_n258), .B2(G33), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n591), .A2(new_n303), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n532), .B(new_n222), .C1(G33), .C2(new_n210), .ZN(new_n595));
  XNOR2_X1  g0395(.A(new_n595), .B(KEYINPUT79), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n348), .B1(G20), .B2(new_n591), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n596), .A2(new_n597), .A3(KEYINPUT20), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT20), .B1(new_n596), .B2(new_n597), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n594), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OR2_X1    g0401(.A1(new_n590), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n601), .A2(new_n588), .A3(G169), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT21), .ZN(new_n604));
  OAI211_X1 g0404(.A(KEYINPUT21), .B(G169), .C1(new_n585), .C2(new_n587), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n588), .B2(new_n292), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n603), .A2(new_n604), .B1(new_n606), .B2(new_n601), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  AND4_X1   g0409(.A1(new_n448), .A2(new_n504), .A3(new_n580), .A4(new_n609), .ZN(G372));
  NAND3_X1  g0410(.A1(new_n344), .A2(new_n354), .A3(new_n366), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n339), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n432), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n445), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n291), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n615), .A2(KEYINPUT85), .A3(new_n297), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT85), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n613), .A2(new_n445), .B1(new_n290), .B2(new_n289), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n617), .B1(new_n618), .B2(new_n296), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n570), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n579), .A2(new_n498), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n479), .A2(new_n501), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n607), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n621), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n570), .A2(new_n574), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n576), .A2(new_n577), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n517), .A2(new_n519), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n626), .A2(KEYINPUT84), .A3(KEYINPUT26), .A4(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n629), .A2(new_n570), .A3(new_n574), .A4(KEYINPUT26), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT84), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT26), .ZN(new_n634));
  INV_X1    g0434(.A(new_n520), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n517), .A2(KEYINPUT76), .A3(new_n519), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n577), .B(new_n576), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n570), .A2(new_n574), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n634), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n630), .A2(new_n633), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n625), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n448), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n620), .A2(new_n642), .ZN(G369));
  INV_X1    g0443(.A(new_n601), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n472), .A2(new_n222), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n645), .A2(KEYINPUT27), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(KEYINPUT27), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(G213), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(G343), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n608), .B1(new_n644), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n607), .A2(new_n601), .A3(new_n650), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n655), .A2(G330), .ZN(new_n656));
  INV_X1    g0456(.A(new_n479), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n504), .B1(new_n657), .B2(new_n651), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n503), .A2(new_n479), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n658), .B1(new_n659), .B2(new_n651), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n607), .A2(new_n650), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n479), .A2(new_n501), .A3(new_n651), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n661), .A2(new_n665), .ZN(G399));
  INV_X1    g0466(.A(new_n225), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(G41), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NOR4_X1   g0469(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(G1), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n220), .B2(new_n669), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT28), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n494), .A2(new_n495), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n588), .A2(new_n292), .ZN(new_n675));
  INV_X1    g0475(.A(new_n540), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n674), .A2(new_n675), .A3(new_n569), .A4(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT30), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n496), .A2(new_n540), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n588), .A2(new_n292), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT86), .ZN(new_n682));
  OR3_X1    g0482(.A1(new_n569), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n682), .B1(new_n569), .B2(new_n681), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n680), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n650), .B1(new_n679), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT31), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI211_X1 g0488(.A(KEYINPUT31), .B(new_n650), .C1(new_n679), .C2(new_n685), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n690), .A2(KEYINPUT87), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n609), .A2(new_n504), .A3(new_n580), .A4(new_n651), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n690), .B2(KEYINPUT87), .ZN(new_n693));
  OAI21_X1  g0493(.A(G330), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n650), .B1(new_n625), .B2(new_n640), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n695), .A2(KEYINPUT29), .ZN(new_n696));
  AOI211_X1 g0496(.A(new_n498), .B(new_n579), .C1(new_n659), .C2(new_n607), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT26), .B1(new_n637), .B2(new_n638), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n626), .A2(new_n634), .A3(new_n629), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(new_n699), .A3(new_n570), .ZN(new_n700));
  OAI211_X1 g0500(.A(KEYINPUT29), .B(new_n651), .C1(new_n697), .C2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n694), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n673), .B1(new_n703), .B2(G1), .ZN(G364));
  NAND2_X1  g0504(.A1(new_n222), .A2(G13), .ZN(new_n705));
  XOR2_X1   g0505(.A(new_n705), .B(KEYINPUT88), .Z(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(new_n480), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n707), .A2(new_n258), .A3(new_n668), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n656), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(G330), .B2(new_n655), .ZN(new_n710));
  NOR2_X1   g0510(.A1(G13), .A2(G33), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G20), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n655), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n270), .A2(new_n225), .ZN(new_n716));
  INV_X1    g0516(.A(G355), .ZN(new_n717));
  OAI22_X1  g0517(.A1(new_n716), .A2(new_n717), .B1(G116), .B2(new_n225), .ZN(new_n718));
  MUX2_X1   g0518(.A(new_n221), .B(new_n242), .S(G45), .Z(new_n719));
  NOR2_X1   g0519(.A1(new_n399), .A2(new_n400), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n667), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n718), .B1(new_n719), .B2(new_n722), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n575), .A2(KEYINPUT89), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n575), .A2(KEYINPUT89), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n222), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n223), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n713), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n708), .B1(new_n723), .B2(new_n729), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n730), .A2(KEYINPUT90), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(KEYINPUT90), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n222), .A2(new_n266), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n341), .A2(G179), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(G303), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n222), .A2(G190), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n292), .A2(G200), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G311), .ZN(new_n740));
  OAI22_X1  g0540(.A1(new_n735), .A2(new_n736), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n733), .A2(new_n738), .ZN(new_n742));
  INV_X1    g0542(.A(G322), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n377), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n292), .A2(new_n341), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT94), .ZN(new_n746));
  AND3_X1   g0546(.A1(new_n745), .A2(new_n746), .A3(new_n737), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n746), .B1(new_n745), .B2(new_n737), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  XNOR2_X1  g0550(.A(KEYINPUT33), .B(G317), .ZN(new_n751));
  AOI211_X1 g0551(.A(new_n741), .B(new_n744), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n737), .A2(new_n734), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G179), .A2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n737), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI22_X1  g0557(.A1(G283), .A2(new_n754), .B1(new_n757), .B2(G329), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT96), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n733), .A2(new_n745), .ZN(new_n760));
  INV_X1    g0560(.A(G326), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n222), .B1(new_n755), .B2(G190), .ZN(new_n762));
  INV_X1    g0562(.A(G294), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n760), .A2(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT95), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n752), .A2(new_n759), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n760), .A2(new_n202), .B1(new_n739), .B2(new_n215), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n742), .A2(new_n371), .B1(new_n753), .B2(new_n357), .ZN(new_n770));
  INV_X1    g0570(.A(new_n762), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n769), .B(new_n770), .C1(G97), .C2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n270), .B1(new_n735), .B2(new_n208), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT93), .Z(new_n774));
  OAI211_X1 g0574(.A(new_n772), .B(new_n774), .C1(new_n313), .C2(new_n749), .ZN(new_n775));
  XOR2_X1   g0575(.A(KEYINPUT91), .B(G159), .Z(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n756), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT92), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT32), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n768), .B1(new_n775), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(new_n727), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n731), .A2(new_n732), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n710), .B1(new_n715), .B2(new_n782), .ZN(G396));
  NAND3_X1  g0583(.A1(new_n354), .A2(new_n366), .A3(new_n651), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n354), .A2(new_n650), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n364), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n785), .B1(new_n787), .B2(new_n367), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n695), .B(new_n788), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n694), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n708), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n694), .A2(new_n789), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n776), .ZN(new_n794));
  INV_X1    g0594(.A(new_n739), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(G143), .ZN(new_n797));
  INV_X1    g0597(.A(new_n760), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n750), .A2(G150), .B1(G137), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n799), .A2(KEYINPUT99), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(KEYINPUT99), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n796), .B1(new_n797), .B2(new_n742), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n802), .B(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n735), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G50), .A2(new_n805), .B1(new_n757), .B2(G132), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n806), .B1(new_n371), .B2(new_n762), .C1(new_n313), .C2(new_n753), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n804), .A2(new_n720), .A3(new_n807), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n760), .A2(new_n736), .B1(new_n742), .B2(new_n763), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G87), .A2(new_n754), .B1(new_n795), .B2(G116), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n210), .B2(new_n762), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n809), .B(new_n811), .C1(G311), .C2(new_n757), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n377), .B1(new_n735), .B2(new_n357), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT97), .ZN(new_n814));
  INV_X1    g0614(.A(G283), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n812), .B(new_n814), .C1(new_n815), .C2(new_n749), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT98), .Z(new_n817));
  OAI21_X1  g0617(.A(new_n727), .B1(new_n808), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n727), .A2(new_n711), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n791), .B1(new_n215), .B2(new_n819), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n818), .B(new_n820), .C1(new_n788), .C2(new_n712), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n793), .A2(new_n821), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT101), .Z(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(G384));
  AND2_X1   g0624(.A1(new_n511), .A2(new_n512), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n825), .A2(KEYINPUT35), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(KEYINPUT35), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n223), .A2(new_n222), .A3(new_n591), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT36), .Z(new_n830));
  OR3_X1    g0630(.A1(new_n372), .A2(new_n220), .A3(new_n215), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n202), .A2(G68), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n258), .B(G13), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n338), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n835), .A2(new_n329), .A3(new_n332), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n836), .A2(new_n317), .A3(new_n651), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n431), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n415), .A2(new_n376), .ZN(new_n840));
  INV_X1    g0640(.A(new_n404), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n412), .B1(new_n841), .B2(new_n411), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n370), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n843), .A2(KEYINPUT103), .A3(new_n253), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n416), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n405), .A2(new_n376), .A3(new_n415), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n348), .B1(new_n846), .B2(new_n370), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n847), .A2(KEYINPUT103), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n430), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n839), .B1(new_n849), .B2(new_n442), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT104), .ZN(new_n851));
  INV_X1    g0651(.A(new_n430), .ZN(new_n852));
  INV_X1    g0652(.A(new_n416), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n847), .B2(KEYINPUT103), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n843), .A2(new_n253), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT103), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n852), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n851), .B1(new_n858), .B2(new_n648), .ZN(new_n859));
  INV_X1    g0659(.A(new_n648), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n849), .A2(KEYINPUT104), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n850), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT37), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n434), .A2(new_n442), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n434), .A2(new_n860), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT37), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n864), .A2(new_n865), .A3(new_n866), .A4(new_n431), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n445), .A2(new_n432), .B1(new_n859), .B2(new_n861), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n868), .A2(KEYINPUT38), .A3(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n865), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n446), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n864), .A2(new_n865), .A3(new_n431), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(KEYINPUT37), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n867), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT38), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT39), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n871), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT38), .ZN(new_n881));
  INV_X1    g0681(.A(new_n867), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(new_n862), .B2(KEYINPUT37), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n881), .B1(new_n883), .B2(new_n869), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n871), .A2(new_n884), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n880), .A2(KEYINPUT105), .B1(new_n885), .B2(KEYINPUT39), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT105), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n887), .B(new_n879), .C1(new_n871), .C2(new_n884), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n838), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n885), .ZN(new_n890));
  INV_X1    g0690(.A(new_n344), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n317), .B(new_n650), .C1(new_n836), .C2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n317), .A2(new_n650), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n339), .A2(new_n344), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  AOI211_X1 g0695(.A(KEYINPUT102), .B(new_n785), .C1(new_n695), .C2(new_n788), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT102), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n641), .A2(new_n651), .A3(new_n788), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n897), .B1(new_n898), .B2(new_n784), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n895), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  OAI22_X1  g0700(.A1(new_n890), .A2(new_n900), .B1(new_n445), .B2(new_n860), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n889), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n448), .A2(new_n701), .A3(new_n696), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n620), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n903), .B(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n788), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n892), .B2(new_n894), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n692), .A2(new_n688), .A3(new_n689), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT38), .B1(new_n868), .B2(new_n870), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n883), .A2(new_n881), .A3(new_n869), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT40), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n908), .A2(new_n909), .A3(KEYINPUT40), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n913), .B2(new_n877), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n448), .A2(new_n909), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n919), .A2(new_n920), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n921), .A2(G330), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n906), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n706), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n924), .B1(new_n258), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n906), .A2(new_n923), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n834), .B1(new_n926), .B2(new_n927), .ZN(G367));
  XOR2_X1   g0728(.A(new_n668), .B(KEYINPUT41), .Z(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n637), .A2(new_n651), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n650), .B1(new_n635), .B2(new_n636), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(new_n578), .A3(new_n542), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n665), .A2(new_n935), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT44), .Z(new_n937));
  NOR2_X1   g0737(.A1(new_n665), .A2(new_n935), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT45), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n661), .ZN(new_n941));
  INV_X1    g0741(.A(new_n661), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n937), .A2(new_n942), .A3(new_n939), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n663), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n656), .B(new_n660), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n945), .B1(new_n946), .B2(new_n662), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n703), .A2(KEYINPUT108), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n703), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT108), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n944), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n703), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n930), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n707), .A2(new_n258), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n661), .A2(new_n934), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT107), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n573), .A2(new_n651), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n621), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n638), .A2(new_n959), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n958), .B(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n663), .A2(new_n933), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT106), .Z(new_n968));
  INV_X1    g0768(.A(KEYINPUT42), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n578), .B1(new_n935), .B2(new_n659), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n651), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n968), .A2(new_n969), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n966), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n965), .B(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n956), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n722), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n728), .B1(new_n225), .B2(new_n350), .C1(new_n979), .C2(new_n238), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n980), .A2(new_n708), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n749), .A2(new_n776), .B1(new_n202), .B2(new_n739), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT110), .Z(new_n983));
  INV_X1    g0783(.A(G150), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n270), .B1(new_n762), .B2(new_n313), .C1(new_n984), .C2(new_n742), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n735), .A2(new_n371), .B1(new_n753), .B2(new_n215), .ZN(new_n986));
  INV_X1    g0786(.A(G137), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n760), .A2(new_n797), .B1(new_n756), .B2(new_n987), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n985), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n735), .A2(new_n591), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT46), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n749), .A2(new_n763), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n760), .A2(new_n740), .B1(new_n742), .B2(new_n736), .ZN(new_n993));
  INV_X1    g0793(.A(G317), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n753), .A2(new_n210), .B1(new_n756), .B2(new_n994), .ZN(new_n995));
  NOR4_X1   g0795(.A1(new_n991), .A2(new_n992), .A3(new_n993), .A4(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(G283), .A2(new_n795), .B1(new_n771), .B2(G107), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n997), .A2(KEYINPUT109), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n997), .A2(KEYINPUT109), .ZN(new_n999));
  NOR3_X1   g0799(.A1(new_n998), .A2(new_n999), .A3(new_n721), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n983), .A2(new_n989), .B1(new_n996), .B2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1001), .A2(KEYINPUT47), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(KEYINPUT47), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n727), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n981), .B1(new_n1002), .B2(new_n1004), .C1(new_n963), .C2(new_n714), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n978), .A2(new_n1005), .ZN(G387));
  INV_X1    g0806(.A(new_n955), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n660), .A2(new_n714), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n716), .A2(new_n670), .B1(G107), .B2(new_n225), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n234), .A2(G45), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n249), .A2(G50), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT50), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n670), .B(new_n480), .C1(new_n313), .C2(new_n215), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT111), .Z(new_n1014));
  AOI21_X1  g0814(.A(new_n979), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1009), .B1(new_n1010), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n708), .B1(new_n1016), .B2(new_n729), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n805), .A2(G77), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n984), .B2(new_n756), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n1019), .A2(KEYINPUT112), .B1(G97), .B2(new_n754), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1020), .B(new_n721), .C1(KEYINPUT112), .C2(new_n1019), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT113), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n762), .A2(new_n350), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G159), .A2(new_n798), .B1(new_n795), .B2(G68), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n202), .B2(new_n742), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1023), .B(new_n1025), .C1(new_n352), .C2(new_n750), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1022), .A2(new_n1026), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n735), .A2(new_n763), .B1(new_n762), .B2(new_n815), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G322), .A2(new_n798), .B1(new_n795), .B2(G303), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n994), .B2(new_n742), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(new_n750), .B2(G311), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1028), .B1(new_n1031), .B2(KEYINPUT48), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(KEYINPUT48), .B2(new_n1031), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT49), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n720), .B1(new_n591), .B2(new_n753), .C1(new_n761), .C2(new_n756), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT114), .Z(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1027), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1017), .B1(new_n1039), .B2(new_n727), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n947), .A2(new_n1007), .B1(new_n1008), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n949), .A2(new_n668), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n947), .A2(new_n703), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1041), .B1(new_n1042), .B2(new_n1043), .ZN(G393));
  AOI21_X1  g0844(.A(new_n669), .B1(new_n944), .B2(new_n949), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n951), .A2(new_n948), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1045), .B1(new_n944), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n941), .A2(new_n943), .A3(new_n1007), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n728), .B1(new_n210), .B2(new_n225), .C1(new_n979), .C2(new_n245), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n708), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n771), .A2(G77), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n249), .B2(new_n739), .C1(new_n749), .C2(new_n202), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT115), .Z(new_n1053));
  OAI22_X1  g0853(.A1(new_n760), .A2(new_n984), .B1(new_n742), .B2(new_n374), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT51), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n753), .A2(new_n208), .B1(new_n756), .B2(new_n797), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G68), .B2(new_n805), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1053), .A2(new_n721), .A3(new_n1055), .A4(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT116), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n760), .A2(new_n994), .B1(new_n742), .B2(new_n740), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT52), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n750), .A2(G303), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n735), .A2(new_n815), .B1(new_n739), .B2(new_n763), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(G322), .B2(new_n757), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n377), .B1(new_n753), .B2(new_n357), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(G116), .B2(new_n771), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .A4(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1060), .A2(new_n1061), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1050), .B1(new_n1070), .B2(new_n727), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n934), .B2(new_n714), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1047), .A2(new_n1048), .A3(new_n1072), .ZN(G390));
  AOI21_X1  g0873(.A(new_n791), .B1(new_n249), .B2(new_n819), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT118), .Z(new_n1075));
  OAI22_X1  g0875(.A1(new_n742), .A2(new_n591), .B1(new_n753), .B2(new_n313), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n270), .B(new_n1076), .C1(G87), .C2(new_n805), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n750), .A2(G107), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n739), .A2(new_n210), .B1(new_n756), .B2(new_n763), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(G283), .B2(new_n798), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1077), .A2(new_n1051), .A3(new_n1078), .A4(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(KEYINPUT54), .B(G143), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n798), .A2(G128), .B1(new_n795), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(G132), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1084), .B1(new_n1085), .B2(new_n742), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n735), .A2(new_n984), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT53), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n1088), .A2(new_n1089), .B1(new_n374), .B2(new_n762), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n1089), .B2(new_n1088), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1087), .B(new_n1091), .C1(new_n987), .C2(new_n749), .ZN(new_n1092));
  INV_X1    g0892(.A(G125), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n270), .B1(new_n756), .B2(new_n1093), .C1(new_n202), .C2(new_n753), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT119), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1081), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1075), .B1(new_n727), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(KEYINPUT39), .B1(new_n912), .B2(new_n913), .ZN(new_n1098));
  NOR3_X1   g0898(.A1(new_n913), .A2(KEYINPUT39), .A3(new_n877), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1098), .B1(new_n1099), .B2(new_n887), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n885), .A2(KEYINPUT105), .A3(KEYINPUT39), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1097), .B1(new_n1102), .B2(new_n712), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n900), .A2(new_n837), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n869), .B1(new_n863), .B2(new_n867), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n877), .B1(new_n1105), .B2(KEYINPUT38), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n887), .B1(new_n1106), .B2(new_n879), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n879), .B1(new_n871), .B2(new_n884), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1104), .B(new_n1101), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n697), .A2(new_n700), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1110), .A2(new_n650), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n787), .A2(new_n367), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n785), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n895), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n837), .B1(new_n913), .B2(new_n877), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1109), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n908), .A2(new_n909), .A3(G330), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g0919(.A(G330), .B(new_n908), .C1(new_n691), .C2(new_n693), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1109), .A2(new_n1115), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1103), .B1(new_n1122), .B2(new_n955), .ZN(new_n1123));
  AND3_X1   g0923(.A1(new_n909), .A2(G330), .A3(new_n788), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1120), .B(new_n1113), .C1(new_n895), .C2(new_n1124), .ZN(new_n1125));
  OAI211_X1 g0925(.A(G330), .B(new_n788), .C1(new_n691), .C2(new_n693), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1118), .B1(new_n1126), .B2(new_n1114), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n896), .A2(new_n899), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1125), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n369), .A2(G330), .A3(new_n909), .A4(new_n447), .ZN(new_n1130));
  OR2_X1    g0930(.A1(new_n1130), .A2(KEYINPUT117), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(KEYINPUT117), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1131), .A2(new_n620), .A3(new_n904), .A4(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1129), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1119), .A2(new_n1136), .A3(new_n1121), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n669), .B1(new_n1122), .B2(new_n1135), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1123), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(G378));
  INV_X1    g0940(.A(KEYINPUT57), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n910), .B1(new_n871), .B2(new_n884), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n918), .B(G330), .C1(new_n1142), .C2(KEYINPUT40), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n261), .A2(new_n860), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n298), .B(new_n1144), .ZN(new_n1145));
  XOR2_X1   g0945(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1146));
  XNOR2_X1  g0946(.A(new_n1145), .B(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1143), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1147), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n916), .A2(G330), .A3(new_n918), .A4(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n903), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT122), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n889), .A2(new_n1148), .A3(new_n1150), .A4(new_n902), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n889), .A2(new_n902), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(KEYINPUT122), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n1109), .A2(new_n1115), .A3(new_n1120), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1117), .B1(new_n1109), .B2(new_n1115), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1133), .B1(new_n1161), .B2(new_n1129), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1141), .B1(new_n1158), .B2(new_n1162), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n901), .B1(new_n1102), .B2(new_n838), .ZN(new_n1165));
  OAI21_X1  g0965(.A(KEYINPUT123), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT123), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n903), .A2(new_n1151), .A3(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1166), .A2(new_n1168), .A3(new_n1154), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT124), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1137), .A2(new_n1134), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .A4(KEYINPUT57), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1163), .A2(new_n1172), .A3(new_n668), .ZN(new_n1173));
  AND4_X1   g0973(.A1(new_n889), .A2(new_n902), .A3(new_n1148), .A4(new_n1150), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n1167), .B2(new_n1156), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1141), .B1(new_n1175), .B2(new_n1166), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1170), .B1(new_n1176), .B2(new_n1171), .ZN(new_n1177));
  OR2_X1    g0977(.A1(new_n1173), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1158), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1147), .A2(new_n711), .ZN(new_n1180));
  AOI211_X1 g0980(.A(G33), .B(G41), .C1(new_n794), .C2(new_n754), .ZN(new_n1181));
  INV_X1    g0981(.A(G124), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1181), .B1(new_n1182), .B2(new_n756), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n735), .A2(new_n1082), .B1(new_n739), .B2(new_n987), .ZN(new_n1184));
  INV_X1    g0984(.A(G128), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n760), .A2(new_n1093), .B1(new_n742), .B2(new_n1185), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1184), .B(new_n1186), .C1(G150), .C2(new_n771), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n1085), .B2(new_n749), .ZN(new_n1188));
  XOR2_X1   g0988(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1189));
  AOI21_X1  g0989(.A(new_n1183), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1018), .B1(new_n313), .B2(new_n762), .C1(new_n357), .C2(new_n742), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n739), .A2(new_n350), .B1(new_n756), .B2(new_n815), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n760), .A2(new_n591), .B1(new_n753), .B2(new_n371), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n721), .A2(G41), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1195), .B(new_n1196), .C1(new_n210), .C2(new_n749), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT58), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1196), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1201), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1202));
  AND4_X1   g1002(.A1(new_n1191), .A2(new_n1199), .A3(new_n1200), .A4(new_n1202), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1203), .A2(KEYINPUT121), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(KEYINPUT121), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n1204), .A2(new_n727), .A3(new_n1205), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n791), .B(new_n1206), .C1(new_n202), .C2(new_n819), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1179), .A2(new_n1007), .B1(new_n1180), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1178), .A2(new_n1208), .ZN(G375));
  OAI211_X1 g1009(.A(new_n1133), .B(new_n1125), .C1(new_n1128), .C2(new_n1127), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1135), .A2(new_n930), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1114), .A2(new_n711), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n750), .A2(new_n1083), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n371), .A2(new_n753), .B1(new_n739), .B2(new_n984), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(G50), .B2(new_n771), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n760), .A2(new_n1085), .B1(new_n742), .B2(new_n987), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n735), .A2(new_n374), .B1(new_n756), .B2(new_n1185), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1213), .A2(new_n721), .A3(new_n1215), .A4(new_n1218), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n760), .A2(new_n763), .B1(new_n735), .B2(new_n210), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n742), .A2(new_n815), .B1(new_n756), .B2(new_n736), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n739), .A2(new_n357), .ZN(new_n1222));
  NOR4_X1   g1022(.A1(new_n1220), .A2(new_n1221), .A3(new_n1023), .A4(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n591), .B2(new_n749), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n377), .B1(new_n753), .B2(new_n215), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1225), .B(KEYINPUT125), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1219), .B1(new_n1224), .B2(new_n1226), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n1227), .A2(new_n727), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n791), .B(new_n1228), .C1(new_n313), .C2(new_n819), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1129), .A2(new_n1007), .B1(new_n1212), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1211), .A2(new_n1230), .ZN(G381));
  NAND3_X1  g1031(.A1(new_n1178), .A2(new_n1139), .A3(new_n1208), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n976), .B1(new_n954), .B2(new_n955), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1005), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1234), .A2(new_n1235), .A3(G390), .ZN(new_n1236));
  NOR4_X1   g1036(.A1(G384), .A2(G396), .A3(G393), .A4(G381), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1233), .A2(new_n1236), .A3(new_n1237), .ZN(G407));
  OAI211_X1 g1038(.A(G407), .B(G213), .C1(G343), .C2(new_n1232), .ZN(G409));
  NAND2_X1  g1039(.A1(new_n649), .A2(G213), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(G378), .B(new_n1208), .C1(new_n1173), .C2(new_n1177), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1158), .A2(new_n1162), .A3(new_n929), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1169), .A2(new_n1007), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1180), .A2(new_n1207), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1139), .B1(new_n1243), .B2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1241), .B1(new_n1242), .B2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n669), .B1(new_n1129), .B2(new_n1134), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1210), .A2(KEYINPUT60), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1210), .A2(KEYINPUT60), .ZN(new_n1251));
  OAI211_X1 g1051(.A(KEYINPUT126), .B(new_n1249), .C1(new_n1250), .C2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1230), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1210), .B(KEYINPUT60), .ZN(new_n1254));
  AOI21_X1  g1054(.A(KEYINPUT126), .B1(new_n1254), .B2(new_n1249), .ZN(new_n1255));
  OAI21_X1  g1055(.A(G384), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1249), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT126), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1259), .A2(new_n823), .A3(new_n1230), .A4(new_n1252), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1256), .A2(new_n1260), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1240), .A2(KEYINPUT127), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n1261), .A2(new_n1263), .B1(G2897), .B2(new_n1241), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1241), .A2(G2897), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n1265), .B(new_n1262), .C1(new_n1256), .C2(new_n1260), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(KEYINPUT63), .B1(new_n1248), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1248), .A2(new_n1261), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1248), .A2(KEYINPUT63), .A3(new_n1261), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(G387), .A2(G390), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1236), .ZN(new_n1273));
  XOR2_X1   g1073(.A(G393), .B(G396), .Z(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1272), .A2(new_n1273), .A3(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(G390), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(new_n978), .B2(new_n1005), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1274), .B1(new_n1278), .B2(new_n1236), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1276), .A2(new_n1279), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1280), .A2(KEYINPUT61), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1270), .A2(new_n1271), .A3(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT62), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1248), .A2(new_n1283), .A3(new_n1261), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT61), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1285), .B1(new_n1248), .B2(new_n1267), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1283), .B1(new_n1248), .B2(new_n1261), .ZN(new_n1287));
  NOR3_X1   g1087(.A1(new_n1284), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1280), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1282), .B1(new_n1288), .B2(new_n1289), .ZN(G405));
  INV_X1    g1090(.A(new_n1261), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1139), .B1(new_n1178), .B2(new_n1208), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1291), .B1(new_n1233), .B2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1292), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1294), .A2(new_n1232), .A3(new_n1261), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1280), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1293), .A2(new_n1295), .A3(new_n1289), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(G402));
endmodule


