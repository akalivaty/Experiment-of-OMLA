//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1285,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G250), .ZN(new_n206));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G257), .ZN(new_n213));
  INV_X1    g0013(.A(G264), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n206), .B(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n215), .A2(KEYINPUT0), .ZN(new_n216));
  AND2_X1   g0016(.A1(KEYINPUT64), .A2(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(KEYINPUT64), .A2(G20), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n202), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(G50), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(new_n215), .A2(KEYINPUT0), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n227));
  INV_X1    g0027(.A(G77), .ZN(new_n228));
  INV_X1    g0028(.A(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G107), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n227), .B1(new_n228), .B2(new_n229), .C1(new_n230), .C2(new_n214), .ZN(new_n231));
  AOI22_X1  g0031(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  INV_X1    g0033(.A(G97), .ZN(new_n234));
  OAI221_X1 g0034(.A(new_n232), .B1(new_n202), .B2(new_n233), .C1(new_n234), .C2(new_n213), .ZN(new_n235));
  OAI21_X1  g0035(.A(new_n210), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  OR2_X1    g0036(.A1(new_n236), .A2(KEYINPUT1), .ZN(new_n237));
  NAND3_X1  g0037(.A1(new_n216), .A2(new_n226), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g0038(.A(new_n238), .B1(KEYINPUT1), .B2(new_n236), .ZN(G361));
  XOR2_X1   g0039(.A(G238), .B(G244), .Z(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT65), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n244), .B(KEYINPUT66), .Z(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G264), .B(G270), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G358));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT67), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(G68), .B(G77), .Z(new_n254));
  XOR2_X1   g0054(.A(G50), .B(G58), .Z(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n253), .B(new_n256), .ZN(G351));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  AOI21_X1  g0061(.A(G1698), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G222), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n260), .A2(new_n261), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(G223), .A3(G1698), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n263), .B(new_n265), .C1(new_n228), .C2(new_n264), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n220), .B1(G33), .B2(G41), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G41), .ZN(new_n269));
  OAI211_X1 g0069(.A(G1), .B(G13), .C1(new_n259), .C2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT68), .B(G45), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n269), .ZN(new_n274));
  INV_X1    g0074(.A(G274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n275), .A2(G1), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n272), .A2(G226), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n268), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G179), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G150), .ZN(new_n283));
  OAI21_X1  g0083(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n219), .A2(G33), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n283), .B(new_n284), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n220), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(new_n289), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n201), .B1(new_n207), .B2(G20), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n293), .A2(new_n294), .B1(new_n201), .B2(new_n292), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n290), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n281), .B(new_n296), .C1(G169), .C2(new_n279), .ZN(new_n297));
  INV_X1    g0097(.A(new_n289), .ZN(new_n298));
  INV_X1    g0098(.A(new_n286), .ZN(new_n299));
  OR2_X1    g0099(.A1(KEYINPUT64), .A2(G20), .ZN(new_n300));
  NAND2_X1  g0100(.A1(KEYINPUT64), .A2(G20), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n299), .A2(new_n282), .B1(new_n302), .B2(G77), .ZN(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT15), .B(G87), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n305), .A2(G33), .A3(new_n219), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n298), .B1(new_n303), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n207), .A2(G20), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n293), .A2(G77), .A3(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(G77), .B2(new_n291), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n274), .A2(new_n276), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n270), .A2(new_n271), .ZN(new_n314));
  NOR2_X1   g0114(.A1(G232), .A2(G1698), .ZN(new_n315));
  INV_X1    g0115(.A(G238), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n315), .B1(new_n316), .B2(G1698), .ZN(new_n317));
  AND2_X1   g0117(.A1(KEYINPUT3), .A2(G33), .ZN(new_n318));
  NOR2_X1   g0118(.A1(KEYINPUT3), .A2(G33), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n267), .B1(new_n264), .B2(G107), .ZN(new_n322));
  OAI221_X1 g0122(.A(new_n313), .B1(new_n229), .B2(new_n314), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n323), .A2(G179), .ZN(new_n324));
  INV_X1    g0124(.A(G169), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n312), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n323), .A2(G200), .ZN(new_n328));
  INV_X1    g0128(.A(G190), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n311), .B(new_n328), .C1(new_n329), .C2(new_n323), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  OR2_X1    g0131(.A1(new_n296), .A2(KEYINPUT9), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n296), .A2(KEYINPUT9), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n332), .A2(new_n333), .B1(G200), .B2(new_n278), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT10), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT69), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n336), .B1(new_n279), .B2(G190), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n334), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n335), .B1(new_n334), .B2(new_n337), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n297), .B(new_n331), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT70), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n340), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n338), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n345), .A2(KEYINPUT70), .A3(new_n297), .A4(new_n331), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n282), .A2(G50), .B1(G20), .B2(new_n222), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(new_n285), .B2(new_n228), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n348), .A2(KEYINPUT11), .A3(new_n289), .ZN(new_n349));
  AOI21_X1  g0149(.A(KEYINPUT11), .B1(new_n348), .B2(new_n289), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n293), .A2(G68), .A3(new_n308), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT12), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(new_n292), .B2(new_n222), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n291), .A2(KEYINPUT12), .A3(G68), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n351), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OR3_X1    g0155(.A1(new_n349), .A2(new_n350), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n233), .A2(G1698), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n264), .B(new_n357), .C1(G226), .C2(G1698), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G33), .A2(G97), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n270), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT13), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n272), .A2(G238), .B1(new_n274), .B2(new_n276), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n313), .B1(new_n316), .B2(new_n314), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT13), .B1(new_n365), .B2(new_n360), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT72), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT14), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(G169), .A3(new_n369), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n361), .A2(new_n363), .B1(KEYINPUT71), .B2(KEYINPUT13), .ZN(new_n371));
  NAND2_X1  g0171(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n372));
  NOR3_X1   g0172(.A1(new_n365), .A2(new_n360), .A3(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n370), .B1(new_n280), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n369), .B1(new_n367), .B2(G169), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n356), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n356), .B1(G200), .B2(new_n367), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n329), .B2(new_n374), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n343), .A2(new_n346), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n293), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n299), .A2(new_n308), .ZN(new_n383));
  OAI22_X1  g0183(.A1(new_n382), .A2(new_n383), .B1(new_n291), .B2(new_n299), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(G223), .ZN(new_n386));
  INV_X1    g0186(.A(G1698), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n264), .B(new_n388), .C1(G226), .C2(new_n387), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G87), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n267), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n272), .A2(G232), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n392), .A2(G190), .A3(new_n393), .A4(new_n313), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n313), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n270), .B1(new_n389), .B2(new_n390), .ZN(new_n396));
  OAI21_X1  g0196(.A(G200), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT76), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n300), .A2(new_n260), .A3(new_n301), .A4(new_n261), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT7), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n219), .A2(new_n320), .A3(KEYINPUT76), .A4(KEYINPUT7), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT75), .ZN(new_n405));
  NOR3_X1   g0205(.A1(new_n318), .A2(new_n319), .A3(G20), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n405), .B1(new_n406), .B2(KEYINPUT7), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n260), .A2(new_n208), .A3(new_n261), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n408), .A2(KEYINPUT75), .A3(new_n401), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n404), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G68), .ZN(new_n412));
  INV_X1    g0212(.A(G159), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n413), .A2(G20), .A3(G33), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(G58), .A2(G68), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n208), .B1(new_n223), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n415), .B1(new_n417), .B2(KEYINPUT73), .ZN(new_n418));
  AND2_X1   g0218(.A1(G58), .A2(G68), .ZN(new_n419));
  NOR2_X1   g0219(.A1(G58), .A2(G68), .ZN(new_n420));
  OAI211_X1 g0220(.A(KEYINPUT73), .B(G20), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT16), .B1(new_n412), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n219), .A2(new_n320), .A3(new_n401), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n408), .A2(KEYINPUT7), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(new_n426), .A3(G68), .ZN(new_n427));
  OAI21_X1  g0227(.A(G20), .B1(new_n419), .B2(new_n420), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT73), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AND4_X1   g0230(.A1(KEYINPUT74), .A2(new_n430), .A3(new_n421), .A4(new_n415), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n414), .B1(new_n428), .B2(new_n429), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT74), .B1(new_n432), .B2(new_n421), .ZN(new_n433));
  OAI211_X1 g0233(.A(KEYINPUT16), .B(new_n427), .C1(new_n431), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n289), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n385), .B(new_n398), .C1(new_n424), .C2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT17), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(KEYINPUT77), .A3(new_n437), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n425), .A2(new_n426), .A3(G68), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT74), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n418), .B2(new_n422), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n432), .A2(KEYINPUT74), .A3(new_n421), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n298), .B1(new_n443), .B2(KEYINPUT16), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT16), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n222), .B1(new_n404), .B2(new_n410), .ZN(new_n446));
  INV_X1    g0246(.A(new_n423), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n384), .B1(new_n444), .B2(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n392), .A2(G179), .A3(new_n393), .A4(new_n313), .ZN(new_n450));
  OAI21_X1  g0250(.A(G169), .B1(new_n395), .B2(new_n396), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT18), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n385), .B1(new_n424), .B2(new_n435), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT18), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(new_n456), .A3(new_n452), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n437), .A2(KEYINPUT77), .ZN(new_n458));
  OR2_X1    g0258(.A1(new_n437), .A2(KEYINPUT77), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n449), .A2(new_n458), .A3(new_n459), .A4(new_n398), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n438), .A2(new_n454), .A3(new_n457), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n259), .A2(G97), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n219), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G116), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n288), .A2(new_n220), .B1(G20), .B2(new_n465), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n464), .A2(new_n466), .B1(KEYINPUT84), .B2(KEYINPUT20), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT84), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT20), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n291), .A2(new_n465), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n207), .A2(G33), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n291), .A2(new_n473), .A3(new_n220), .A4(new_n288), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n472), .B1(new_n475), .B2(new_n465), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n464), .A2(new_n468), .A3(new_n466), .A4(new_n469), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n471), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G45), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(G1), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT5), .B(G41), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n267), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n481), .A2(new_n480), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n267), .A2(new_n275), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n482), .A2(G270), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(G264), .B(G1698), .C1(new_n318), .C2(new_n319), .ZN(new_n486));
  OAI211_X1 g0286(.A(G257), .B(new_n387), .C1(new_n318), .C2(new_n319), .ZN(new_n487));
  INV_X1    g0287(.A(G303), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n486), .B(new_n487), .C1(new_n488), .C2(new_n264), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n267), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n325), .B1(new_n485), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n478), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT21), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n478), .A2(new_n491), .A3(KEYINPUT21), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n485), .A2(G179), .A3(new_n490), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n478), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n485), .A2(new_n490), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n478), .B1(G200), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(new_n329), .B2(new_n499), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n300), .B(new_n301), .C1(new_n318), .C2(new_n319), .ZN(new_n503));
  INV_X1    g0303(.A(G87), .ZN(new_n504));
  OAI21_X1  g0304(.A(KEYINPUT22), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT22), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n264), .A2(new_n219), .A3(new_n506), .A4(G87), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(KEYINPUT23), .B1(new_n208), .B2(G107), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G116), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n509), .B1(G20), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(KEYINPUT23), .A2(G107), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n511), .B1(new_n302), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g0314(.A(KEYINPUT85), .B(KEYINPUT24), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n515), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n508), .A2(new_n513), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n298), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(G13), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n520), .A2(G1), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n521), .A2(G20), .A3(new_n230), .ZN(new_n522));
  XNOR2_X1  g0322(.A(new_n522), .B(KEYINPUT25), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n474), .A2(new_n230), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(KEYINPUT86), .B1(new_n519), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n518), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n517), .B1(new_n508), .B2(new_n513), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n289), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT86), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(new_n531), .A3(new_n525), .ZN(new_n532));
  OAI211_X1 g0332(.A(G257), .B(G1698), .C1(new_n318), .C2(new_n319), .ZN(new_n533));
  OAI211_X1 g0333(.A(G250), .B(new_n387), .C1(new_n318), .C2(new_n319), .ZN(new_n534));
  INV_X1    g0334(.A(G294), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n533), .B(new_n534), .C1(new_n259), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n267), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n481), .A2(new_n480), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n538), .A2(G264), .A3(new_n270), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n483), .A2(new_n484), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n537), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G169), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n539), .A2(KEYINPUT87), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT87), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n482), .A2(new_n544), .A3(G264), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n537), .A2(new_n543), .A3(new_n545), .A4(new_n540), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n542), .B1(new_n280), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n527), .A2(new_n532), .A3(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n519), .A2(new_n526), .ZN(new_n549));
  INV_X1    g0349(.A(G200), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(G190), .B2(new_n541), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n502), .A2(new_n548), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT80), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT78), .ZN(new_n556));
  INV_X1    g0356(.A(new_n282), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n556), .B1(new_n557), .B2(new_n228), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n282), .A2(KEYINPUT78), .A3(G77), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g0360(.A(G97), .B(G107), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT6), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NOR3_X1   g0363(.A1(new_n562), .A2(new_n234), .A3(G107), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n560), .B1(new_n565), .B2(new_n219), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n411), .A2(G107), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n566), .B1(new_n567), .B2(KEYINPUT79), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT79), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n411), .A2(new_n569), .A3(G107), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n298), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n291), .A2(G97), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n475), .B2(G97), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n555), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n402), .A2(new_n403), .B1(new_n407), .B2(new_n409), .ZN(new_n576));
  OAI21_X1  g0376(.A(KEYINPUT79), .B1(new_n576), .B2(new_n230), .ZN(new_n577));
  INV_X1    g0377(.A(new_n566), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n577), .A2(new_n570), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n289), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(KEYINPUT80), .A3(new_n573), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n264), .A2(G250), .A3(G1698), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n462), .ZN(new_n583));
  XOR2_X1   g0383(.A(KEYINPUT81), .B(KEYINPUT4), .Z(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(G244), .B2(new_n262), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n264), .A2(KEYINPUT4), .A3(G244), .A4(new_n387), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT82), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n262), .A2(KEYINPUT82), .A3(KEYINPUT4), .A4(G244), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n267), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n482), .A2(G257), .B1(new_n483), .B2(new_n484), .ZN(new_n594));
  OR2_X1    g0394(.A1(new_n594), .A2(KEYINPUT83), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(KEYINPUT83), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n593), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n270), .B1(new_n586), .B2(new_n591), .ZN(new_n598));
  INV_X1    g0398(.A(new_n594), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n597), .A2(G200), .B1(new_n600), .B2(G190), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n575), .A2(new_n581), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n580), .A2(new_n573), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n593), .A2(new_n280), .A3(new_n595), .A4(new_n596), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n325), .B1(new_n598), .B2(new_n599), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n504), .A2(new_n234), .A3(new_n230), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT19), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n359), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n608), .B1(new_n302), .B2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n300), .A2(G33), .A3(G97), .A4(new_n301), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n609), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n611), .B(new_n613), .C1(new_n222), .C2(new_n503), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n289), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n480), .A2(new_n275), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n206), .B1(new_n479), .B2(G1), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(new_n270), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n316), .A2(new_n387), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n229), .A2(G1698), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n619), .B(new_n620), .C1(new_n318), .C2(new_n319), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n621), .A2(new_n510), .ZN(new_n622));
  OAI211_X1 g0422(.A(G190), .B(new_n618), .C1(new_n622), .C2(new_n270), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n305), .A2(new_n291), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n474), .A2(new_n504), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n615), .A2(new_n623), .A3(new_n625), .A4(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n270), .B1(new_n621), .B2(new_n510), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n616), .A2(new_n270), .A3(new_n617), .ZN(new_n631));
  OAI21_X1  g0431(.A(G200), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n615), .B(new_n625), .C1(new_n304), .C2(new_n474), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n280), .B(new_n618), .C1(new_n622), .C2(new_n270), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n325), .B1(new_n630), .B2(new_n631), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n629), .A2(new_n632), .B1(new_n633), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n602), .A2(new_n607), .A3(new_n638), .ZN(new_n639));
  NOR4_X1   g0439(.A1(new_n381), .A2(new_n461), .A3(new_n554), .A4(new_n639), .ZN(G372));
  NOR2_X1   g0440(.A1(new_n381), .A2(new_n461), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT88), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n632), .A2(new_n642), .ZN(new_n643));
  OAI211_X1 g0443(.A(KEYINPUT88), .B(G200), .C1(new_n630), .C2(new_n631), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n474), .A2(new_n304), .ZN(new_n646));
  AOI211_X1 g0446(.A(new_n624), .B(new_n646), .C1(new_n614), .C2(new_n289), .ZN(new_n647));
  OAI22_X1  g0447(.A1(new_n628), .A2(new_n645), .B1(new_n647), .B2(new_n636), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT89), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI221_X1 g0450(.A(KEYINPUT89), .B1(new_n647), .B2(new_n636), .C1(new_n645), .C2(new_n628), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n650), .A2(new_n651), .B1(new_n549), .B2(new_n552), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n547), .B1(new_n519), .B2(new_n526), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n498), .A2(new_n653), .ZN(new_n654));
  AND4_X1   g0454(.A1(new_n602), .A2(new_n607), .A3(new_n652), .A4(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n604), .A2(new_n605), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n650), .B2(new_n651), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  AOI21_X1  g0458(.A(KEYINPUT80), .B1(new_n580), .B2(new_n573), .ZN(new_n659));
  AOI211_X1 g0459(.A(new_n555), .B(new_n574), .C1(new_n579), .C2(new_n289), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n657), .B(new_n658), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n633), .A2(new_n637), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n603), .A2(new_n606), .A3(new_n638), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n663), .B1(new_n664), .B2(KEYINPUT26), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n641), .B1(new_n655), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n297), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n438), .A2(new_n460), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n327), .A2(KEYINPUT90), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n327), .A2(KEYINPUT90), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n377), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n669), .A2(new_n673), .A3(new_n379), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n454), .A2(new_n457), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n668), .B1(new_n676), .B2(new_n345), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n667), .A2(new_n677), .ZN(G369));
  NAND2_X1  g0478(.A1(new_n219), .A2(new_n521), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G213), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(G343), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n478), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n502), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n498), .A2(new_n685), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT91), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G330), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n548), .A2(new_n553), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n527), .A2(new_n532), .A3(new_n684), .ZN(new_n692));
  INV_X1    g0492(.A(new_n684), .ZN(new_n693));
  OAI22_X1  g0493(.A1(new_n691), .A2(new_n692), .B1(new_n548), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT92), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n690), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n653), .A2(new_n684), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n694), .B(KEYINPUT92), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n498), .A2(new_n684), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n698), .A2(new_n702), .ZN(G399));
  NOR2_X1   g0503(.A1(new_n212), .A2(G41), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n608), .A2(G116), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(G1), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n224), .B2(new_n705), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT28), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n548), .A2(new_n498), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n602), .A2(new_n607), .A3(new_n652), .A4(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n659), .A2(new_n660), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n650), .A2(new_n651), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n606), .ZN(new_n714));
  OAI21_X1  g0514(.A(KEYINPUT26), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n603), .A2(new_n638), .A3(new_n606), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n663), .B1(new_n716), .B2(new_n658), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n711), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(KEYINPUT29), .A3(new_n693), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n655), .A2(new_n666), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n684), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n719), .B1(new_n721), .B2(KEYINPUT29), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT31), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n630), .A2(new_n631), .ZN(new_n724));
  AND4_X1   g0524(.A1(new_n537), .A2(new_n724), .A3(new_n543), .A4(new_n545), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n593), .A2(new_n725), .A3(new_n496), .A4(new_n594), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n724), .A2(G179), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n546), .A2(new_n499), .A3(new_n728), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n726), .A2(new_n727), .B1(new_n597), .B2(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n600), .A2(KEYINPUT30), .A3(new_n496), .A4(new_n725), .ZN(new_n731));
  AOI211_X1 g0531(.A(new_n723), .B(new_n693), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n726), .A2(new_n727), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n597), .A2(new_n729), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(new_n734), .A3(new_n731), .ZN(new_n735));
  AOI21_X1  g0535(.A(KEYINPUT31), .B1(new_n735), .B2(new_n684), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n502), .A2(new_n548), .A3(new_n553), .A4(new_n693), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n737), .B1(new_n639), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G330), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT93), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n739), .A2(KEYINPUT93), .A3(G330), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n722), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n709), .B1(new_n746), .B2(G1), .ZN(G364));
  INV_X1    g0547(.A(new_n690), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n302), .A2(new_n520), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G45), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G1), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n704), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(G330), .B2(new_n689), .ZN(new_n754));
  INV_X1    g0554(.A(new_n752), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n220), .B1(G20), .B2(new_n325), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n329), .A2(G200), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n219), .A2(new_n280), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT96), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n759), .A2(new_n760), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n758), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT97), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G58), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G179), .A2(G190), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n302), .A2(G200), .A3(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n230), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR4_X1   g0571(.A1(new_n208), .A2(new_n329), .A3(new_n550), .A4(G179), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n771), .B(new_n264), .C1(new_n504), .C2(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n302), .A2(new_n550), .A3(new_n768), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G159), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT32), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n329), .B(new_n550), .C1(new_n762), .C2(new_n763), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n774), .B(new_n778), .C1(G77), .C2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n759), .A2(G200), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G190), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n219), .B1(new_n280), .B2(new_n758), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n784), .A2(new_n222), .B1(new_n234), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT99), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT98), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(new_n782), .B2(new_n329), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n759), .A2(KEYINPUT98), .A3(G190), .A4(G200), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n786), .A2(new_n787), .B1(new_n792), .B2(G50), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n767), .A2(new_n781), .A3(new_n788), .A4(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n264), .B1(new_n772), .B2(G303), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT100), .ZN(new_n796));
  INV_X1    g0596(.A(new_n785), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n797), .A2(G294), .B1(new_n776), .B2(G329), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n799), .B2(new_n769), .ZN(new_n800));
  XNOR2_X1  g0600(.A(KEYINPUT33), .B(G317), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n796), .B(new_n800), .C1(new_n783), .C2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n764), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n780), .A2(G311), .B1(new_n803), .B2(G322), .ZN(new_n804));
  INV_X1    g0604(.A(G326), .ZN(new_n805));
  INV_X1    g0605(.A(new_n792), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n802), .B(new_n804), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n757), .B1(new_n794), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n520), .A2(new_n259), .A3(KEYINPUT95), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT95), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(G13), .B2(G33), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(G20), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n756), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n256), .A2(G45), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n212), .A2(new_n264), .ZN(new_n817));
  INV_X1    g0617(.A(new_n273), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n816), .B(new_n817), .C1(new_n224), .C2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n211), .A2(new_n264), .ZN(new_n820));
  INV_X1    g0620(.A(G355), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n820), .A2(new_n821), .B1(G116), .B2(new_n211), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT94), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n819), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n755), .B(new_n808), .C1(new_n815), .C2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n814), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n827), .B1(new_n688), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n754), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(G396));
  NAND4_X1  g0631(.A1(new_n670), .A2(new_n312), .A3(new_n671), .A4(new_n684), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n331), .B1(new_n311), .B2(new_n693), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n721), .B(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n752), .B1(new_n835), .B2(new_n744), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n744), .B2(new_n835), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n812), .A2(new_n756), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n755), .B1(new_n228), .B2(new_n838), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n779), .A2(new_n465), .B1(new_n764), .B2(new_n535), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n320), .B1(new_n773), .B2(new_n230), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(G97), .B2(new_n797), .ZN(new_n842));
  INV_X1    g0642(.A(new_n769), .ZN(new_n843));
  AOI22_X1  g0643(.A1(G87), .A2(new_n843), .B1(new_n776), .B2(G311), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n842), .B(new_n844), .C1(new_n799), .C2(new_n784), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n840), .B(new_n845), .C1(G303), .C2(new_n792), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n780), .A2(G159), .B1(G150), .B2(new_n783), .ZN(new_n847));
  INV_X1    g0647(.A(G137), .ZN(new_n848));
  INV_X1    g0648(.A(G143), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n847), .B1(new_n848), .B2(new_n806), .C1(new_n765), .C2(new_n849), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT34), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n264), .B1(new_n773), .B2(new_n201), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n785), .A2(new_n202), .B1(new_n769), .B2(new_n222), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n852), .B(new_n853), .C1(G132), .C2(new_n776), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n846), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n839), .B1(new_n813), .B2(new_n834), .C1(new_n855), .C2(new_n757), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n837), .A2(new_n856), .ZN(G384));
  NOR2_X1   g0657(.A1(new_n749), .A2(new_n207), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n427), .B1(new_n431), .B2(new_n433), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n445), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n384), .B1(new_n444), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT101), .B1(new_n861), .B2(new_n682), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n441), .A2(new_n442), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT16), .B1(new_n863), .B2(new_n427), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n385), .B1(new_n435), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT101), .ZN(new_n866));
  INV_X1    g0666(.A(new_n682), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n862), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n461), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT37), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n865), .A2(new_n452), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT102), .B1(new_n872), .B2(new_n436), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n872), .A2(KEYINPUT102), .A3(new_n436), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n871), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n455), .A2(new_n452), .ZN(new_n877));
  XOR2_X1   g0677(.A(new_n682), .B(KEYINPUT103), .Z(new_n878));
  NAND2_X1  g0678(.A1(new_n455), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n877), .A2(new_n879), .A3(new_n871), .A4(new_n436), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(KEYINPUT38), .B(new_n870), .C1(new_n876), .C2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n878), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n449), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n436), .B1(new_n449), .B2(new_n453), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT37), .B1(new_n885), .B2(new_n884), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n461), .A2(new_n884), .B1(new_n886), .B2(new_n880), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT104), .B1(new_n887), .B2(KEYINPUT38), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n461), .A2(new_n884), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n886), .A2(new_n880), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT104), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT38), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n882), .A2(new_n888), .A3(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT39), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n377), .A2(new_n684), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n862), .A2(new_n868), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n872), .A2(new_n436), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT102), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n899), .A2(new_n875), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n881), .B1(new_n903), .B2(KEYINPUT37), .ZN(new_n904));
  INV_X1    g0704(.A(new_n870), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n893), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n906), .A2(KEYINPUT39), .A3(new_n882), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n897), .A2(new_n898), .A3(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n675), .A2(new_n878), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n356), .A2(new_n684), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n380), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n377), .A2(new_n379), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n912), .A2(new_n356), .A3(new_n684), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n693), .B(new_n834), .C1(new_n655), .C2(new_n666), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n327), .A2(new_n684), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n915), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n906), .A2(new_n882), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n909), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n908), .A2(new_n921), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n641), .B(new_n719), .C1(new_n721), .C2(KEYINPUT29), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n677), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n922), .B(new_n924), .Z(new_n925));
  INV_X1    g0725(.A(G330), .ZN(new_n926));
  INV_X1    g0726(.A(new_n834), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n911), .B2(new_n913), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n739), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n920), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT40), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n928), .A2(KEYINPUT40), .A3(new_n739), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n895), .A2(new_n934), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n641), .A2(new_n739), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n926), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n937), .B2(new_n936), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n858), .B1(new_n925), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n925), .B2(new_n939), .ZN(new_n941));
  INV_X1    g0741(.A(new_n565), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n942), .A2(KEYINPUT35), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(KEYINPUT35), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n943), .A2(G116), .A3(new_n221), .A4(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT36), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n225), .A2(G77), .A3(new_n416), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(G50), .B2(new_n222), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n948), .A2(G1), .A3(new_n520), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n941), .A2(new_n946), .A3(new_n949), .ZN(G367));
  AOI21_X1  g0750(.A(new_n624), .B1(new_n614), .B2(new_n289), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n693), .B1(new_n951), .B2(new_n627), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n650), .B2(new_n651), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n663), .B2(new_n952), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n814), .ZN(new_n955));
  INV_X1    g0755(.A(new_n815), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(new_n212), .B2(new_n305), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n817), .A2(new_n248), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n755), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(G150), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n779), .A2(new_n201), .B1(new_n764), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n264), .B1(new_n773), .B2(new_n202), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(G137), .B2(new_n776), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n797), .A2(G68), .B1(new_n843), .B2(G77), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n963), .B(new_n964), .C1(new_n413), .C2(new_n784), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n961), .B(new_n965), .C1(G143), .C2(new_n792), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT113), .Z(new_n967));
  INV_X1    g0767(.A(KEYINPUT46), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n773), .B2(new_n465), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n772), .A2(KEYINPUT46), .A3(G116), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n969), .B(new_n970), .C1(new_n784), .C2(new_n535), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(KEYINPUT111), .Z(new_n972));
  NAND2_X1  g0772(.A1(new_n766), .A2(G303), .ZN(new_n973));
  INV_X1    g0773(.A(G317), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n320), .B1(new_n769), .B2(new_n234), .C1(new_n974), .C2(new_n775), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT112), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n779), .A2(new_n799), .B1(new_n230), .B2(new_n785), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(G311), .B2(new_n792), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n972), .A2(new_n973), .A3(new_n976), .A4(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n967), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT47), .Z(new_n981));
  OAI211_X1 g0781(.A(new_n955), .B(new_n959), .C1(new_n981), .C2(new_n757), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n751), .B(KEYINPUT110), .Z(new_n983));
  INV_X1    g0783(.A(KEYINPUT106), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n684), .B1(new_n659), .B2(new_n660), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n985), .A2(new_n602), .A3(new_n607), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT105), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n985), .A2(new_n602), .A3(KEYINPUT105), .A4(new_n607), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n606), .B(new_n684), .C1(new_n659), .C2(new_n660), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n984), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n991), .ZN(new_n993));
  AOI211_X1 g0793(.A(KEYINPUT106), .B(new_n993), .C1(new_n988), .C2(new_n989), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n701), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n696), .A2(new_n996), .B1(new_n653), .B2(new_n684), .ZN(new_n997));
  AOI21_X1  g0797(.A(KEYINPUT44), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n990), .A2(new_n991), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(KEYINPUT106), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n990), .A2(new_n984), .A3(new_n991), .ZN(new_n1001));
  AND4_X1   g0801(.A1(KEYINPUT44), .A2(new_n1000), .A3(new_n997), .A4(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n995), .B2(new_n997), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1007), .A2(new_n702), .A3(new_n1004), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g0809(.A(KEYINPUT109), .B(new_n697), .C1(new_n1003), .C2(new_n1009), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT44), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n1007), .B2(new_n702), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n995), .A2(KEYINPUT44), .A3(new_n997), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1011), .A2(new_n698), .A3(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n696), .B(new_n701), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(new_n748), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1018), .A2(new_n745), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1010), .A2(new_n1016), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1011), .A2(new_n1015), .ZN(new_n1021));
  AOI21_X1  g0821(.A(KEYINPUT109), .B1(new_n1021), .B2(new_n697), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n746), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n704), .B(KEYINPUT41), .Z(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n983), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1000), .A2(KEYINPUT107), .A3(new_n1001), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT107), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n992), .B2(new_n994), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n697), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT43), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n954), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n954), .A2(new_n1032), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n548), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n607), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n693), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT42), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n696), .A2(new_n996), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1007), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1039), .B1(new_n1007), .B2(new_n1040), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1034), .B(new_n1035), .C1(new_n1038), .C2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1038), .A2(new_n1044), .A3(new_n1032), .A4(new_n954), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1031), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1035), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n1033), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1031), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1050), .A2(new_n1051), .A3(new_n1046), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1048), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n982), .B1(new_n1026), .B2(new_n1053), .ZN(G387));
  INV_X1    g0854(.A(new_n983), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1018), .A2(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT114), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n820), .A2(new_n706), .B1(G107), .B2(new_n211), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT115), .Z(new_n1059));
  NAND2_X1  g0859(.A1(new_n244), .A2(new_n818), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n706), .ZN(new_n1061));
  AOI211_X1 g0861(.A(G45), .B(new_n1061), .C1(G68), .C2(G77), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n286), .A2(G50), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT50), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n212), .B(new_n264), .C1(new_n1062), .C2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1059), .B1(new_n1060), .B2(new_n1065), .ZN(new_n1066));
  XOR2_X1   g0866(.A(KEYINPUT116), .B(G150), .Z(new_n1067));
  OAI22_X1  g0867(.A1(new_n785), .A2(new_n304), .B1(new_n775), .B2(new_n1067), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n264), .B1(new_n769), .B2(new_n234), .C1(new_n773), .C2(new_n228), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(new_n299), .C2(new_n783), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1070), .B1(new_n201), .B2(new_n764), .C1(new_n222), .C2(new_n779), .ZN(new_n1071));
  OR3_X1    g0871(.A1(new_n806), .A2(KEYINPUT117), .A3(new_n413), .ZN(new_n1072));
  OAI21_X1  g0872(.A(KEYINPUT117), .B1(new_n806), .B2(new_n413), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1071), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n780), .A2(G303), .B1(G311), .B2(new_n783), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n792), .A2(G322), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1075), .B(new_n1076), .C1(new_n765), .C2(new_n974), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT48), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n797), .A2(G283), .B1(new_n772), .B2(G294), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT49), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n320), .B1(new_n775), .B2(new_n805), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G116), .B2(new_n843), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1074), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n752), .B1(new_n956), .B2(new_n1066), .C1(new_n1086), .C2(new_n757), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n696), .B2(new_n814), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1057), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1019), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1018), .A2(new_n745), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1090), .A2(new_n704), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1089), .A2(new_n1092), .ZN(G393));
  NAND2_X1  g0893(.A1(new_n1021), .A2(new_n697), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1094), .A2(new_n1016), .A3(new_n983), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n253), .A2(new_n817), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n815), .B1(new_n234), .B2(new_n211), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n752), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n803), .A2(G159), .B1(new_n792), .B2(G150), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(KEYINPUT118), .B(KEYINPUT51), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n780), .A2(new_n299), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n797), .A2(G77), .B1(new_n776), .B2(G143), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n320), .B1(new_n772), .B2(G68), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1104), .B(new_n1105), .C1(new_n504), .C2(new_n769), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(G50), .B2(new_n783), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .A4(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n783), .A2(G303), .B1(G116), .B2(new_n797), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n779), .B2(new_n535), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT120), .Z(new_n1111));
  NAND2_X1  g0911(.A1(new_n776), .A2(G322), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n264), .B1(new_n772), .B2(G283), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1111), .A2(new_n771), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n803), .A2(G311), .B1(new_n792), .B2(G317), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(KEYINPUT119), .B(KEYINPUT52), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1115), .B(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1108), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1098), .B1(new_n1118), .B2(new_n756), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n1030), .B2(new_n828), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1095), .A2(new_n1120), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1094), .A2(new_n1016), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n705), .B1(new_n1123), .B2(new_n1090), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1121), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(G390));
  NAND2_X1  g0926(.A1(new_n897), .A2(new_n907), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n812), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n838), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n752), .B1(new_n299), .B2(new_n1129), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n780), .A2(G97), .B1(new_n803), .B2(G116), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n785), .A2(new_n228), .B1(new_n775), .B2(new_n535), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n320), .B1(new_n769), .B2(new_n222), .C1(new_n773), .C2(new_n504), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1132), .B(new_n1133), .C1(G107), .C2(new_n783), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1131), .B(new_n1134), .C1(new_n799), .C2(new_n806), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n773), .A2(new_n1067), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT53), .Z(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(new_n803), .B2(G132), .ZN(new_n1138));
  INV_X1    g0938(.A(G125), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n264), .B1(new_n769), .B2(new_n201), .C1(new_n1139), .C2(new_n775), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT124), .Z(new_n1141));
  INV_X1    g0941(.A(G128), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1138), .B(new_n1141), .C1(new_n1142), .C2(new_n806), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n783), .A2(G137), .B1(G159), .B2(new_n797), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(KEYINPUT54), .B(G143), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1144), .B1(new_n779), .B2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT123), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1135), .B1(new_n1143), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1130), .B1(new_n1148), .B2(new_n756), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1128), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n916), .A2(new_n918), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n914), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n898), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1127), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n742), .A2(new_n743), .A3(new_n834), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1156), .A2(new_n915), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n718), .A2(new_n693), .A3(new_n834), .ZN(new_n1159));
  AND2_X1   g0959(.A1(new_n1159), .A2(new_n918), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1153), .B(new_n895), .C1(new_n1160), .C2(new_n915), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1155), .A2(new_n1158), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n740), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n928), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n897), .A2(new_n907), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n882), .A2(new_n888), .A3(new_n894), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n915), .B1(new_n1159), .B2(new_n918), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n1167), .A2(new_n1168), .A3(new_n898), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1165), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1162), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1150), .B1(new_n1171), .B2(new_n1055), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1163), .A2(new_n641), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n923), .A2(new_n677), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(KEYINPUT121), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT121), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n923), .A2(new_n1176), .A3(new_n677), .A4(new_n1173), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1151), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1156), .A2(new_n915), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1165), .B1(new_n1181), .B2(KEYINPUT122), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT122), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1156), .A2(new_n1183), .A3(new_n915), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1180), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n915), .B1(new_n740), .B2(new_n927), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1160), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1157), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1179), .B1(new_n1185), .B2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n705), .B1(new_n1189), .B2(new_n1171), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1188), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n1156), .A2(new_n1183), .A3(new_n915), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1183), .B1(new_n1156), .B2(new_n915), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1192), .A2(new_n1193), .A3(new_n1165), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1191), .B1(new_n1194), .B2(new_n1180), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1164), .B1(new_n1155), .B2(new_n1161), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n1166), .A2(new_n1169), .A3(new_n1157), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1195), .A2(new_n1198), .A3(new_n1179), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1172), .B1(new_n1190), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(G378));
  AOI21_X1  g1001(.A(new_n929), .B1(new_n906), .B2(new_n882), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n935), .B(G330), .C1(new_n1202), .C2(KEYINPUT40), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n345), .A2(new_n297), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n867), .A2(new_n296), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1204), .B(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1206), .B(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1203), .A2(new_n1209), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n933), .A2(G330), .A3(new_n935), .A4(new_n1208), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n922), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n922), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1209), .A2(new_n812), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n752), .B1(G50), .B2(new_n1129), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n202), .A2(new_n769), .B1(new_n775), .B2(new_n799), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n264), .A2(G41), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n773), .B2(new_n228), .C1(new_n222), .C2(new_n785), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1219), .B(new_n1221), .C1(G97), .C2(new_n783), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n780), .A2(new_n305), .B1(new_n803), .B2(G107), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1222), .B(new_n1223), .C1(new_n465), .C2(new_n806), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT58), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1220), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1227), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n797), .A2(G150), .ZN(new_n1230));
  INV_X1    g1030(.A(G132), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1230), .B1(new_n773), .B2(new_n1145), .C1(new_n784), .C2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(G137), .B2(new_n780), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n1139), .B2(new_n806), .C1(new_n1142), .C2(new_n764), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT125), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(KEYINPUT59), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n843), .A2(G159), .ZN(new_n1237));
  AOI211_X1 g1037(.A(G33), .B(G41), .C1(new_n776), .C2(G124), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1235), .A2(KEYINPUT59), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n1229), .B1(new_n1225), .B2(new_n1224), .C1(new_n1239), .C2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1218), .B1(new_n1241), .B2(new_n756), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1216), .A2(new_n983), .B1(new_n1217), .B2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1178), .B1(new_n1195), .B2(new_n1198), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n922), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n1210), .A2(new_n1211), .B1(new_n908), .B2(new_n921), .ZN(new_n1246));
  OAI21_X1  g1046(.A(KEYINPUT57), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n704), .B1(new_n1244), .B2(new_n1247), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n739), .A2(KEYINPUT93), .A3(G330), .ZN(new_n1249));
  AOI21_X1  g1049(.A(KEYINPUT93), .B1(new_n739), .B2(G330), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1249), .A2(new_n1250), .A3(new_n927), .ZN(new_n1251));
  OAI21_X1  g1051(.A(KEYINPUT122), .B1(new_n1251), .B2(new_n914), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1252), .A2(new_n1164), .A3(new_n1184), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1188), .B1(new_n1253), .B2(new_n1151), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1179), .B1(new_n1254), .B2(new_n1171), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT57), .B1(new_n1255), .B2(new_n1216), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1243), .B1(new_n1248), .B2(new_n1256), .ZN(G375));
  OAI211_X1 g1057(.A(new_n1178), .B(new_n1191), .C1(new_n1194), .C2(new_n1180), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1189), .A2(new_n1258), .A3(new_n1025), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n915), .A2(new_n812), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n752), .B1(G68), .B2(new_n1129), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n784), .A2(new_n1145), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n797), .A2(G50), .B1(new_n776), .B2(G128), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n320), .B1(new_n772), .B2(G159), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1263), .B(new_n1264), .C1(new_n202), .C2(new_n769), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n1262), .B(new_n1265), .C1(G150), .C2(new_n780), .ZN(new_n1266));
  OAI221_X1 g1066(.A(new_n1266), .B1(new_n1231), .B2(new_n806), .C1(new_n848), .C2(new_n765), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n780), .A2(G107), .B1(new_n803), .B2(G283), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n785), .A2(new_n304), .B1(new_n775), .B2(new_n488), .ZN(new_n1269));
  OAI221_X1 g1069(.A(new_n320), .B1(new_n769), .B2(new_n228), .C1(new_n773), .C2(new_n234), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n1269), .B(new_n1270), .C1(G116), .C2(new_n783), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1268), .B(new_n1271), .C1(new_n535), .C2(new_n806), .ZN(new_n1272));
  OR2_X1    g1072(.A1(new_n1272), .A2(KEYINPUT126), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(KEYINPUT126), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1267), .A2(new_n1273), .A3(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1261), .B1(new_n1275), .B2(new_n756), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n1195), .A2(new_n983), .B1(new_n1260), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1259), .A2(new_n1277), .ZN(G381));
  OAI211_X1 g1078(.A(new_n1125), .B(new_n982), .C1(new_n1026), .C2(new_n1053), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(G375), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1089), .A2(new_n830), .A3(new_n1092), .ZN(new_n1282));
  NOR3_X1   g1082(.A1(new_n1282), .A2(G384), .A3(G381), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1280), .A2(new_n1200), .A3(new_n1281), .A4(new_n1283), .ZN(G407));
  NAND2_X1  g1084(.A1(new_n1200), .A2(new_n683), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G407), .B(G213), .C1(G375), .C2(new_n1285), .ZN(G409));
  NAND3_X1  g1086(.A1(new_n1255), .A2(new_n1025), .A3(new_n1216), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1243), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1200), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1289), .B1(G375), .B2(new_n1200), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n683), .A2(G213), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1254), .A2(KEYINPUT60), .A3(new_n1178), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1293), .A2(new_n704), .A3(new_n1189), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT60), .B1(new_n1254), .B2(new_n1178), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1277), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(G384), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  OAI211_X1 g1098(.A(G384), .B(new_n1277), .C1(new_n1294), .C2(new_n1295), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n683), .A2(G213), .A3(G2897), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(KEYINPUT127), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT127), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1298), .A2(new_n1303), .A3(new_n1299), .A4(new_n1300), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1300), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1292), .A2(new_n1302), .A3(new_n1304), .A4(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1299), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT60), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1258), .A2(new_n1310), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1311), .A2(new_n704), .A3(new_n1189), .A4(new_n1293), .ZN(new_n1312));
  AOI21_X1  g1112(.A(G384), .B1(new_n1312), .B2(new_n1277), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1309), .A2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1290), .A2(new_n1291), .A3(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(KEYINPUT62), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT61), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT62), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1290), .A2(new_n1314), .A3(new_n1318), .A4(new_n1291), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1308), .A2(new_n1316), .A3(new_n1317), .A4(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(G393), .A2(G396), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1282), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(G387), .A2(G390), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1322), .B1(new_n1323), .B2(new_n1279), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1323), .A2(new_n1279), .A3(new_n1322), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1320), .A2(new_n1327), .ZN(new_n1328));
  AND3_X1   g1128(.A1(new_n1323), .A2(new_n1279), .A3(new_n1322), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1329), .A2(new_n1324), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1315), .A2(KEYINPUT63), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT63), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1290), .A2(new_n1314), .A3(new_n1332), .A4(new_n1291), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1331), .A2(new_n1333), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1330), .A2(new_n1334), .A3(new_n1317), .A4(new_n1308), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1328), .A2(new_n1335), .ZN(G405));
  NAND2_X1  g1136(.A1(new_n1281), .A2(G378), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(G375), .A2(new_n1200), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(new_n1314), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1337), .A2(new_n1305), .A3(new_n1338), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1330), .A2(new_n1340), .A3(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1327), .A2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1342), .A2(new_n1344), .ZN(G402));
endmodule


