//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1 0 1 0 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n814, new_n816, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OR2_X1    g003(.A1(new_n204), .A2(KEYINPUT90), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n202), .A2(G1gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(KEYINPUT90), .ZN(new_n207));
  XNOR2_X1  g006(.A(KEYINPUT91), .B(G8gat), .ZN(new_n208));
  NAND4_X1  g007(.A1(new_n205), .A2(new_n206), .A3(new_n207), .A4(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n206), .A2(new_n204), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G8gat), .ZN(new_n211));
  AND2_X1   g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT21), .ZN(new_n213));
  XOR2_X1   g012(.A(G57gat), .B(G64gat), .Z(new_n214));
  INV_X1    g013(.A(KEYINPUT9), .ZN(new_n215));
  INV_X1    g014(.A(G71gat), .ZN(new_n216));
  INV_X1    g015(.A(G78gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  XOR2_X1   g018(.A(G71gat), .B(G78gat), .Z(new_n220));
  OR2_X1    g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n220), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n212), .B1(new_n213), .B2(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(new_n224), .B(KEYINPUT100), .Z(new_n225));
  AOI21_X1  g024(.A(KEYINPUT21), .B1(new_n221), .B2(new_n222), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n226), .B(KEYINPUT98), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n227), .B(KEYINPUT99), .ZN(new_n228));
  XOR2_X1   g027(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n228), .A2(new_n230), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n225), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n233), .ZN(new_n235));
  INV_X1    g034(.A(new_n225), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(new_n231), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G127gat), .B(G155gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(G231gat), .A2(G233gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G183gat), .B(G211gat), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n241), .B(new_n242), .Z(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n238), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n234), .A2(new_n237), .A3(new_n243), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G120gat), .B(G148gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(G176gat), .B(G204gat), .ZN(new_n249));
  XOR2_X1   g048(.A(new_n248), .B(new_n249), .Z(new_n250));
  NAND2_X1  g049(.A1(G230gat), .A2(G233gat), .ZN(new_n251));
  INV_X1    g050(.A(G85gat), .ZN(new_n252));
  INV_X1    g051(.A(G92gat), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT102), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT102), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(G85gat), .A3(G92gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n254), .A2(new_n256), .A3(KEYINPUT7), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT7), .ZN(new_n258));
  OAI211_X1 g057(.A(KEYINPUT102), .B(new_n258), .C1(new_n252), .C2(new_n253), .ZN(new_n259));
  NAND2_X1  g058(.A1(G99gat), .A2(G106gat), .ZN(new_n260));
  AOI22_X1  g059(.A1(KEYINPUT8), .A2(new_n260), .B1(new_n252), .B2(new_n253), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n257), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(G99gat), .B(G106gat), .Z(new_n263));
  OR2_X1    g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n263), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(new_n223), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n264), .A2(new_n222), .A3(new_n221), .A4(new_n265), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n251), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n250), .B1(new_n270), .B2(KEYINPUT105), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n271), .B1(KEYINPUT105), .B2(new_n270), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT10), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n267), .A2(new_n273), .A3(new_n268), .ZN(new_n274));
  OR2_X1    g073(.A1(new_n268), .A2(new_n273), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(new_n251), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n272), .A2(new_n277), .ZN(new_n278));
  OR2_X1    g077(.A1(new_n277), .A2(KEYINPUT106), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(KEYINPUT106), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n269), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n278), .B1(new_n281), .B2(new_n250), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT88), .ZN(new_n284));
  INV_X1    g083(.A(G29gat), .ZN(new_n285));
  INV_X1    g084(.A(G36gat), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT14), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT14), .ZN(new_n288));
  NOR3_X1   g087(.A1(new_n288), .A2(G29gat), .A3(G36gat), .ZN(new_n289));
  AOI211_X1 g088(.A(new_n287), .B(new_n289), .C1(G29gat), .C2(G36gat), .ZN(new_n290));
  INV_X1    g089(.A(G43gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(G50gat), .ZN(new_n292));
  INV_X1    g091(.A(G50gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G43gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n292), .A2(new_n294), .A3(KEYINPUT15), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n284), .B1(new_n290), .B2(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(KEYINPUT86), .B(KEYINPUT15), .Z(new_n297));
  INV_X1    g096(.A(new_n294), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n292), .B1(new_n298), .B2(KEYINPUT87), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT87), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n297), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n302), .A2(new_n290), .A3(new_n295), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n296), .A2(new_n303), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n302), .A2(new_n290), .A3(new_n284), .A4(new_n295), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(KEYINPUT17), .A3(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n306), .B(KEYINPUT92), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n304), .A2(new_n305), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT89), .B1(new_n309), .B2(KEYINPUT17), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT89), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT17), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n308), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n307), .A2(new_n310), .A3(new_n313), .A4(new_n266), .ZN(new_n314));
  OR2_X1    g113(.A1(new_n314), .A2(KEYINPUT103), .ZN(new_n315));
  NAND2_X1  g114(.A1(G232gat), .A2(G233gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT41), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n318), .B1(new_n309), .B2(new_n266), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n319), .B1(new_n314), .B2(KEYINPUT103), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  XOR2_X1   g120(.A(G190gat), .B(G218gat), .Z(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n317), .A2(KEYINPUT41), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n324), .B(KEYINPUT101), .ZN(new_n325));
  XOR2_X1   g124(.A(G134gat), .B(G162gat), .Z(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n328), .A2(KEYINPUT104), .ZN(new_n329));
  INV_X1    g128(.A(new_n322), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n315), .A2(new_n320), .A3(new_n330), .ZN(new_n331));
  AND3_X1   g130(.A1(new_n323), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n327), .B(KEYINPUT104), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n334), .B1(new_n323), .B2(new_n331), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n247), .B(new_n283), .C1(new_n332), .C2(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(KEYINPUT93), .B(KEYINPUT18), .Z(new_n337));
  NAND4_X1  g136(.A1(new_n307), .A2(new_n310), .A3(new_n313), .A4(new_n212), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n209), .A2(new_n211), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n308), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G229gat), .A2(G233gat), .ZN(new_n341));
  AND2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n337), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT97), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n338), .A2(KEYINPUT18), .A3(new_n342), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n212), .A2(new_n304), .A3(new_n305), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT94), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n346), .A2(new_n340), .A3(new_n347), .ZN(new_n348));
  XOR2_X1   g147(.A(new_n341), .B(KEYINPUT13), .Z(new_n349));
  NAND3_X1  g148(.A1(new_n308), .A2(KEYINPUT94), .A3(new_n339), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT95), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n351), .B(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n344), .A2(new_n345), .A3(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G113gat), .B(G141gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(G197gat), .ZN(new_n356));
  XOR2_X1   g155(.A(KEYINPUT11), .B(G169gat), .Z(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  XOR2_X1   g157(.A(new_n358), .B(KEYINPUT12), .Z(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n360), .B1(new_n343), .B2(KEYINPUT97), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n354), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n343), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n363), .A2(new_n353), .A3(new_n345), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n359), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT96), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n364), .A2(KEYINPUT96), .A3(new_n359), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n362), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n336), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(G228gat), .A2(G233gat), .ZN(new_n371));
  AND2_X1   g170(.A1(G155gat), .A2(G162gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(G155gat), .A2(G162gat), .ZN(new_n373));
  OR2_X1    g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(G141gat), .ZN(new_n375));
  INV_X1    g174(.A(G148gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(G141gat), .A2(G148gat), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(G162gat), .ZN(new_n380));
  OR2_X1    g179(.A1(KEYINPUT75), .A2(G155gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(KEYINPUT75), .A2(G155gat), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT2), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n374), .B(new_n379), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT74), .B1(new_n372), .B2(new_n373), .ZN(new_n386));
  OR2_X1    g185(.A1(new_n373), .A2(KEYINPUT74), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n377), .A2(new_n384), .A3(new_n378), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G197gat), .B(G204gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(G211gat), .A2(G218gat), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT22), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(G211gat), .ZN(new_n396));
  INV_X1    g195(.A(G218gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n395), .A2(new_n392), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n392), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n400), .A2(new_n391), .A3(new_n394), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT29), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n390), .B1(new_n402), .B2(KEYINPUT3), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT80), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n371), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n403), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n399), .A2(new_n401), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT3), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n385), .A2(new_n408), .A3(new_n389), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT29), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n407), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n405), .B1(new_n406), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n411), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n413), .B(new_n403), .C1(new_n404), .C2(new_n371), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(G22gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n412), .A2(new_n414), .A3(G22gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G78gat), .B(G106gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(KEYINPUT31), .B(G50gat), .ZN(new_n421));
  XOR2_X1   g220(.A(new_n420), .B(new_n421), .Z(new_n422));
  AOI21_X1  g221(.A(G22gat), .B1(new_n412), .B2(new_n414), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT81), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n417), .A2(new_n424), .A3(new_n418), .A4(new_n422), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT36), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT70), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT1), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n431), .B1(G113gat), .B2(G120gat), .ZN(new_n432));
  AND2_X1   g231(.A1(G113gat), .A2(G120gat), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n430), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(G127gat), .B(G134gat), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n435), .B(new_n430), .C1(new_n433), .C2(new_n432), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT25), .ZN(new_n440));
  NAND2_X1  g239(.A1(G169gat), .A2(G176gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT23), .ZN(new_n442));
  INV_X1    g241(.A(G169gat), .ZN(new_n443));
  INV_X1    g242(.A(G176gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n440), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n443), .A2(new_n444), .A3(KEYINPUT67), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT67), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n448), .B1(G169gat), .B2(G176gat), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n449), .A3(KEYINPUT23), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT68), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(G183gat), .A2(G190gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n452), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n451), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n455), .A2(new_n452), .A3(new_n456), .ZN(new_n459));
  NAND4_X1  g258(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT65), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n455), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n442), .A2(new_n445), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT23), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n465), .A2(G176gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n443), .A2(KEYINPUT66), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT66), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(G169gat), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n466), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n463), .A2(new_n464), .A3(new_n470), .ZN(new_n471));
  AOI22_X1  g270(.A1(new_n458), .A2(new_n459), .B1(new_n440), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(KEYINPUT27), .B(G183gat), .ZN(new_n473));
  INV_X1    g272(.A(G190gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT69), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT28), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n475), .A2(new_n478), .B1(G183gat), .B2(G190gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n445), .A2(KEYINPUT26), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n447), .A2(new_n449), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n441), .B(new_n480), .C1(new_n481), .C2(KEYINPUT26), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n473), .A2(new_n476), .A3(new_n477), .A4(new_n474), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n479), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n439), .B1(new_n472), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(G227gat), .A2(G233gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(KEYINPUT64), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n455), .A2(new_n456), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT68), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n489), .A2(new_n459), .A3(new_n450), .A4(new_n446), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n455), .A2(new_n460), .A3(new_n462), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n470), .A2(new_n464), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n440), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n439), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n479), .A2(new_n482), .A3(new_n483), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n485), .A2(new_n487), .A3(new_n497), .ZN(new_n498));
  XOR2_X1   g297(.A(G71gat), .B(G99gat), .Z(new_n499));
  XNOR2_X1  g298(.A(G15gat), .B(G43gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT33), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n498), .A2(KEYINPUT32), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT71), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n498), .A2(KEYINPUT71), .A3(KEYINPUT32), .A4(new_n502), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n485), .A2(new_n497), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT34), .ZN(new_n509));
  INV_X1    g308(.A(new_n487), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n509), .B1(new_n508), .B2(new_n510), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n498), .A2(KEYINPUT32), .ZN(new_n515));
  INV_X1    g314(.A(new_n498), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n515), .B(new_n501), .C1(new_n516), .C2(KEYINPUT33), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n507), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n514), .B1(new_n507), .B2(new_n517), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n429), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n507), .A2(new_n517), .ZN(new_n521));
  INV_X1    g320(.A(new_n514), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n514), .A3(new_n517), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(KEYINPUT36), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n428), .B1(new_n520), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT85), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT37), .ZN(new_n528));
  NAND2_X1  g327(.A1(G226gat), .A2(G233gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT72), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n494), .A2(new_n496), .A3(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n530), .A2(KEYINPUT29), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n533), .B1(new_n494), .B2(new_n496), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n407), .B1(new_n531), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n532), .B1(new_n472), .B2(new_n484), .ZN(new_n536));
  INV_X1    g335(.A(new_n407), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n494), .A2(new_n496), .A3(new_n530), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n528), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G8gat), .B(G36gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(G64gat), .B(G92gat), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n541), .B(new_n542), .Z(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n531), .A2(new_n534), .A3(new_n407), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n537), .B1(new_n536), .B2(new_n538), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n544), .A2(KEYINPUT37), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n540), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT38), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n527), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n539), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n544), .B1(new_n552), .B2(KEYINPUT37), .ZN(new_n553));
  OAI211_X1 g352(.A(KEYINPUT85), .B(KEYINPUT38), .C1(new_n553), .C2(new_n540), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n535), .A2(KEYINPUT84), .A3(new_n539), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n555), .B(KEYINPUT37), .C1(KEYINPUT84), .C2(new_n535), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n547), .A2(new_n548), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n550), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n535), .A2(new_n539), .A3(new_n543), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G1gat), .B(G29gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT0), .ZN(new_n562));
  XNOR2_X1  g361(.A(G57gat), .B(G85gat), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n562), .B(new_n563), .Z(new_n564));
  OAI211_X1 g363(.A(new_n377), .B(new_n378), .C1(new_n372), .C2(new_n373), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n381), .A2(new_n382), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(G162gat), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n565), .B1(new_n567), .B2(KEYINPUT2), .ZN(new_n568));
  AND3_X1   g367(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT3), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n570), .A2(new_n495), .A3(new_n409), .ZN(new_n571));
  NAND2_X1  g370(.A1(G225gat), .A2(G233gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n573), .A2(KEYINPUT5), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n439), .A2(new_n385), .A3(new_n389), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT4), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT77), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT4), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n439), .A2(new_n578), .A3(new_n385), .A4(new_n389), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n577), .B1(new_n576), .B2(new_n579), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n571), .B(new_n574), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT5), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n495), .A2(new_n390), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(new_n575), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n583), .B1(new_n585), .B2(new_n573), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT76), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n576), .A2(new_n587), .A3(new_n579), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n575), .A2(KEYINPUT76), .A3(KEYINPUT4), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n589), .A2(new_n571), .A3(new_n572), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n586), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n564), .B1(new_n582), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n560), .B1(new_n592), .B2(KEYINPUT6), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n551), .A2(new_n554), .A3(new_n558), .A4(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n582), .A2(new_n591), .A3(new_n564), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT78), .ZN(new_n596));
  INV_X1    g395(.A(new_n592), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT6), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT78), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n582), .A2(new_n591), .A3(new_n599), .A4(new_n564), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n596), .A2(new_n597), .A3(new_n598), .A4(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT83), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n598), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n605), .A2(KEYINPUT83), .A3(new_n597), .A4(new_n596), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n594), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n571), .B1(new_n580), .B2(new_n581), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT39), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n608), .A2(new_n609), .A3(new_n573), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n608), .A2(new_n573), .ZN(new_n611));
  OAI21_X1  g410(.A(KEYINPUT39), .B1(new_n585), .B2(new_n573), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n564), .B(new_n610), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(KEYINPUT82), .A2(KEYINPUT40), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n560), .A2(KEYINPUT30), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT30), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n559), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT73), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n618), .A2(KEYINPUT73), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n547), .B(new_n616), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n592), .B1(new_n613), .B2(new_n614), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n615), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n526), .B1(new_n607), .B2(new_n624), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n595), .A2(KEYINPUT78), .ZN(new_n626));
  OAI21_X1  g425(.A(KEYINPUT79), .B1(new_n626), .B2(new_n604), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT79), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n596), .A2(new_n628), .A3(new_n598), .A4(new_n600), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n627), .A2(new_n597), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n592), .A2(KEYINPUT6), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n622), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n426), .A2(new_n427), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n633), .B1(new_n520), .B2(new_n525), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT35), .ZN(new_n635));
  NOR4_X1   g434(.A1(new_n428), .A2(new_n518), .A3(new_n519), .A4(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n632), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  AOI22_X1  g436(.A1(new_n603), .A2(new_n606), .B1(KEYINPUT6), .B2(new_n592), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n518), .A2(new_n519), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n616), .A2(new_n547), .ZN(new_n640));
  INV_X1    g439(.A(new_n621), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n640), .B1(new_n641), .B2(new_n619), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n633), .A2(new_n639), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n635), .B1(new_n638), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n625), .A2(new_n637), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n370), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n630), .A2(new_n631), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g449(.A(KEYINPUT16), .B(G8gat), .Z(new_n651));
  NAND3_X1  g450(.A1(new_n647), .A2(new_n622), .A3(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(G8gat), .B1(new_n646), .B2(new_n642), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  MUX2_X1   g453(.A(new_n652), .B(new_n654), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g454(.A1(new_n520), .A2(new_n525), .ZN(new_n656));
  OAI21_X1  g455(.A(G15gat), .B1(new_n646), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(G15gat), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n639), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n657), .B1(new_n646), .B2(new_n659), .ZN(G1326gat));
  NOR2_X1   g459(.A1(new_n646), .A2(new_n633), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT43), .B(G22gat), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(G1327gat));
  NOR2_X1   g462(.A1(new_n332), .A2(new_n335), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n645), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n369), .A2(new_n247), .A3(new_n282), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n668), .A2(new_n285), .A3(new_n648), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT45), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n666), .A2(KEYINPUT44), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n665), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n667), .ZN(new_n675));
  INV_X1    g474(.A(new_n648), .ZN(new_n676));
  OAI21_X1  g475(.A(G29gat), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n670), .A2(new_n677), .ZN(G1328gat));
  NAND3_X1  g477(.A1(new_n668), .A2(new_n286), .A3(new_n622), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n679), .B(KEYINPUT46), .Z(new_n680));
  OAI21_X1  g479(.A(G36gat), .B1(new_n675), .B2(new_n642), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(G1329gat));
  NAND2_X1  g481(.A1(new_n668), .A2(new_n639), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT107), .ZN(new_n684));
  AOI22_X1  g483(.A1(new_n683), .A2(new_n291), .B1(new_n684), .B2(KEYINPUT47), .ZN(new_n685));
  INV_X1    g484(.A(new_n656), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n674), .A2(G43gat), .A3(new_n686), .A4(new_n667), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n684), .A2(KEYINPUT47), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n685), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n688), .B1(new_n685), .B2(new_n687), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(G1330gat));
  NAND4_X1  g490(.A1(new_n671), .A2(new_n428), .A3(new_n673), .A4(new_n667), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(G50gat), .ZN(new_n693));
  NOR2_X1   g492(.A1(KEYINPUT108), .A2(KEYINPUT48), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n633), .A2(G50gat), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n694), .B1(new_n668), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(KEYINPUT108), .A2(KEYINPUT48), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT109), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n697), .B(new_n699), .ZN(G1331gat));
  OR2_X1    g499(.A1(new_n354), .A2(new_n361), .ZN(new_n701));
  INV_X1    g500(.A(new_n368), .ZN(new_n702));
  AOI21_X1  g501(.A(KEYINPUT96), .B1(new_n364), .B2(new_n359), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n247), .ZN(new_n705));
  NOR4_X1   g504(.A1(new_n704), .A2(new_n664), .A3(new_n705), .A4(new_n283), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n645), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n648), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g509(.A1(new_n707), .A2(new_n642), .ZN(new_n711));
  NOR2_X1   g510(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n712));
  AND2_X1   g511(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n714), .B1(new_n711), .B2(new_n712), .ZN(G1333gat));
  OAI21_X1  g514(.A(G71gat), .B1(new_n707), .B2(new_n656), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n639), .A2(new_n216), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(new_n707), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1334gat));
  NOR2_X1   g519(.A1(new_n707), .A2(new_n633), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(new_n217), .ZN(G1335gat));
  NAND2_X1  g521(.A1(new_n369), .A2(new_n705), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n723), .A2(new_n283), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n671), .A2(new_n673), .A3(new_n724), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n725), .A2(new_n648), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT51), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n645), .A2(KEYINPUT111), .A3(new_n664), .ZN(new_n728));
  INV_X1    g527(.A(new_n723), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT111), .B1(new_n645), .B2(new_n664), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n727), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT111), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n665), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n734), .A2(KEYINPUT51), .A3(new_n729), .A4(new_n728), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n648), .A2(new_n252), .A3(new_n282), .ZN(new_n738));
  OAI22_X1  g537(.A1(new_n726), .A2(new_n252), .B1(new_n737), .B2(new_n738), .ZN(G1336gat));
  INV_X1    g538(.A(KEYINPUT112), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n732), .A2(new_n740), .A3(new_n735), .ZN(new_n741));
  OAI211_X1 g540(.A(KEYINPUT112), .B(new_n727), .C1(new_n730), .C2(new_n731), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n283), .A2(G92gat), .A3(new_n642), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n671), .A2(new_n622), .A3(new_n673), .A4(new_n724), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G92gat), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT52), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n736), .A2(new_n743), .ZN(new_n749));
  XOR2_X1   g548(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n750));
  NAND3_X1  g549(.A1(new_n749), .A2(new_n746), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n748), .A2(new_n751), .ZN(G1337gat));
  INV_X1    g551(.A(KEYINPUT114), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n283), .A2(G99gat), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n736), .A2(new_n639), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(G99gat), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n757), .B1(new_n725), .B2(new_n686), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n753), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n725), .A2(new_n686), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n755), .B(KEYINPUT114), .C1(new_n760), .C2(new_n757), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(G1338gat));
  NOR3_X1   g561(.A1(new_n283), .A2(G106gat), .A3(new_n633), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n741), .A2(new_n742), .A3(new_n763), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n671), .A2(new_n428), .A3(new_n673), .A4(new_n724), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G106gat), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(KEYINPUT53), .ZN(new_n768));
  XNOR2_X1  g567(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT115), .B1(new_n736), .B2(new_n763), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT115), .ZN(new_n771));
  INV_X1    g570(.A(new_n763), .ZN(new_n772));
  AOI211_X1 g571(.A(new_n771), .B(new_n772), .C1(new_n732), .C2(new_n735), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n766), .B(new_n769), .C1(new_n770), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n768), .A2(new_n774), .ZN(G1339gat));
  NAND2_X1  g574(.A1(new_n323), .A2(new_n331), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n333), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n323), .A2(new_n329), .A3(new_n331), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n369), .A2(new_n779), .A3(new_n247), .A4(new_n283), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n341), .B1(new_n338), .B2(new_n340), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n349), .B1(new_n348), .B2(new_n350), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n358), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n282), .B(new_n783), .C1(new_n354), .C2(new_n361), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n332), .B2(new_n335), .ZN(new_n785));
  INV_X1    g584(.A(new_n278), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n274), .A2(new_n275), .A3(G230gat), .A4(G233gat), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT117), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n789), .A2(KEYINPUT54), .A3(new_n277), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n279), .A2(new_n791), .A3(new_n280), .ZN(new_n792));
  INV_X1    g591(.A(new_n250), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n790), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n786), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n790), .A2(new_n792), .A3(KEYINPUT55), .A4(new_n793), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n785), .B1(new_n704), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n783), .B1(new_n354), .B2(new_n361), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n705), .B1(new_n802), .B2(new_n779), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n780), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n622), .A2(new_n519), .A3(new_n518), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n804), .A2(new_n648), .A3(new_n633), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n369), .A2(G113gat), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT118), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(G113gat), .B1(new_n806), .B2(new_n369), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n811), .B(new_n812), .ZN(G1340gat));
  NOR2_X1   g612(.A1(new_n806), .A2(new_n283), .ZN(new_n814));
  XOR2_X1   g613(.A(new_n814), .B(G120gat), .Z(G1341gat));
  NOR2_X1   g614(.A1(new_n806), .A2(new_n705), .ZN(new_n816));
  XOR2_X1   g615(.A(new_n816), .B(G127gat), .Z(G1342gat));
  NOR2_X1   g616(.A1(new_n336), .A2(new_n704), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n779), .B(new_n784), .C1(new_n369), .C2(new_n798), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n701), .A2(new_n797), .A3(new_n796), .A4(new_n783), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n247), .B1(new_n820), .B2(new_n664), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n818), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n822), .A2(new_n428), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n823), .A2(new_n648), .A3(new_n639), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n664), .A2(new_n642), .ZN(new_n825));
  XOR2_X1   g624(.A(new_n825), .B(KEYINPUT120), .Z(new_n826));
  INV_X1    g625(.A(G134gat), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OR3_X1    g627(.A1(new_n824), .A2(KEYINPUT56), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(G134gat), .B1(new_n824), .B2(new_n825), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT56), .B1(new_n824), .B2(new_n828), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(G1343gat));
  NOR3_X1   g631(.A1(new_n676), .A2(new_n622), .A3(new_n686), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n369), .A2(new_n375), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n822), .A2(new_n835), .A3(new_n633), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT57), .B1(new_n804), .B2(new_n428), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n833), .B(new_n834), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n839));
  NOR2_X1   g638(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n648), .B1(new_n634), .B2(KEYINPUT121), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n841), .B1(KEYINPUT121), .B2(new_n634), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n804), .A2(new_n842), .A3(new_n642), .A4(new_n704), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n840), .B1(new_n843), .B2(new_n375), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n838), .A2(new_n839), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n839), .B1(new_n838), .B2(new_n844), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(G1344gat));
  AND2_X1   g646(.A1(new_n804), .A2(new_n842), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n848), .A2(new_n642), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n849), .A2(new_n376), .A3(new_n282), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n282), .B(new_n833), .C1(new_n836), .C2(new_n837), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n851), .A2(new_n852), .A3(G148gat), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n851), .B2(G148gat), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n850), .B1(new_n853), .B2(new_n854), .ZN(G1345gat));
  AOI21_X1  g654(.A(new_n566), .B1(new_n849), .B2(new_n247), .ZN(new_n856));
  INV_X1    g655(.A(new_n833), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n835), .B1(new_n822), .B2(new_n633), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n804), .A2(KEYINPUT57), .A3(new_n428), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n247), .A2(new_n566), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n861), .B(KEYINPUT123), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n856), .B1(new_n860), .B2(new_n862), .ZN(G1346gat));
  NAND3_X1  g662(.A1(new_n848), .A2(new_n380), .A3(new_n826), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n860), .A2(new_n664), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(new_n865), .B2(new_n380), .ZN(G1347gat));
  NOR2_X1   g665(.A1(new_n822), .A2(new_n648), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n639), .A2(new_n633), .A3(new_n622), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n869), .A2(new_n467), .A3(new_n469), .A4(new_n704), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n648), .A2(new_n642), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n639), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT124), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n823), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(G169gat), .B1(new_n874), .B2(new_n369), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n870), .A2(new_n875), .ZN(G1348gat));
  NAND3_X1  g675(.A1(new_n869), .A2(new_n444), .A3(new_n282), .ZN(new_n877));
  OAI21_X1  g676(.A(G176gat), .B1(new_n874), .B2(new_n283), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(G1349gat));
  OAI21_X1  g678(.A(G183gat), .B1(new_n874), .B2(new_n705), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n867), .A2(new_n473), .A3(new_n247), .A4(new_n868), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n880), .A2(new_n883), .A3(new_n881), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(G1350gat));
  NAND3_X1  g686(.A1(new_n869), .A2(new_n474), .A3(new_n664), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT126), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n823), .A2(new_n664), .A3(new_n873), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT61), .ZN(new_n891));
  AND4_X1   g690(.A1(new_n889), .A2(new_n890), .A3(new_n891), .A4(G190gat), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n474), .B1(KEYINPUT126), .B2(KEYINPUT61), .ZN(new_n893));
  AOI22_X1  g692(.A1(new_n890), .A2(new_n893), .B1(new_n889), .B2(new_n891), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n888), .B1(new_n892), .B2(new_n894), .ZN(G1351gat));
  AND2_X1   g694(.A1(new_n634), .A2(new_n622), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n867), .A2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(G197gat), .B1(new_n898), .B2(new_n704), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n871), .A2(new_n656), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n900), .B1(new_n858), .B2(new_n859), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n704), .A2(G197gat), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(G1352gat));
  INV_X1    g702(.A(G204gat), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n867), .A2(new_n904), .A3(new_n282), .A4(new_n896), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT62), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n905), .A2(KEYINPUT62), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n901), .A2(new_n282), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n906), .B(new_n907), .C1(new_n908), .C2(new_n904), .ZN(G1353gat));
  NAND3_X1  g708(.A1(new_n898), .A2(new_n396), .A3(new_n247), .ZN(new_n910));
  INV_X1    g709(.A(new_n900), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n247), .B(new_n911), .C1(new_n836), .C2(new_n837), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n912), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT63), .B1(new_n912), .B2(G211gat), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n910), .B1(new_n913), .B2(new_n914), .ZN(G1354gat));
  OAI21_X1  g714(.A(new_n397), .B1(new_n897), .B2(new_n779), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g717(.A(KEYINPUT127), .B(new_n397), .C1(new_n897), .C2(new_n779), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n779), .A2(new_n397), .ZN(new_n920));
  AOI22_X1  g719(.A1(new_n918), .A2(new_n919), .B1(new_n901), .B2(new_n920), .ZN(G1355gat));
endmodule


