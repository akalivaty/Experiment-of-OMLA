//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 1 0 1 0 1 0 1 0 1 0 0 1 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI21_X1  g0005(.A(G50), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  AND2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  XNOR2_X1  g0010(.A(KEYINPUT66), .B(G244), .ZN(new_n211));
  AND2_X1   g0011(.A1(new_n211), .A2(G77), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G107), .A2(G264), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n210), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT1), .Z(new_n219));
  INV_X1    g0019(.A(new_n210), .ZN(new_n220));
  INV_X1    g0020(.A(G13), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n220), .A2(KEYINPUT65), .A3(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT65), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n223), .B1(new_n210), .B2(G13), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  INV_X1    g0026(.A(KEYINPUT0), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n204), .A2(new_n205), .ZN(new_n231));
  INV_X1    g0031(.A(G50), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI22_X1  g0033(.A1(new_n226), .A2(new_n227), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n219), .B(new_n234), .C1(new_n227), .C2(new_n226), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(KEYINPUT67), .Z(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G226), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n239), .B(G232), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  NOR2_X1   g0051(.A1(G41), .A2(G45), .ZN(new_n252));
  INV_X1    g0052(.A(G274), .ZN(new_n253));
  NOR3_X1   g0053(.A1(new_n252), .A2(G1), .A3(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n255), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G223), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(new_n259), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(G222), .A3(new_n255), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n261), .B(new_n263), .C1(new_n207), .C2(new_n262), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n254), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(KEYINPUT68), .A2(G1), .ZN(new_n267));
  NOR2_X1   g0067(.A1(KEYINPUT68), .A2(G1), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n267), .A2(new_n252), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT69), .ZN(new_n270));
  NOR3_X1   g0070(.A1(new_n269), .A2(new_n270), .A3(new_n265), .ZN(new_n271));
  INV_X1    g0071(.A(new_n252), .ZN(new_n272));
  OR2_X1    g0072(.A1(KEYINPUT68), .A2(G1), .ZN(new_n273));
  NAND2_X1  g0073(.A1(KEYINPUT68), .A2(G1), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n228), .ZN(new_n276));
  INV_X1    g0076(.A(G41), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n276), .B1(new_n257), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(KEYINPUT69), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(G226), .B1(new_n271), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n266), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G200), .ZN(new_n282));
  XNOR2_X1  g0082(.A(new_n282), .B(KEYINPUT75), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT9), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n273), .A2(G13), .A3(G20), .A4(new_n274), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT71), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n267), .A2(new_n268), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT71), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n287), .A2(new_n288), .A3(G13), .A4(G20), .ZN(new_n289));
  AND2_X1   g0089(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT70), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(new_n229), .A3(G33), .ZN(new_n292));
  OAI21_X1  g0092(.A(KEYINPUT70), .B1(new_n257), .B2(G20), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n292), .B(new_n293), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G150), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n296), .B(new_n298), .C1(new_n206), .C2(new_n229), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n228), .B1(new_n210), .B2(new_n257), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n290), .A2(new_n232), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n286), .A2(new_n289), .ZN(new_n302));
  INV_X1    g0102(.A(new_n300), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n232), .B1(new_n287), .B2(G20), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(KEYINPUT74), .B1(new_n301), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n293), .A2(new_n292), .ZN(new_n307));
  XNOR2_X1  g0107(.A(KEYINPUT8), .B(G58), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n298), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n229), .B1(new_n231), .B2(new_n232), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n300), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n286), .A2(new_n289), .A3(new_n232), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n305), .A2(new_n311), .A3(KEYINPUT74), .A4(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n284), .B1(new_n306), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n305), .A2(new_n312), .A3(new_n311), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT74), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n318), .A2(KEYINPUT9), .A3(new_n313), .ZN(new_n319));
  INV_X1    g0119(.A(new_n281), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G190), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n315), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  OR3_X1    g0122(.A1(new_n283), .A2(new_n322), .A3(KEYINPUT10), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT76), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n318), .A2(new_n313), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n326), .A2(new_n284), .B1(G190), .B2(new_n320), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n327), .A2(KEYINPUT76), .A3(new_n319), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n325), .A2(new_n328), .B1(G200), .B2(new_n281), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT10), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n323), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n281), .A2(G169), .ZN(new_n332));
  INV_X1    g0132(.A(G179), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n332), .B1(new_n333), .B2(new_n281), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n316), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n302), .A2(new_n303), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT73), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n273), .A2(new_n274), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(new_n229), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n302), .A2(KEYINPUT73), .A3(new_n303), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n338), .A2(G68), .A3(new_n341), .A4(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT12), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n290), .A2(new_n344), .A3(new_n203), .ZN(new_n345));
  OAI21_X1  g0145(.A(KEYINPUT12), .B1(new_n302), .B2(G68), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n297), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(new_n307), .B2(new_n207), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n300), .ZN(new_n349));
  XNOR2_X1  g0149(.A(KEYINPUT77), .B(KEYINPUT11), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n348), .A2(new_n300), .A3(new_n350), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n345), .A2(new_n346), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n343), .A2(new_n354), .ZN(new_n355));
  AND2_X1   g0155(.A1(KEYINPUT3), .A2(G33), .ZN(new_n356));
  NOR2_X1   g0156(.A1(KEYINPUT3), .A2(G33), .ZN(new_n357));
  OAI211_X1 g0157(.A(G232), .B(G1698), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  OAI211_X1 g0158(.A(G226), .B(new_n255), .C1(new_n356), .C2(new_n357), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G33), .A2(G97), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n265), .ZN(new_n362));
  INV_X1    g0162(.A(new_n254), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G238), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n270), .B1(new_n269), .B2(new_n265), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n275), .A2(KEYINPUT69), .A3(new_n278), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT13), .B1(new_n364), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(G238), .B1(new_n271), .B2(new_n279), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT13), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n254), .B1(new_n361), .B2(new_n265), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n369), .A2(G179), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G169), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n375), .B1(new_n369), .B2(new_n373), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT14), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n374), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  AOI211_X1 g0178(.A(KEYINPUT14), .B(new_n375), .C1(new_n369), .C2(new_n373), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n355), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT73), .B1(new_n302), .B2(new_n303), .ZN(new_n381));
  AOI211_X1 g0181(.A(new_n337), .B(new_n300), .C1(new_n286), .C2(new_n289), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n341), .A2(G77), .ZN(new_n383));
  NOR3_X1   g0183(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n290), .A2(KEYINPUT72), .A3(new_n207), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT72), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n302), .B2(G77), .ZN(new_n388));
  INV_X1    g0188(.A(new_n308), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n389), .A2(new_n297), .B1(G20), .B2(G77), .ZN(new_n390));
  XNOR2_X1  g0190(.A(KEYINPUT15), .B(G87), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n390), .B1(new_n307), .B2(new_n391), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n386), .A2(new_n388), .B1(new_n392), .B2(new_n300), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n260), .A2(G238), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n262), .A2(G232), .A3(new_n255), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n356), .A2(new_n357), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G107), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n394), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n254), .B1(new_n398), .B2(new_n265), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n211), .B1(new_n271), .B2(new_n279), .ZN(new_n400));
  INV_X1    g0200(.A(G190), .ZN(new_n401));
  AND3_X1   g0201(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(G200), .B1(new_n399), .B2(new_n400), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n385), .B(new_n393), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(G200), .ZN(new_n405));
  INV_X1    g0205(.A(new_n373), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n371), .B1(new_n370), .B2(new_n372), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n369), .A2(new_n401), .A3(new_n373), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n355), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n386), .A2(new_n388), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n392), .A2(new_n300), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AND3_X1   g0214(.A1(new_n399), .A2(new_n400), .A3(G179), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n375), .B1(new_n399), .B2(new_n400), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n414), .A2(new_n384), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n380), .A2(new_n404), .A3(new_n411), .A4(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT78), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n229), .A2(new_n257), .ZN(new_n420));
  INV_X1    g0220(.A(G159), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(G58), .A2(G68), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n204), .A2(new_n205), .A3(new_n423), .ZN(new_n424));
  AOI211_X1 g0224(.A(new_n419), .B(new_n422), .C1(new_n424), .C2(G20), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n258), .A2(new_n229), .A3(new_n259), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT7), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n396), .A2(KEYINPUT7), .A3(new_n229), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n203), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n424), .A2(G20), .ZN(new_n431));
  INV_X1    g0231(.A(new_n422), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI22_X1  g0233(.A1(new_n425), .A2(KEYINPUT16), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT7), .B1(new_n396), .B2(new_n229), .ZN(new_n435));
  NOR4_X1   g0235(.A1(new_n356), .A2(new_n357), .A3(new_n427), .A4(G20), .ZN(new_n436));
  OAI21_X1  g0236(.A(G68), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT16), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n422), .B1(new_n424), .B2(G20), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n437), .A2(new_n419), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n434), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n300), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n340), .A2(new_n308), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n302), .A2(new_n443), .A3(new_n303), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(new_n302), .B2(new_n389), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  OAI211_X1 g0246(.A(G223), .B(new_n255), .C1(new_n356), .C2(new_n357), .ZN(new_n447));
  OAI211_X1 g0247(.A(G226), .B(G1698), .C1(new_n356), .C2(new_n357), .ZN(new_n448));
  INV_X1    g0248(.A(G87), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n447), .B(new_n448), .C1(new_n257), .C2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n265), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n265), .B1(new_n272), .B2(new_n287), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n254), .B1(new_n452), .B2(G232), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n451), .A2(new_n453), .A3(new_n401), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n451), .A2(new_n453), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n454), .B1(new_n455), .B2(G200), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n442), .A2(new_n446), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT17), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n451), .A2(new_n453), .A3(new_n333), .ZN(new_n460));
  AOI21_X1  g0260(.A(G169), .B1(new_n451), .B2(new_n453), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n303), .B1(new_n434), .B2(new_n440), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(new_n463), .B2(new_n445), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT18), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n442), .A2(KEYINPUT17), .A3(new_n446), .A4(new_n456), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT18), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n462), .B(new_n467), .C1(new_n463), .C2(new_n445), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n459), .A2(new_n465), .A3(new_n466), .A4(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n418), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n331), .A2(new_n335), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT79), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT79), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n331), .A2(new_n473), .A3(new_n335), .A4(new_n470), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT6), .ZN(new_n477));
  INV_X1    g0277(.A(G97), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n477), .A2(new_n478), .A3(G107), .ZN(new_n479));
  XNOR2_X1  g0279(.A(G97), .B(G107), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n479), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  OAI22_X1  g0281(.A1(new_n481), .A2(new_n229), .B1(new_n207), .B2(new_n420), .ZN(new_n482));
  INV_X1    g0282(.A(G107), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n483), .B1(new_n428), .B2(new_n429), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n300), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n287), .A2(G33), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n302), .A2(G97), .A3(new_n303), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n290), .A2(new_n478), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n485), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT82), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n260), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n491));
  OAI211_X1 g0291(.A(G244), .B(new_n255), .C1(new_n356), .C2(new_n357), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT80), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT4), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n493), .B1(new_n492), .B2(new_n494), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n491), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT81), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n492), .B2(new_n494), .ZN(new_n499));
  INV_X1    g0299(.A(G244), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n500), .B1(new_n258), .B2(new_n259), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n501), .A2(KEYINPUT81), .A3(KEYINPUT4), .A4(new_n255), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n490), .B1(new_n497), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n492), .A2(new_n494), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT80), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n499), .A2(new_n502), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n508), .A2(KEYINPUT82), .A3(new_n509), .A4(new_n491), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n504), .A2(new_n265), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(G45), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n339), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g0313(.A(KEYINPUT5), .B(G41), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n513), .A2(G274), .A3(new_n278), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n287), .A2(G45), .ZN(new_n516));
  INV_X1    g0316(.A(new_n514), .ZN(new_n517));
  OAI211_X1 g0317(.A(G257), .B(new_n278), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  AND2_X1   g0318(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n511), .A2(G179), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n375), .B1(new_n511), .B2(new_n519), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n489), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT83), .B1(new_n511), .B2(new_n519), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n511), .A2(KEYINPUT83), .A3(new_n519), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n405), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n489), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n511), .A2(new_n519), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n527), .B1(new_n528), .B2(new_n401), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n522), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(G116), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n531), .B1(new_n287), .B2(G33), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n338), .A2(new_n342), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n257), .A2(G97), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G33), .A2(G283), .ZN(new_n535));
  AOI21_X1  g0335(.A(G20), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n229), .A2(new_n531), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n300), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT20), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(KEYINPUT20), .B(new_n300), .C1(new_n536), .C2(new_n537), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n290), .A2(new_n531), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(G264), .B(G1698), .C1(new_n356), .C2(new_n357), .ZN(new_n543));
  OAI211_X1 g0343(.A(G257), .B(new_n255), .C1(new_n356), .C2(new_n357), .ZN(new_n544));
  XNOR2_X1  g0344(.A(KEYINPUT85), .B(G303), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n543), .B(new_n544), .C1(new_n262), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n265), .ZN(new_n547));
  OAI211_X1 g0347(.A(G270), .B(new_n278), .C1(new_n516), .C2(new_n517), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(new_n515), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n549), .A2(KEYINPUT21), .A3(G169), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n547), .A2(G179), .A3(new_n515), .A4(new_n548), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n533), .A2(new_n542), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n549), .A2(new_n405), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n547), .A2(new_n401), .A3(new_n515), .A4(new_n548), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n555), .A2(new_n533), .A3(new_n542), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n549), .A2(G169), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(new_n533), .B2(new_n542), .ZN(new_n558));
  OAI21_X1  g0358(.A(KEYINPUT86), .B1(new_n558), .B2(KEYINPUT21), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT86), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT21), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n540), .A2(new_n541), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(G116), .B2(new_n302), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n381), .A2(new_n382), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n563), .B1(new_n564), .B2(new_n532), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n560), .B(new_n561), .C1(new_n565), .C2(new_n557), .ZN(new_n566));
  AOI211_X1 g0366(.A(new_n552), .B(new_n556), .C1(new_n559), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n290), .A2(new_n391), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n302), .A2(G87), .A3(new_n303), .A4(new_n486), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n262), .A2(new_n229), .A3(G68), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT19), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n229), .B1(new_n360), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(G87), .A2(G97), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n483), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n293), .A2(new_n292), .A3(G97), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n571), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT84), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT84), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n577), .A2(new_n580), .A3(new_n571), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n576), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n568), .B(new_n569), .C1(new_n582), .C2(new_n303), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n287), .A2(G45), .A3(new_n253), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n278), .B(new_n585), .C1(new_n513), .C2(G250), .ZN(new_n586));
  OAI211_X1 g0386(.A(G238), .B(new_n255), .C1(new_n356), .C2(new_n357), .ZN(new_n587));
  OAI211_X1 g0387(.A(G244), .B(G1698), .C1(new_n356), .C2(new_n357), .ZN(new_n588));
  NAND2_X1  g0388(.A1(G33), .A2(G116), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n265), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n405), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(G190), .B2(new_n592), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(G169), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n333), .B2(new_n592), .ZN(new_n596));
  INV_X1    g0396(.A(new_n391), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n302), .A2(new_n303), .A3(new_n597), .A4(new_n486), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n568), .B(new_n598), .C1(new_n582), .C2(new_n303), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n584), .A2(new_n594), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n229), .B(G87), .C1(new_n356), .C2(new_n357), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT87), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n262), .A2(KEYINPUT87), .A3(new_n229), .A4(G87), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(new_n604), .A3(KEYINPUT22), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT22), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n601), .A2(new_n602), .A3(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT23), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(G20), .B2(new_n483), .ZN(new_n609));
  NOR3_X1   g0409(.A1(new_n229), .A2(KEYINPUT23), .A3(G107), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n589), .A2(G20), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n605), .A2(new_n607), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT24), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n605), .A2(KEYINPUT24), .A3(new_n607), .A4(new_n612), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n300), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(KEYINPUT25), .B1(new_n302), .B2(G107), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n302), .A2(G107), .A3(new_n303), .A4(new_n486), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT25), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n286), .A2(new_n289), .A3(new_n620), .A4(new_n483), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n618), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n617), .A2(new_n623), .ZN(new_n624));
  OAI211_X1 g0424(.A(G250), .B(new_n255), .C1(new_n356), .C2(new_n357), .ZN(new_n625));
  OAI211_X1 g0425(.A(G257), .B(G1698), .C1(new_n356), .C2(new_n357), .ZN(new_n626));
  NAND2_X1  g0426(.A1(G33), .A2(G294), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n265), .ZN(new_n629));
  OAI211_X1 g0429(.A(G264), .B(new_n278), .C1(new_n516), .C2(new_n517), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(new_n515), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(G169), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n333), .B2(new_n631), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n624), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n631), .A2(new_n405), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n629), .A2(new_n515), .A3(new_n630), .A4(new_n401), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n617), .A2(new_n623), .A3(new_n637), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n600), .A2(new_n634), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n567), .A2(new_n639), .ZN(new_n640));
  NOR3_X1   g0440(.A1(new_n476), .A2(new_n530), .A3(new_n640), .ZN(G372));
  INV_X1    g0441(.A(new_n335), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT89), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n417), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n385), .A2(new_n393), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n415), .A2(new_n416), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(new_n646), .A3(KEYINPUT89), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n411), .A2(new_n644), .A3(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n648), .A2(new_n380), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n459), .A2(new_n466), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n465), .B(new_n468), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n642), .B1(new_n651), .B2(new_n331), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n600), .B(new_n489), .C1(new_n520), .C2(new_n521), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(KEYINPUT88), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n528), .A2(G169), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n511), .A2(G179), .A3(new_n519), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n658), .A2(KEYINPUT26), .A3(new_n489), .A4(new_n600), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(KEYINPUT88), .B1(new_n653), .B2(new_n654), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n596), .A2(new_n599), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n559), .A2(new_n566), .ZN(new_n664));
  INV_X1    g0464(.A(new_n552), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(new_n665), .A3(new_n634), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n600), .A2(new_n638), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n663), .B1(new_n669), .B2(new_n530), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n662), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n652), .B1(new_n476), .B2(new_n671), .ZN(G369));
  NAND2_X1  g0472(.A1(new_n664), .A2(new_n665), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n221), .A2(G20), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT27), .B1(new_n339), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT27), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n287), .A2(new_n677), .A3(new_n674), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n676), .A2(G213), .A3(new_n678), .A4(G343), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT90), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n565), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n673), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n552), .B1(new_n559), .B2(new_n566), .ZN(new_n683));
  INV_X1    g0483(.A(new_n556), .ZN(new_n684));
  INV_X1    g0484(.A(new_n681), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT91), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT91), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n682), .A2(new_n686), .A3(new_n689), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n624), .A2(new_n633), .A3(new_n680), .ZN(new_n691));
  INV_X1    g0491(.A(new_n680), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n624), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n638), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n691), .B1(new_n694), .B2(new_n634), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n688), .A2(G330), .A3(new_n690), .A4(new_n695), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n617), .A2(new_n623), .A3(new_n637), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n680), .B1(new_n617), .B2(new_n623), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n634), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n624), .A2(new_n633), .A3(new_n680), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n701), .A2(new_n683), .A3(new_n692), .ZN(new_n702));
  OAI21_X1  g0502(.A(KEYINPUT92), .B1(new_n702), .B2(new_n691), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n695), .A2(new_n673), .A3(new_n680), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT92), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(new_n705), .A3(new_n700), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n696), .A2(new_n707), .ZN(G399));
  INV_X1    g0508(.A(new_n225), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  INV_X1    g0510(.A(G1), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n573), .A2(new_n483), .A3(new_n531), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(KEYINPUT93), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT93), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n715), .B1(new_n710), .B2(new_n233), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n714), .B1(new_n713), .B2(new_n716), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT28), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n680), .B1(new_n662), .B2(new_n670), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT29), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n667), .B1(new_n683), .B2(new_n634), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n511), .A2(KEYINPUT83), .A3(new_n519), .ZN(new_n723));
  OAI21_X1  g0523(.A(G200), .B1(new_n723), .B2(new_n523), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n511), .A2(new_n519), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n489), .B1(new_n725), .B2(G190), .ZN(new_n726));
  AOI22_X1  g0526(.A1(new_n724), .A2(new_n726), .B1(new_n658), .B2(new_n489), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n722), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n653), .A2(new_n654), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT96), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n729), .A2(new_n659), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n653), .A2(KEYINPUT96), .A3(new_n654), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n728), .A2(new_n731), .A3(new_n663), .A4(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(KEYINPUT29), .A3(new_n680), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n721), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n549), .A2(new_n631), .A3(new_n333), .A4(new_n592), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(KEYINPUT95), .B1(new_n528), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT95), .ZN(new_n739));
  AOI211_X1 g0539(.A(new_n739), .B(new_n736), .C1(new_n511), .C2(new_n519), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n629), .A2(new_n630), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n551), .A2(new_n742), .A3(new_n592), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n511), .A2(new_n743), .A3(new_n519), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT30), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n511), .A2(new_n743), .A3(KEYINPUT30), .A4(new_n519), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n692), .B1(new_n741), .B2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT31), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n680), .A2(new_n750), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n725), .A2(new_n736), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n752), .B1(new_n748), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(KEYINPUT94), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT94), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n756), .B(new_n752), .C1(new_n748), .C2(new_n753), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n751), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n727), .A2(new_n567), .A3(new_n639), .A4(new_n680), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(G330), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n735), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n718), .B1(new_n763), .B2(G1), .ZN(G364));
  NAND2_X1  g0564(.A1(new_n688), .A2(new_n690), .ZN(new_n765));
  INV_X1    g0565(.A(G330), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n688), .A2(G330), .A3(new_n690), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n711), .B1(new_n674), .B2(G45), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OR3_X1    g0570(.A1(new_n710), .A2(KEYINPUT97), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(KEYINPUT97), .B1(new_n710), .B2(new_n770), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n767), .A2(new_n768), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n765), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n228), .B1(G20), .B2(new_n375), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n333), .A2(new_n405), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n229), .A2(G190), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n229), .A2(new_n401), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n784), .A2(new_n333), .A3(G200), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n262), .B1(new_n783), .B2(new_n203), .C1(new_n449), .C2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G179), .A2(G200), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n782), .A2(new_n787), .ZN(new_n788));
  OR3_X1    g0588(.A1(new_n788), .A2(KEYINPUT32), .A3(new_n421), .ZN(new_n789));
  OAI21_X1  g0589(.A(KEYINPUT32), .B1(new_n788), .B2(new_n421), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n787), .A2(G190), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n789), .B(new_n790), .C1(new_n478), .C2(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n782), .A2(new_n333), .A3(G200), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT99), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n786), .B(new_n794), .C1(G107), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n781), .A2(new_n784), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n333), .A2(G200), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n784), .A2(new_n799), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n798), .A2(new_n232), .B1(new_n800), .B2(new_n202), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n782), .A2(new_n799), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n801), .B1(G77), .B2(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT98), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n797), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G322), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n396), .B1(new_n800), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(G294), .B2(new_n792), .ZN(new_n809));
  INV_X1    g0609(.A(new_n798), .ZN(new_n810));
  INV_X1    g0610(.A(new_n788), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n810), .A2(G326), .B1(new_n811), .B2(G329), .ZN(new_n812));
  INV_X1    g0612(.A(new_n785), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n813), .A2(G303), .B1(new_n803), .B2(G311), .ZN(new_n814));
  AND3_X1   g0614(.A1(new_n809), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(KEYINPUT33), .B(G317), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n783), .B1(new_n817), .B2(KEYINPUT100), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(KEYINPUT100), .B2(new_n817), .ZN(new_n819));
  INV_X1    g0619(.A(G283), .ZN(new_n820));
  INV_X1    g0620(.A(new_n796), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n815), .B(new_n819), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n780), .B1(new_n806), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n777), .A2(new_n779), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n709), .A2(new_n262), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n247), .A2(G45), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n233), .A2(G45), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n709), .A2(new_n396), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n829), .A2(G355), .B1(new_n531), .B2(new_n709), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n773), .B(new_n823), .C1(new_n824), .C2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n778), .A2(new_n832), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n774), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(G396));
  INV_X1    g0635(.A(KEYINPUT102), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n647), .A2(new_n644), .A3(new_n645), .A4(new_n692), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n645), .A2(new_n692), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n838), .A2(new_n404), .A3(new_n417), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n836), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n837), .A2(new_n836), .A3(new_n839), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n843), .B(new_n680), .C1(new_n662), .C2(new_n670), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n722), .A2(new_n727), .B1(new_n599), .B2(new_n596), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT88), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n729), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n848), .A2(new_n655), .A3(new_n659), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n692), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n850), .A2(new_n843), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n761), .B1(new_n845), .B2(new_n851), .ZN(new_n852));
  OR2_X1    g0652(.A1(new_n852), .A2(KEYINPUT103), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(KEYINPUT103), .ZN(new_n854));
  OR3_X1    g0654(.A1(new_n845), .A2(new_n851), .A3(new_n761), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n853), .A2(new_n773), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n779), .A2(new_n775), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n773), .B1(new_n207), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n800), .ZN(new_n859));
  INV_X1    g0659(.A(new_n783), .ZN(new_n860));
  AOI22_X1  g0660(.A1(G143), .A2(new_n859), .B1(new_n860), .B2(G150), .ZN(new_n861));
  INV_X1    g0661(.A(G137), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n861), .B1(new_n862), .B2(new_n798), .C1(new_n421), .C2(new_n802), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT34), .ZN(new_n864));
  INV_X1    g0664(.A(G132), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n262), .B1(new_n788), .B2(new_n865), .C1(new_n785), .C2(new_n232), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(G58), .B2(new_n792), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n864), .B(new_n867), .C1(new_n203), .C2(new_n821), .ZN(new_n868));
  INV_X1    g0668(.A(G294), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n793), .A2(new_n478), .B1(new_n800), .B2(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT101), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n796), .A2(G87), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n813), .A2(G107), .B1(new_n810), .B2(G303), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n262), .B1(new_n811), .B2(G311), .ZN(new_n874));
  AOI22_X1  g0674(.A1(G283), .A2(new_n860), .B1(new_n803), .B2(G116), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n871), .A2(new_n872), .A3(new_n876), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n868), .A2(new_n877), .ZN(new_n878));
  OAI221_X1 g0678(.A(new_n858), .B1(new_n780), .B2(new_n878), .C1(new_n843), .C2(new_n776), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n856), .A2(new_n879), .ZN(G384));
  INV_X1    g0680(.A(KEYINPUT110), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n380), .A2(KEYINPUT106), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n410), .B1(new_n355), .B2(new_n692), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT106), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n884), .B(new_n355), .C1(new_n378), .C2(new_n379), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n882), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT107), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT107), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n882), .A2(new_n883), .A3(new_n888), .A4(new_n885), .ZN(new_n889));
  OR2_X1    g0689(.A1(new_n883), .A2(new_n380), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT109), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n749), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n746), .B(new_n747), .C1(new_n738), .C2(new_n740), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(KEYINPUT109), .A3(new_n692), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT31), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n894), .A2(new_n752), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n759), .A2(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n891), .B(new_n843), .C1(new_n896), .C2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT37), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n678), .A2(G213), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n901), .A2(new_n676), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT16), .B1(new_n430), .B2(new_n433), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n303), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n462), .A2(new_n902), .B1(new_n905), .B2(new_n445), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n900), .B1(new_n457), .B2(new_n906), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n457), .A2(new_n464), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT108), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n902), .B1(new_n463), .B2(new_n445), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n908), .A2(new_n909), .A3(new_n900), .A4(new_n910), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n457), .A2(new_n464), .A3(new_n910), .A4(new_n900), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(KEYINPUT108), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n907), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n905), .A2(new_n445), .ZN(new_n915));
  INV_X1    g0715(.A(new_n902), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n469), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT38), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n914), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n457), .A2(new_n464), .A3(new_n910), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT37), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n912), .A2(KEYINPUT108), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n912), .A2(KEYINPUT108), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n910), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n469), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT38), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT40), .B1(new_n921), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n881), .B1(new_n899), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT40), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n911), .A2(new_n913), .B1(KEYINPUT37), .B2(new_n922), .ZN(new_n933));
  INV_X1    g0733(.A(new_n928), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n920), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n912), .B(new_n909), .ZN(new_n936));
  OAI211_X1 g0736(.A(KEYINPUT38), .B(new_n918), .C1(new_n936), .C2(new_n907), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n932), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n894), .A2(KEYINPUT109), .A3(new_n692), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT109), .B1(new_n894), .B2(new_n692), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n750), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(new_n759), .A3(new_n897), .ZN(new_n942));
  AND3_X1   g0742(.A1(new_n837), .A2(new_n836), .A3(new_n839), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n943), .A2(new_n840), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n889), .A2(new_n890), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n944), .B1(new_n945), .B2(new_n887), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n938), .A2(new_n942), .A3(new_n946), .A4(KEYINPUT110), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n920), .B1(new_n914), .B2(new_n919), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n937), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n942), .A2(new_n946), .A3(new_n949), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n931), .A2(new_n947), .B1(new_n932), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n475), .A2(new_n942), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n951), .B(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(G330), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT39), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n948), .B2(new_n937), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n935), .A2(new_n955), .A3(new_n937), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n882), .A2(new_n885), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n960), .A2(new_n692), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n891), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n645), .A2(new_n646), .A3(new_n680), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT105), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n963), .B1(new_n844), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n949), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n465), .A2(new_n468), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n916), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n962), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n475), .A2(new_n721), .A3(new_n734), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n972), .A2(new_n652), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n971), .B(new_n973), .Z(new_n974));
  AOI22_X1  g0774(.A1(new_n954), .A2(new_n974), .B1(new_n339), .B2(new_n675), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n974), .B2(new_n954), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT35), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n481), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n978), .A2(G116), .A3(new_n230), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n979), .A2(KEYINPUT104), .B1(new_n977), .B2(new_n481), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n980), .B1(KEYINPUT104), .B2(new_n979), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT36), .Z(new_n982));
  NAND2_X1  g0782(.A1(G50), .A2(G77), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n424), .A2(new_n983), .B1(G50), .B2(new_n203), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n984), .A2(new_n221), .A3(new_n339), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n976), .A2(new_n982), .A3(new_n985), .ZN(G367));
  NAND2_X1  g0786(.A1(new_n692), .A2(new_n489), .ZN(new_n987));
  INV_X1    g0787(.A(new_n522), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n727), .A2(new_n987), .B1(new_n988), .B2(new_n692), .ZN(new_n989));
  INV_X1    g0789(.A(new_n600), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n692), .A2(new_n583), .ZN(new_n991));
  MUX2_X1   g0791(.A(new_n663), .B(new_n990), .S(new_n991), .Z(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n994));
  OR3_X1    g0794(.A1(new_n696), .A2(new_n989), .A3(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n994), .B1(new_n696), .B2(new_n989), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(KEYINPUT111), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT111), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n995), .A2(new_n999), .A3(new_n996), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n989), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n702), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1003), .A2(KEYINPUT42), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n634), .B1(new_n724), .B2(new_n726), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1005), .A2(new_n988), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n1003), .A2(KEYINPUT42), .B1(new_n680), .B2(new_n1006), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n1004), .A2(new_n1007), .B1(KEYINPUT43), .B2(new_n993), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1001), .B(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n710), .B(KEYINPUT41), .Z(new_n1010));
  INV_X1    g0810(.A(KEYINPUT45), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT112), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n707), .B2(new_n1002), .ZN(new_n1013));
  AOI211_X1 g0813(.A(KEYINPUT112), .B(new_n989), .C1(new_n703), .C2(new_n706), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1011), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NOR3_X1   g0815(.A1(new_n702), .A2(KEYINPUT92), .A3(new_n691), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n705), .B1(new_n704), .B2(new_n700), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1002), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(KEYINPUT112), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n707), .A2(new_n1012), .A3(new_n1002), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1019), .A2(KEYINPUT45), .A3(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n703), .A2(new_n706), .A3(new_n989), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT44), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1015), .A2(new_n1021), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n696), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1015), .A2(new_n1021), .A3(new_n1024), .A4(new_n696), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n695), .B1(new_n673), .B2(new_n680), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1029), .A2(new_n702), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n768), .B(new_n1030), .Z(new_n1031));
  NOR2_X1   g0831(.A1(new_n762), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1027), .A2(new_n1028), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1010), .B1(new_n1033), .B2(new_n763), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1009), .B1(new_n1034), .B2(new_n770), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT113), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1009), .B(KEYINPUT113), .C1(new_n1034), .C2(new_n770), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n824), .B1(new_n225), .B2(new_n391), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n825), .B2(new_n243), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n773), .A2(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G294), .A2(new_n860), .B1(new_n811), .B2(G317), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT114), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n785), .B2(new_n531), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1043), .B1(new_n478), .B2(new_n795), .C1(KEYINPUT46), .C2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(KEYINPUT46), .B2(new_n1045), .ZN(new_n1047));
  INV_X1    g0847(.A(G311), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n396), .B1(new_n798), .B2(new_n1048), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n800), .A2(new_n545), .B1(new_n802), .B2(new_n820), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(G107), .C2(new_n792), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n795), .A2(new_n207), .B1(new_n802), .B2(new_n232), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n396), .B(new_n1053), .C1(G137), .C2(new_n811), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G150), .A2(new_n859), .B1(new_n860), .B2(G159), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n813), .A2(G58), .B1(new_n810), .B2(G143), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n792), .A2(G68), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(KEYINPUT47), .B1(new_n1052), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1052), .A2(KEYINPUT47), .A3(new_n1058), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n779), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n777), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1042), .B1(new_n1059), .B2(new_n1061), .C1(new_n993), .C2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1039), .A2(new_n1063), .ZN(G387));
  INV_X1    g0864(.A(new_n1031), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n770), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n396), .B1(new_n795), .B2(new_n531), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n545), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n810), .A2(G322), .B1(new_n803), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(G317), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1069), .B1(new_n1048), .B2(new_n783), .C1(new_n1070), .C2(new_n800), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT48), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n813), .A2(G294), .B1(G283), .B2(new_n792), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT49), .Z(new_n1077));
  AOI211_X1 g0877(.A(new_n1067), .B(new_n1077), .C1(G326), .C2(new_n811), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(G50), .A2(new_n859), .B1(new_n811), .B2(G150), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n396), .B1(new_n860), .B2(new_n389), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n597), .A2(new_n792), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n813), .A2(G77), .B1(new_n803), .B2(G68), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n421), .B2(new_n798), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1082), .B(new_n1084), .C1(G97), .C2(new_n796), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n779), .B1(new_n1078), .B2(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n829), .A2(new_n712), .B1(new_n483), .B2(new_n709), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n240), .A2(G45), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n308), .A2(G50), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT115), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1090), .A2(KEYINPUT50), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(KEYINPUT50), .ZN(new_n1092));
  AOI211_X1 g0892(.A(G45), .B(new_n712), .C1(G68), .C2(G77), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n825), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1087), .B1(new_n1088), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n773), .B1(new_n1096), .B2(new_n824), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1086), .B(new_n1097), .C1(new_n695), .C2(new_n1062), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1032), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1099), .A2(KEYINPUT116), .A3(new_n710), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n763), .B2(new_n1065), .ZN(new_n1101));
  AOI21_X1  g0901(.A(KEYINPUT116), .B1(new_n1099), .B2(new_n710), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1066), .B(new_n1098), .C1(new_n1101), .C2(new_n1102), .ZN(G393));
  NAND2_X1  g0903(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n1099), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1105), .A2(new_n710), .A3(new_n1033), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1027), .A2(new_n770), .A3(new_n1028), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n773), .ZN(new_n1108));
  NOR3_X1   g0908(.A1(new_n250), .A2(new_n709), .A3(new_n262), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n824), .B1(new_n225), .B2(new_n478), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1108), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n785), .A2(new_n820), .B1(new_n788), .B2(new_n807), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT117), .Z(new_n1113));
  OAI22_X1  g0913(.A1(new_n798), .A2(new_n1070), .B1(new_n800), .B2(new_n1048), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT52), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n396), .B1(new_n802), .B2(new_n869), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n1068), .B2(new_n860), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1118), .B1(new_n531), .B2(new_n793), .C1(new_n821), .C2(new_n483), .ZN(new_n1119));
  INV_X1    g0919(.A(G150), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n798), .A2(new_n1120), .B1(new_n800), .B2(new_n421), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT51), .Z(new_n1122));
  OAI21_X1  g0922(.A(new_n262), .B1(new_n785), .B2(new_n203), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(G77), .B2(new_n792), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n803), .A2(new_n389), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(G50), .A2(new_n860), .B1(new_n811), .B2(G143), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n872), .A2(new_n1124), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n1116), .A2(new_n1119), .B1(new_n1122), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1111), .B1(new_n1128), .B2(new_n779), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n1002), .B2(new_n1062), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1106), .A2(new_n1107), .A3(new_n1130), .ZN(G390));
  AOI21_X1  g0931(.A(new_n773), .B1(new_n308), .B2(new_n857), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT118), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n785), .A2(new_n1120), .ZN(new_n1134));
  XOR2_X1   g0934(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n1135));
  OAI221_X1 g0935(.A(new_n262), .B1(new_n865), .B2(new_n800), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n795), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n810), .A2(G128), .B1(new_n1137), .B2(G50), .ZN(new_n1138));
  INV_X1    g0938(.A(G125), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1138), .B1(new_n1139), .B2(new_n788), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1136), .B(new_n1140), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT54), .B(G143), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n783), .A2(new_n862), .B1(new_n802), .B2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G159), .B2(new_n792), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT119), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n396), .B1(new_n785), .B2(new_n449), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n798), .A2(new_n820), .B1(new_n800), .B2(new_n531), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1146), .B(new_n1147), .C1(G77), .C2(new_n792), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(G97), .A2(new_n803), .B1(new_n811), .B2(G294), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n483), .B2(new_n783), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(G68), .B2(new_n796), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1141), .A2(new_n1145), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT121), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n779), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1133), .B1(new_n1154), .B2(new_n1156), .C1(new_n959), .C2(new_n776), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n921), .A2(new_n929), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n956), .B1(new_n1158), .B2(new_n955), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n967), .B2(new_n961), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n733), .A2(new_n680), .A3(new_n843), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n966), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n891), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n961), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n921), .B2(new_n929), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n946), .B(G330), .C1(new_n760), .C2(new_n758), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1160), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1165), .B1(new_n1162), .B2(new_n891), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n965), .B1(new_n850), .B2(new_n843), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1164), .B1(new_n1171), .B2(new_n963), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1170), .B1(new_n1159), .B2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n944), .A2(new_n766), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n942), .A2(new_n891), .A3(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1169), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1157), .B1(new_n1176), .B2(new_n769), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT122), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(KEYINPUT76), .B1(new_n327), .B2(new_n319), .ZN(new_n1180));
  AND4_X1   g0980(.A1(KEYINPUT76), .A2(new_n315), .A3(new_n319), .A4(new_n321), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n282), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(KEYINPUT10), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n642), .B1(new_n1183), .B2(new_n323), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n473), .B1(new_n1184), .B2(new_n470), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n474), .ZN(new_n1186));
  OAI211_X1 g0986(.A(G330), .B(new_n942), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n942), .A2(new_n1174), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n963), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1162), .ZN(new_n1190));
  AND3_X1   g0990(.A1(new_n1189), .A2(new_n1168), .A3(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n963), .B1(new_n761), .B2(new_n944), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1171), .B1(new_n1192), .B2(new_n1175), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n973), .B(new_n1187), .C1(new_n1191), .C2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1176), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n972), .A2(new_n1187), .A3(new_n652), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1192), .A2(new_n1175), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n844), .A2(new_n966), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1189), .A2(new_n1190), .A3(new_n1168), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1196), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1175), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1198), .A2(new_n891), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n959), .B1(new_n1203), .B2(new_n1164), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1202), .B1(new_n1204), .B2(new_n1170), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1201), .A2(new_n1205), .A3(new_n1169), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1195), .A2(new_n710), .A3(new_n1206), .ZN(new_n1207));
  OAI211_X1 g1007(.A(KEYINPUT122), .B(new_n1157), .C1(new_n1176), .C2(new_n769), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1179), .A2(new_n1207), .A3(new_n1208), .ZN(G378));
  NAND2_X1  g1009(.A1(new_n931), .A2(new_n947), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n950), .A2(new_n932), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1210), .A2(G330), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n326), .A2(new_n902), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1184), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n331), .A2(new_n335), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1213), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1214), .A2(new_n1217), .ZN(new_n1218));
  XOR2_X1   g1018(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1219), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1214), .A2(new_n1217), .A3(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1212), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n971), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n951), .A2(G330), .A3(new_n1223), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1226), .B1(new_n1225), .B2(new_n1227), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n770), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1224), .A2(new_n775), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n857), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1108), .B1(G50), .B2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n232), .B1(G33), .B2(G41), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(new_n396), .B2(new_n277), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n813), .A2(G77), .B1(new_n860), .B2(G97), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n202), .B2(new_n795), .C1(new_n531), .C2(new_n798), .ZN(new_n1237));
  AOI211_X1 g1037(.A(G41), .B(new_n262), .C1(new_n859), .C2(G107), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1238), .B1(new_n820), .B2(new_n788), .C1(new_n391), .C2(new_n802), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1237), .B(new_n1239), .C1(G68), .C2(new_n792), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1235), .B1(new_n1240), .B2(KEYINPUT58), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n785), .A2(new_n1142), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1242), .A2(KEYINPUT123), .B1(G150), .B2(new_n792), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(KEYINPUT123), .B2(new_n1242), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n798), .A2(new_n1139), .B1(new_n802), .B2(new_n862), .ZN(new_n1245));
  INV_X1    g1045(.A(G128), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n1246), .A2(new_n800), .B1(new_n783), .B2(new_n865), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(new_n1244), .A2(new_n1245), .A3(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1249), .A2(KEYINPUT59), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n257), .B(new_n277), .C1(new_n795), .C2(new_n421), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(G124), .B2(new_n811), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT59), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1252), .B1(new_n1248), .B2(new_n1253), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n1241), .B1(KEYINPUT58), .B2(new_n1240), .C1(new_n1250), .C2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1233), .B1(new_n1255), .B2(new_n779), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1231), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1230), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n710), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT124), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1196), .A2(new_n1260), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n972), .A2(new_n1187), .A3(KEYINPUT124), .A4(new_n652), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n1176), .B2(new_n1194), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT57), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1259), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1266), .B1(new_n1206), .B2(new_n1263), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n1229), .B2(KEYINPUT125), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT125), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n1271), .B(new_n1226), .C1(new_n1225), .C2(new_n1227), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1268), .B1(new_n1270), .B2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1258), .B1(new_n1267), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(G375));
  XNOR2_X1  g1075(.A(new_n769), .B(KEYINPUT126), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n963), .A2(new_n775), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1108), .B1(G68), .B2(new_n1232), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(G116), .A2(new_n860), .B1(new_n811), .B2(G303), .ZN(new_n1280));
  OAI221_X1 g1080(.A(new_n1280), .B1(new_n869), .B2(new_n798), .C1(new_n821), .C2(new_n207), .ZN(new_n1281));
  AOI22_X1  g1081(.A1(new_n813), .A2(G97), .B1(new_n803), .B2(G107), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n262), .B1(new_n859), .B2(G283), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1282), .A2(new_n1081), .A3(new_n1283), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(G150), .A2(new_n803), .B1(new_n811), .B2(G128), .ZN(new_n1285));
  OAI221_X1 g1085(.A(new_n1285), .B1(new_n421), .B2(new_n785), .C1(new_n783), .C2(new_n1142), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(G132), .A2(new_n810), .B1(new_n859), .B2(G137), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n396), .B1(new_n1137), .B2(G58), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1287), .B(new_n1288), .C1(new_n232), .C2(new_n793), .ZN(new_n1289));
  OAI22_X1  g1089(.A1(new_n1281), .A2(new_n1284), .B1(new_n1286), .B2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1279), .B1(new_n779), .B2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1277), .B1(new_n1278), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1010), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1199), .A2(new_n1196), .A3(new_n1200), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1194), .A2(new_n1293), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1292), .A2(new_n1295), .ZN(G381));
  INV_X1    g1096(.A(new_n1063), .ZN(new_n1297));
  AOI211_X1 g1097(.A(new_n1297), .B(G390), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1298));
  INV_X1    g1098(.A(G378), .ZN(new_n1299));
  NOR4_X1   g1099(.A1(G393), .A2(G381), .A3(G384), .A4(G396), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1298), .A2(new_n1299), .A3(new_n1274), .A4(new_n1300), .ZN(G407));
  INV_X1    g1101(.A(G343), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(G213), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1274), .A2(new_n1299), .A3(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(G407), .A2(G213), .A3(new_n1305), .ZN(G409));
  NAND2_X1  g1106(.A1(G387), .A2(G390), .ZN(new_n1307));
  INV_X1    g1107(.A(G390), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1039), .A2(new_n1063), .A3(new_n1308), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(G393), .B(new_n834), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1307), .A2(new_n1309), .A3(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1308), .B1(new_n1039), .B2(new_n1063), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1310), .B1(new_n1313), .B2(new_n1298), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1312), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1304), .A2(G2897), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  AND2_X1   g1117(.A1(new_n1294), .A2(KEYINPUT60), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1294), .A2(KEYINPUT60), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n710), .B(new_n1194), .C1(new_n1318), .C2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1320), .A2(G384), .A3(new_n1292), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(G384), .B1(new_n1320), .B2(new_n1292), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1317), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1323), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1325), .A2(new_n1321), .A3(new_n1316), .ZN(new_n1326));
  AND2_X1   g1126(.A1(new_n1324), .A2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1257), .ZN(new_n1328));
  AND4_X1   g1128(.A1(G330), .A2(new_n1210), .A3(new_n1211), .A4(new_n1223), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1223), .B1(new_n951), .B2(G330), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n971), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  AOI22_X1  g1131(.A1(new_n1331), .A2(new_n1269), .B1(new_n1206), .B2(new_n1263), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1328), .B1(new_n1332), .B2(new_n1293), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1276), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1334), .B1(new_n1270), .B2(new_n1272), .ZN(new_n1335));
  AOI21_X1  g1135(.A(G378), .B1(new_n1333), .B2(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1336), .B1(G378), .B2(new_n1274), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1327), .B1(new_n1337), .B2(new_n1304), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1258), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1264), .A2(KEYINPUT57), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1228), .B1(new_n1271), .B2(new_n1331), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1272), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1340), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n710), .B1(new_n1332), .B2(KEYINPUT57), .ZN(new_n1344));
  OAI211_X1 g1144(.A(G378), .B(new_n1339), .C1(new_n1343), .C2(new_n1344), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1276), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1257), .B1(new_n1265), .B2(new_n1010), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1299), .B1(new_n1346), .B2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1345), .A2(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT62), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1351));
  NAND4_X1  g1151(.A1(new_n1349), .A2(new_n1350), .A3(new_n1303), .A4(new_n1351), .ZN(new_n1352));
  XNOR2_X1  g1152(.A(KEYINPUT127), .B(KEYINPUT61), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1338), .A2(new_n1352), .A3(new_n1353), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1304), .B1(new_n1345), .B2(new_n1348), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1350), .B1(new_n1355), .B2(new_n1351), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1315), .B1(new_n1354), .B2(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1355), .A2(new_n1351), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1324), .A2(new_n1326), .ZN(new_n1359));
  AOI21_X1  g1159(.A(new_n1359), .B1(new_n1349), .B2(new_n1303), .ZN(new_n1360));
  INV_X1    g1160(.A(KEYINPUT63), .ZN(new_n1361));
  OAI21_X1  g1161(.A(new_n1358), .B1(new_n1360), .B2(new_n1361), .ZN(new_n1362));
  INV_X1    g1162(.A(KEYINPUT61), .ZN(new_n1363));
  AND3_X1   g1163(.A1(new_n1312), .A2(new_n1314), .A3(new_n1363), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1355), .A2(KEYINPUT63), .A3(new_n1351), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1362), .A2(new_n1364), .A3(new_n1365), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1357), .A2(new_n1366), .ZN(G405));
  XNOR2_X1  g1167(.A(new_n1274), .B(G378), .ZN(new_n1368));
  INV_X1    g1168(.A(new_n1368), .ZN(new_n1369));
  AND3_X1   g1169(.A1(new_n1312), .A2(new_n1314), .A3(new_n1351), .ZN(new_n1370));
  AOI21_X1  g1170(.A(new_n1351), .B1(new_n1312), .B2(new_n1314), .ZN(new_n1371));
  OAI21_X1  g1171(.A(new_n1369), .B1(new_n1370), .B2(new_n1371), .ZN(new_n1372));
  AOI21_X1  g1172(.A(new_n1311), .B1(new_n1307), .B2(new_n1309), .ZN(new_n1373));
  NOR3_X1   g1173(.A1(new_n1313), .A2(new_n1298), .A3(new_n1310), .ZN(new_n1374));
  OAI22_X1  g1174(.A1(new_n1373), .A2(new_n1374), .B1(new_n1323), .B2(new_n1322), .ZN(new_n1375));
  NAND3_X1  g1175(.A1(new_n1312), .A2(new_n1314), .A3(new_n1351), .ZN(new_n1376));
  NAND3_X1  g1176(.A1(new_n1375), .A2(new_n1368), .A3(new_n1376), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1372), .A2(new_n1377), .ZN(G402));
endmodule


