//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n440, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n578, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n624, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1233,
    new_n1234;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G120), .Z(new_n440));
  INV_X1    g015(.A(new_n440), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(new_n440), .A2(G57), .A3(G69), .A4(G108), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT66), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n462), .A2(new_n464), .A3(G137), .ZN(new_n465));
  NAND2_X1  g040(.A1(G101), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n462), .A2(new_n464), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n467), .B1(G2105), .B2(new_n471), .ZN(G160));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(KEYINPUT67), .A3(G124), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n477));
  INV_X1    g052(.A(G124), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n477), .B1(new_n474), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n469), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n483), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n476), .A2(new_n479), .A3(new_n481), .A4(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  NAND4_X1  g061(.A1(new_n462), .A2(new_n464), .A3(G138), .A4(new_n483), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n473), .A2(KEYINPUT4), .A3(G138), .A4(new_n483), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(new_n483), .B2(G114), .ZN(new_n492));
  INV_X1    g067(.A(G102), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(new_n483), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n462), .A2(new_n464), .A3(G126), .A4(G2105), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n473), .A2(KEYINPUT68), .A3(G126), .A4(G2105), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n494), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n491), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  NAND2_X1  g076(.A1(G75), .A2(G543), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT69), .A2(KEYINPUT5), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT69), .A2(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g079(.A(G543), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT70), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n509));
  OAI211_X1 g084(.A(new_n509), .B(G543), .C1(new_n503), .C2(new_n504), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n506), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G62), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n502), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G50), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n506), .A2(new_n508), .A3(new_n510), .A4(new_n515), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n514), .A2(new_n521), .ZN(G166));
  INV_X1    g097(.A(new_n519), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G89), .ZN(new_n524));
  AND3_X1   g099(.A1(new_n506), .A2(new_n508), .A3(new_n510), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n517), .A2(G51), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT71), .B(KEYINPUT7), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n528), .B(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n524), .A2(new_n526), .A3(new_n527), .A4(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  NAND2_X1  g108(.A1(new_n517), .A2(G52), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n519), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(KEYINPUT72), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT72), .ZN(new_n538));
  OAI211_X1 g113(.A(new_n538), .B(new_n534), .C1(new_n519), .C2(new_n535), .ZN(new_n539));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G64), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n511), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n537), .A2(new_n539), .B1(G651), .B2(new_n542), .ZN(G171));
  NAND4_X1  g118(.A1(new_n506), .A2(G56), .A3(new_n508), .A4(new_n510), .ZN(new_n544));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g121(.A(KEYINPUT73), .B1(new_n546), .B2(G651), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT73), .ZN(new_n548));
  INV_X1    g123(.A(G651), .ZN(new_n549));
  AOI211_X1 g124(.A(new_n548), .B(new_n549), .C1(new_n544), .C2(new_n545), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n517), .A2(G43), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n519), .B2(new_n552), .ZN(new_n553));
  NOR3_X1   g128(.A1(new_n547), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(G188));
  NAND4_X1  g135(.A1(new_n506), .A2(G65), .A3(new_n508), .A4(new_n510), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT75), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT76), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n561), .A2(KEYINPUT76), .A3(new_n563), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n566), .A2(G651), .A3(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT74), .ZN(new_n569));
  AND2_X1   g144(.A1(new_n519), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n519), .A2(new_n569), .ZN(new_n571));
  OAI21_X1  g146(.A(G91), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n517), .A2(G53), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT9), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n568), .A2(new_n572), .A3(new_n574), .ZN(G299));
  INV_X1    g150(.A(G171), .ZN(G301));
  INV_X1    g151(.A(G166), .ZN(G303));
  NAND3_X1  g152(.A1(new_n525), .A2(KEYINPUT74), .A3(new_n515), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n519), .A2(new_n569), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G87), .B1(G49), .B2(new_n517), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G288));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n511), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n586), .A2(G651), .B1(G48), .B2(new_n517), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n570), .A2(new_n571), .ZN(new_n588));
  INV_X1    g163(.A(G86), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(KEYINPUT77), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT77), .ZN(new_n592));
  OAI211_X1 g167(.A(new_n587), .B(new_n592), .C1(new_n588), .C2(new_n589), .ZN(new_n593));
  AND2_X1   g168(.A1(new_n591), .A2(new_n593), .ZN(G305));
  NAND2_X1  g169(.A1(new_n525), .A2(G60), .ZN(new_n595));
  NAND2_X1  g170(.A1(G72), .A2(G543), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n549), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  XNOR2_X1  g173(.A(KEYINPUT78), .B(G47), .ZN(new_n599));
  OAI22_X1  g174(.A1(new_n519), .A2(new_n598), .B1(new_n516), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n604), .B1(new_n580), .B2(G92), .ZN(new_n605));
  INV_X1    g180(.A(G92), .ZN(new_n606));
  AOI211_X1 g181(.A(KEYINPUT10), .B(new_n606), .C1(new_n578), .C2(new_n579), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(G79), .A2(G543), .ZN(new_n609));
  XNOR2_X1  g184(.A(KEYINPUT79), .B(G66), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n511), .B2(new_n610), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n611), .A2(G651), .B1(G54), .B2(new_n517), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n608), .A2(KEYINPUT80), .A3(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(G92), .B1(new_n570), .B2(new_n571), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(KEYINPUT10), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n580), .A2(new_n604), .A3(G92), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n615), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT80), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n613), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n603), .B1(new_n620), .B2(G868), .ZN(G284));
  OAI21_X1  g196(.A(new_n603), .B1(new_n620), .B2(G868), .ZN(G321));
  NAND2_X1  g197(.A1(G286), .A2(G868), .ZN(new_n623));
  AND3_X1   g198(.A1(new_n568), .A2(new_n572), .A3(new_n574), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(G868), .ZN(G297));
  OAI21_X1  g200(.A(new_n623), .B1(new_n624), .B2(G868), .ZN(G280));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n620), .B1(new_n627), .B2(G860), .ZN(G148));
  NAND2_X1  g203(.A1(new_n546), .A2(G651), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(new_n548), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n523), .A2(G81), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n546), .A2(KEYINPUT73), .A3(G651), .ZN(new_n632));
  NAND4_X1  g207(.A1(new_n630), .A2(new_n631), .A3(new_n551), .A4(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(G868), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n620), .A2(new_n627), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n635), .B1(new_n637), .B2(new_n634), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g214(.A1(new_n480), .A2(G2104), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT13), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2100), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n475), .A2(KEYINPUT81), .A3(G123), .ZN(new_n644));
  INV_X1    g219(.A(KEYINPUT81), .ZN(new_n645));
  INV_X1    g220(.A(G123), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n645), .B1(new_n474), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n480), .A2(G135), .ZN(new_n648));
  OR2_X1    g223(.A1(G99), .A2(G2105), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n649), .B(G2104), .C1(G111), .C2(new_n483), .ZN(new_n650));
  NAND4_X1  g225(.A1(new_n644), .A2(new_n647), .A3(new_n648), .A4(new_n650), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n651), .A2(G2096), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(G2096), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n643), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT82), .ZN(G156));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT83), .B(G2438), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2427), .B(G2430), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(KEYINPUT14), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2451), .B(G2454), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT16), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2443), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n661), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(KEYINPUT84), .B(KEYINPUT85), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G1341), .B(G1348), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2446), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n667), .A2(new_n670), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n671), .A2(G14), .A3(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G401));
  XOR2_X1   g249(.A(G2072), .B(G2078), .Z(new_n675));
  XOR2_X1   g250(.A(G2067), .B(G2678), .Z(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT86), .B(KEYINPUT18), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n675), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2096), .B(G2100), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n677), .A2(new_n678), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n685), .A2(new_n679), .A3(KEYINPUT17), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n686), .A2(new_n680), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n684), .B(new_n687), .Z(G227));
  XNOR2_X1  g263(.A(G1971), .B(G1976), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  XOR2_X1   g265(.A(G1956), .B(G2474), .Z(new_n691));
  XOR2_X1   g266(.A(G1961), .B(G1966), .Z(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n692), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT20), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n694), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n690), .A2(new_n693), .A3(new_n695), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n698), .B(new_n699), .C1(new_n697), .C2(new_n696), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT21), .B(G1986), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(G1991), .B(G1996), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT22), .B(G1981), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n704), .B(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(G229));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G23), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G288), .B2(G16), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT33), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n714), .A2(G1976), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G1976), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n712), .A2(new_n713), .ZN(new_n718));
  AOI211_X1 g293(.A(KEYINPUT33), .B(new_n711), .C1(G288), .C2(G16), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n709), .A2(G22), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G166), .B2(new_n709), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n722), .A2(G1971), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(G1971), .ZN(new_n724));
  NAND4_X1  g299(.A1(new_n716), .A2(new_n720), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G1981), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n591), .A2(new_n593), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G16), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT32), .ZN(new_n730));
  NOR2_X1   g305(.A1(G6), .A2(G16), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n709), .B1(new_n591), .B2(new_n593), .ZN(new_n734));
  OAI21_X1  g309(.A(KEYINPUT32), .B1(new_n734), .B2(new_n731), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n727), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n733), .A2(new_n727), .A3(new_n735), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n726), .A2(new_n739), .A3(KEYINPUT34), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT34), .ZN(new_n741));
  AND3_X1   g316(.A1(new_n733), .A2(new_n727), .A3(new_n735), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n742), .A2(new_n736), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n741), .B1(new_n743), .B2(new_n725), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT36), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n746), .A2(KEYINPUT91), .ZN(new_n747));
  INV_X1    g322(.A(G24), .ZN(new_n748));
  OAI21_X1  g323(.A(KEYINPUT90), .B1(new_n748), .B2(G16), .ZN(new_n749));
  OR3_X1    g324(.A1(new_n748), .A2(KEYINPUT90), .A3(G16), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n749), .B(new_n750), .C1(new_n601), .C2(new_n709), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G1986), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  OR3_X1    g328(.A1(KEYINPUT87), .A2(G95), .A3(G2105), .ZN(new_n754));
  INV_X1    g329(.A(G107), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n461), .B1(new_n755), .B2(G2105), .ZN(new_n756));
  OAI21_X1  g331(.A(KEYINPUT87), .B1(G95), .B2(G2105), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n754), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT88), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n475), .A2(G119), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n480), .A2(G131), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n759), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  MUX2_X1   g337(.A(G25), .B(new_n762), .S(G29), .Z(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT89), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT35), .B(G1991), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n745), .A2(new_n747), .A3(new_n753), .A4(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n709), .A2(KEYINPUT23), .A3(G20), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT23), .ZN(new_n769));
  INV_X1    g344(.A(G20), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n770), .B2(G16), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n768), .B(new_n771), .C1(new_n624), .C2(new_n709), .ZN(new_n772));
  INV_X1    g347(.A(G1956), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G29), .A2(G33), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT94), .Z(new_n776));
  NAND3_X1  g351(.A1(new_n483), .A2(G103), .A3(G2104), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT25), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n480), .A2(G139), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n778), .B(new_n779), .C1(new_n483), .C2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(G29), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n776), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(KEYINPUT95), .A2(G2072), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(KEYINPUT95), .A2(G2072), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT24), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n788), .A2(G34), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n788), .A2(G34), .ZN(new_n791));
  AOI21_X1  g366(.A(G29), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n467), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n471), .A2(G2105), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n792), .B1(new_n795), .B2(G29), .ZN(new_n796));
  INV_X1    g371(.A(G2084), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT96), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT26), .ZN(new_n801));
  NAND2_X1  g376(.A1(G105), .A2(G2104), .ZN(new_n802));
  INV_X1    g377(.A(G141), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n469), .B2(new_n803), .ZN(new_n804));
  AOI22_X1  g379(.A1(G129), .A2(new_n475), .B1(new_n804), .B2(new_n483), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n806), .A2(new_n782), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(KEYINPUT97), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT27), .B(G1996), .Z(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT97), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G29), .B2(G32), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n808), .B(new_n810), .C1(new_n807), .C2(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n787), .A2(new_n798), .A3(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT98), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n709), .A2(G5), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G171), .B2(new_n709), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT101), .ZN(new_n818));
  INV_X1    g393(.A(G1961), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n796), .A2(new_n797), .ZN(new_n821));
  NOR2_X1   g396(.A1(G164), .A2(new_n782), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G27), .B2(new_n782), .ZN(new_n823));
  INV_X1    g398(.A(G2078), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n815), .A2(new_n820), .A3(new_n821), .A4(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n818), .A2(new_n819), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n709), .A2(G21), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G168), .B2(new_n709), .ZN(new_n829));
  INV_X1    g404(.A(G1966), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT31), .B(G11), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT99), .B(G28), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT30), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(new_n782), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n832), .B(new_n835), .C1(new_n651), .C2(new_n782), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT100), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n823), .A2(new_n824), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n831), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n826), .A2(new_n827), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n709), .A2(G19), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(new_n554), .B2(new_n709), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(G1341), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n475), .A2(G128), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n480), .A2(G140), .ZN(new_n845));
  NOR2_X1   g420(.A1(G104), .A2(G2105), .ZN(new_n846));
  OAI21_X1  g421(.A(G2104), .B1(new_n483), .B2(G116), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n844), .B(new_n845), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G29), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n782), .A2(G26), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT92), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT28), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(G2067), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n709), .B1(new_n613), .B2(new_n619), .ZN(new_n856));
  NOR2_X1   g431(.A1(G4), .A2(G16), .ZN(new_n857));
  OAI21_X1  g432(.A(G1348), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NOR3_X1   g434(.A1(new_n856), .A2(G1348), .A3(new_n857), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n843), .B(new_n855), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT93), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n860), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(new_n858), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n865), .A2(KEYINPUT93), .A3(new_n843), .A4(new_n855), .ZN(new_n866));
  AND4_X1   g441(.A1(new_n774), .A2(new_n840), .A3(new_n863), .A4(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n808), .B1(new_n807), .B2(new_n812), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(new_n809), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n767), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n782), .A2(G35), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(G162), .B2(new_n782), .ZN(new_n872));
  XOR2_X1   g447(.A(KEYINPUT29), .B(G2090), .Z(new_n873));
  XOR2_X1   g448(.A(new_n872), .B(new_n873), .Z(new_n874));
  INV_X1    g449(.A(new_n747), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n746), .A2(KEYINPUT91), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n752), .B1(new_n740), .B2(new_n744), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n877), .B1(new_n878), .B2(new_n766), .ZN(new_n879));
  NOR3_X1   g454(.A1(new_n870), .A2(new_n874), .A3(new_n879), .ZN(G311));
  AND2_X1   g455(.A1(new_n767), .A2(new_n867), .ZN(new_n881));
  INV_X1    g456(.A(new_n879), .ZN(new_n882));
  INV_X1    g457(.A(new_n874), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n881), .A2(new_n882), .A3(new_n883), .A4(new_n869), .ZN(G150));
  NAND2_X1  g459(.A1(new_n620), .A2(G559), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT39), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n506), .A2(G67), .A3(new_n508), .A4(new_n510), .ZN(new_n887));
  NAND2_X1  g462(.A1(G80), .A2(G543), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(KEYINPUT102), .B1(new_n889), .B2(G651), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT102), .ZN(new_n891));
  AOI211_X1 g466(.A(new_n891), .B(new_n549), .C1(new_n887), .C2(new_n888), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n517), .A2(G55), .ZN(new_n893));
  INV_X1    g468(.A(G93), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n893), .B1(new_n519), .B2(new_n894), .ZN(new_n895));
  NOR3_X1   g470(.A1(new_n890), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n633), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n889), .A2(G651), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n891), .ZN(new_n899));
  INV_X1    g474(.A(new_n895), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n889), .A2(KEYINPUT102), .A3(G651), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n554), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n897), .A2(new_n903), .ZN(new_n904));
  XOR2_X1   g479(.A(new_n904), .B(KEYINPUT38), .Z(new_n905));
  XNOR2_X1  g480(.A(new_n886), .B(new_n905), .ZN(new_n906));
  XOR2_X1   g481(.A(KEYINPUT103), .B(G860), .Z(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT104), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n896), .A2(new_n908), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT37), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(G145));
  XNOR2_X1  g488(.A(new_n762), .B(new_n641), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(new_n781), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n651), .B(G160), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(G162), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n489), .A2(new_n490), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n919), .B1(new_n489), .B2(new_n490), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n499), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n918), .A2(new_n923), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n918), .A2(new_n923), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n916), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n916), .B1(new_n925), .B2(new_n924), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n475), .A2(G130), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n480), .A2(G142), .ZN(new_n930));
  NOR2_X1   g505(.A1(G106), .A2(G2105), .ZN(new_n931));
  OAI21_X1  g506(.A(G2104), .B1(new_n483), .B2(G118), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n929), .B(new_n930), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n806), .B(new_n933), .ZN(new_n934));
  XOR2_X1   g509(.A(new_n934), .B(new_n848), .Z(new_n935));
  NAND2_X1  g510(.A1(new_n928), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G37), .ZN(new_n937));
  INV_X1    g512(.A(new_n935), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(new_n926), .B2(new_n927), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n940), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n608), .A2(new_n624), .A3(new_n942), .A4(new_n612), .ZN(new_n943));
  NAND2_X1  g518(.A1(G299), .A2(KEYINPUT107), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n568), .A2(new_n572), .A3(new_n942), .A4(new_n574), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(new_n617), .A3(new_n945), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n943), .A2(new_n946), .A3(KEYINPUT41), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT41), .B1(new_n943), .B2(new_n946), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n904), .B(KEYINPUT106), .ZN(new_n950));
  OR2_X1    g525(.A1(new_n950), .A2(new_n636), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n636), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT42), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n943), .A2(new_n946), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n951), .A2(new_n952), .A3(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n954), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(G303), .B1(new_n581), .B2(new_n582), .ZN(new_n959));
  NOR2_X1   g534(.A1(G288), .A2(G166), .ZN(new_n960));
  OAI21_X1  g535(.A(G305), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n581), .A2(new_n582), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(G303), .ZN(new_n963));
  NAND2_X1  g538(.A1(G288), .A2(G166), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(new_n728), .A3(new_n964), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n961), .A2(new_n965), .A3(new_n601), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n601), .B1(new_n961), .B2(new_n965), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n951), .A2(new_n952), .A3(new_n956), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT42), .B1(new_n970), .B2(new_n953), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n958), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n969), .B1(new_n958), .B2(new_n971), .ZN(new_n973));
  OAI21_X1  g548(.A(G868), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n902), .A2(new_n634), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(G295));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n975), .ZN(G331));
  INV_X1    g552(.A(KEYINPUT43), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT108), .ZN(new_n979));
  NOR2_X1   g554(.A1(G171), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n542), .A2(G651), .ZN(new_n982));
  XNOR2_X1  g557(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n509), .B1(new_n983), .B2(G543), .ZN(new_n984));
  INV_X1    g559(.A(new_n510), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n986), .A2(G90), .A3(new_n508), .A4(new_n515), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n538), .B1(new_n987), .B2(new_n534), .ZN(new_n988));
  INV_X1    g563(.A(new_n539), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n979), .B(new_n982), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(G168), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n991), .A2(new_n903), .A3(new_n897), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n991), .B1(new_n903), .B2(new_n897), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n981), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n943), .A2(new_n946), .A3(KEYINPUT41), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT41), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n956), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(G286), .B1(G171), .B2(new_n979), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n904), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n991), .A2(new_n897), .A3(new_n903), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n999), .A2(new_n980), .A3(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n994), .A2(new_n995), .A3(new_n997), .A4(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT109), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT109), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n949), .A2(new_n1004), .A3(new_n1001), .A4(new_n994), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n994), .A2(new_n1001), .ZN(new_n1006));
  INV_X1    g581(.A(new_n956), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1003), .A2(new_n1005), .A3(new_n968), .A4(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n937), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n1002), .A2(KEYINPUT109), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n968), .B1(new_n1011), .B2(new_n1005), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n978), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1002), .A2(KEYINPUT110), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT110), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n949), .A2(new_n1015), .A3(new_n1001), .A4(new_n994), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1014), .A2(new_n1008), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n969), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1018), .A2(KEYINPUT43), .A3(new_n937), .A4(new_n1009), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1013), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT44), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT43), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1018), .A2(new_n978), .A3(new_n937), .A4(new_n1009), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT44), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1021), .A2(new_n1026), .ZN(G397));
  INV_X1    g602(.A(G1384), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n923), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT45), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n1032));
  INV_X1    g607(.A(G40), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1032), .B1(new_n795), .B2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(G160), .A2(KEYINPUT111), .A3(G40), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1031), .A2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n848), .B(new_n854), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1996), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1040), .B1(new_n801), .B2(new_n805), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n806), .A2(G1996), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n1039), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n762), .A2(new_n765), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n762), .A2(new_n765), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1047), .B1(G1986), .B2(G290), .ZN(new_n1048));
  INV_X1    g623(.A(G1986), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n601), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1037), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(G8), .B1(new_n1036), .B2(new_n1029), .ZN(new_n1052));
  XNOR2_X1  g627(.A(new_n1052), .B(KEYINPUT112), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n587), .B1(new_n589), .B2(new_n519), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(G1981), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n587), .B(new_n727), .C1(new_n588), .C2(new_n589), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT49), .B1(new_n1058), .B2(KEYINPUT116), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT115), .B1(KEYINPUT116), .B2(KEYINPUT49), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1060), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1053), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  OAI211_X1 g639(.A(KEYINPUT117), .B(new_n1053), .C1(new_n1059), .C2(new_n1061), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n962), .A2(G1976), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1053), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT52), .B1(G288), .B2(new_n717), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n1069), .B(KEYINPUT114), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1064), .A2(new_n1065), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT113), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT52), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1072), .B1(new_n1068), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1067), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G8), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT50), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n923), .A2(new_n1078), .A3(new_n1028), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT111), .B1(G160), .B2(G40), .ZN(new_n1080));
  AND4_X1   g655(.A1(KEYINPUT111), .A2(new_n793), .A3(new_n794), .A4(G40), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n500), .A2(new_n1028), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT50), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1079), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n1085), .A2(G2090), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1083), .A2(new_n1030), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1082), .B(new_n1087), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1088));
  INV_X1    g663(.A(G1971), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1077), .B1(new_n1086), .B2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(G166), .A2(new_n1077), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1092), .B(KEYINPUT55), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1036), .B1(new_n1029), .B2(KEYINPUT50), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT119), .B1(new_n1083), .B2(KEYINPUT50), .ZN(new_n1096));
  AOI21_X1  g671(.A(G1384), .B1(new_n491), .B2(new_n499), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT119), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1097), .A2(new_n1098), .A3(new_n1078), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1095), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1090), .B1(new_n1101), .B2(G2090), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1102), .A2(G8), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(new_n1093), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1071), .A2(new_n1076), .A3(new_n1094), .A4(new_n1105), .ZN(new_n1106));
  XOR2_X1   g681(.A(KEYINPUT56), .B(G2072), .Z(new_n1107));
  OR2_X1    g682(.A1(new_n1088), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT120), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1109), .B1(new_n1101), .B2(new_n773), .ZN(new_n1110));
  AOI211_X1 g685(.A(KEYINPUT120), .B(G1956), .C1(new_n1095), .C2(new_n1100), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1108), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(G299), .B(KEYINPUT57), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1113), .B(KEYINPUT122), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1113), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1115), .B(new_n1108), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1116));
  OAI21_X1  g691(.A(KEYINPUT121), .B1(new_n1036), .B2(new_n1029), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT121), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n489), .A2(new_n490), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT105), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n920), .ZN(new_n1121));
  AOI21_X1  g696(.A(G1384), .B1(new_n1121), .B2(new_n499), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1082), .A2(new_n1118), .A3(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1117), .A2(new_n854), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(G1348), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1085), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n617), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1112), .A2(new_n1114), .B1(new_n1116), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n617), .B(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1130), .A2(KEYINPUT60), .A3(new_n1124), .A4(new_n1126), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1124), .A2(new_n1126), .A3(KEYINPUT60), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT60), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1129), .B1(new_n608), .B2(new_n612), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1131), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1137));
  XNOR2_X1  g712(.A(KEYINPUT58), .B(G1341), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1138), .B1(new_n1117), .B2(new_n1123), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1088), .A2(G1996), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n554), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1142), .A2(KEYINPUT123), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  OAI221_X1 g719(.A(new_n554), .B1(KEYINPUT123), .B2(new_n1142), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1136), .A2(new_n1137), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1116), .A2(KEYINPUT61), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1099), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1098), .B1(new_n1097), .B2(new_n1078), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1082), .B1(new_n1122), .B2(new_n1078), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n773), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT120), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1101), .A2(new_n1109), .A3(new_n773), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1156), .A2(new_n1157), .A3(new_n1115), .A4(new_n1108), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1148), .A2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1128), .B1(new_n1147), .B2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1031), .B(new_n1082), .C1(new_n1030), .C2(new_n1083), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(new_n830), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1162), .B(G168), .C1(G2084), .C2(new_n1085), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(G8), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT51), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(KEYINPUT125), .A2(KEYINPUT51), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1164), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1163), .A2(new_n1165), .A3(new_n1166), .A4(G8), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1085), .ZN(new_n1171));
  AOI22_X1  g746(.A1(new_n1161), .A2(new_n830), .B1(new_n1171), .B2(new_n797), .ZN(new_n1172));
  OR3_X1    g747(.A1(new_n1172), .A2(new_n1077), .A3(G168), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1169), .A2(new_n1170), .A3(new_n1173), .ZN(new_n1174));
  OR2_X1    g749(.A1(new_n1088), .A2(G2078), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT53), .ZN(new_n1176));
  AOI22_X1  g751(.A1(new_n1175), .A2(new_n1176), .B1(new_n819), .B2(new_n1085), .ZN(new_n1177));
  XOR2_X1   g752(.A(G171), .B(KEYINPUT54), .Z(new_n1178));
  INV_X1    g753(.A(new_n1178), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1176), .A2(G2078), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1180), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1181), .B1(new_n1122), .B2(KEYINPUT45), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1182), .A2(new_n1031), .A3(G40), .A4(G160), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1177), .A2(new_n1179), .A3(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1177), .B1(new_n1161), .B2(new_n1181), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(new_n1178), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1160), .A2(new_n1174), .A3(new_n1184), .A4(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1174), .A2(KEYINPUT62), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT62), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1169), .A2(new_n1170), .A3(new_n1189), .A4(new_n1173), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1188), .A2(G171), .A3(new_n1190), .A4(new_n1185), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1106), .B1(new_n1187), .B2(new_n1191), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1172), .A2(new_n1077), .A3(G286), .ZN(new_n1193));
  OR2_X1    g768(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1071), .A2(new_n1076), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1195), .A2(KEYINPUT63), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT63), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1193), .A2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1094), .B1(new_n1104), .B2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1071), .A2(new_n1199), .A3(new_n1076), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1053), .B(KEYINPUT118), .ZN(new_n1201));
  AOI211_X1 g776(.A(G1976), .B(G288), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1056), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1201), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1196), .A2(new_n1200), .A3(new_n1204), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1051), .B1(new_n1192), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(new_n1037), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT46), .ZN(new_n1209));
  OAI22_X1  g784(.A1(new_n1207), .A2(G1996), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1037), .B1(new_n806), .B2(new_n1039), .ZN(new_n1212));
  NAND4_X1  g787(.A1(new_n1037), .A2(KEYINPUT126), .A3(KEYINPUT46), .A4(new_n1040), .ZN(new_n1213));
  NAND4_X1  g788(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  XOR2_X1   g789(.A(new_n1214), .B(KEYINPUT47), .Z(new_n1215));
  NAND2_X1  g790(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1216));
  OR2_X1    g791(.A1(new_n848), .A2(G2067), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1207), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g793(.A1(new_n1037), .A2(new_n1049), .A3(new_n601), .ZN(new_n1219));
  XOR2_X1   g794(.A(new_n1219), .B(KEYINPUT48), .Z(new_n1220));
  INV_X1    g795(.A(new_n1047), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n1220), .B1(new_n1037), .B2(new_n1221), .ZN(new_n1222));
  NOR3_X1   g797(.A1(new_n1215), .A2(new_n1218), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1206), .A2(new_n1223), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g799(.A(G227), .ZN(new_n1226));
  NAND4_X1  g800(.A1(new_n707), .A2(G319), .A3(new_n673), .A4(new_n1226), .ZN(new_n1227));
  INV_X1    g801(.A(KEYINPUT127), .ZN(new_n1228));
  OAI21_X1  g802(.A(new_n940), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g803(.A(new_n1227), .ZN(new_n1230));
  NOR2_X1   g804(.A1(new_n1230), .A2(KEYINPUT127), .ZN(new_n1231));
  AOI211_X1 g805(.A(new_n1229), .B(new_n1231), .C1(new_n1022), .C2(new_n1023), .ZN(G308));
  INV_X1    g806(.A(new_n1231), .ZN(new_n1233));
  NAND2_X1  g807(.A1(new_n1230), .A2(KEYINPUT127), .ZN(new_n1234));
  NAND4_X1  g808(.A1(new_n1024), .A2(new_n1233), .A3(new_n940), .A4(new_n1234), .ZN(G225));
endmodule


