//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 1 1 0 1 0 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 1 0 1 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n446, new_n449, new_n451, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n552, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n599, new_n601, new_n602, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1148,
    new_n1149;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  NAND2_X1  g023(.A1(G94), .A2(G452), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT67), .Z(G173));
  NAND2_X1  g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g027(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  NOR4_X1   g031(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT68), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT69), .Z(G261));
  INV_X1    g035(.A(G261), .ZN(G325));
  INV_X1    g036(.A(G2106), .ZN(new_n462));
  OR2_X1    g037(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G567), .ZN(new_n464));
  OR2_X1    g039(.A1(new_n458), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(G319));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  INV_X1    g043(.A(G113), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(G125), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT70), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n477), .A2(KEYINPUT70), .A3(G125), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n468), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(new_n470), .ZN(new_n481));
  NAND2_X1  g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  AOI21_X1  g057(.A(G2105), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G137), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT71), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n485), .B1(new_n470), .B2(G2105), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n468), .A2(KEYINPUT71), .A3(G2104), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G101), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n479), .A2(new_n490), .ZN(G160));
  NAND2_X1  g066(.A1(new_n483), .A2(G136), .ZN(new_n492));
  OR2_X1    g067(.A1(G100), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n494));
  INV_X1    g069(.A(G124), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n477), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n492), .B(new_n494), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G162));
  NAND2_X1  g073(.A1(G126), .A2(G2105), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n468), .A2(G138), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT72), .A2(KEYINPUT4), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OR2_X1    g077(.A1(new_n468), .A2(G114), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n502), .A2(new_n477), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  OAI211_X1 g081(.A(G138), .B(new_n468), .C1(new_n472), .C2(new_n473), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(new_n501), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(KEYINPUT73), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(KEYINPUT5), .A3(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(new_n518), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n511), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n521), .A2(new_n522), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n516), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n519), .A2(new_n528), .ZN(G166));
  NAND3_X1  g104(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n523), .A2(G51), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n513), .A2(new_n515), .B1(new_n521), .B2(new_n522), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G89), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n534), .A2(new_n536), .ZN(G168));
  AOI22_X1  g112(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT74), .ZN(new_n539));
  OR3_X1    g114(.A1(new_n538), .A2(new_n539), .A3(new_n518), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n538), .B2(new_n518), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n535), .A2(G90), .B1(new_n523), .B2(G52), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  NAND2_X1  g119(.A1(new_n523), .A2(G43), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n526), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n547), .B1(G651), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n552));
  XOR2_X1   g127(.A(new_n552), .B(KEYINPUT75), .Z(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  INV_X1    g131(.A(new_n523), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT76), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G53), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT9), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n523), .A2(new_n558), .A3(new_n561), .A4(G53), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n560), .A2(new_n562), .B1(G91), .B2(new_n535), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n516), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n564), .A2(new_n518), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(G299));
  INV_X1    g141(.A(G168), .ZN(G286));
  INV_X1    g142(.A(G166), .ZN(G303));
  NAND2_X1  g143(.A1(new_n535), .A2(G87), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n523), .A2(G49), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(G288));
  AOI22_X1  g147(.A1(new_n535), .A2(G86), .B1(new_n523), .B2(G48), .ZN(new_n573));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n513), .B2(new_n515), .ZN(new_n575));
  AND2_X1   g150(.A1(G73), .A2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n573), .A2(new_n577), .ZN(G305));
  AOI22_X1  g153(.A1(new_n535), .A2(G85), .B1(new_n523), .B2(G47), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n518), .B2(new_n580), .ZN(G290));
  NAND2_X1  g156(.A1(G301), .A2(G868), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n535), .A2(G92), .ZN(new_n583));
  XOR2_X1   g158(.A(new_n583), .B(KEYINPUT10), .Z(new_n584));
  AOI22_X1  g159(.A1(new_n516), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n518), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n557), .A2(KEYINPUT77), .ZN(new_n587));
  INV_X1    g162(.A(G54), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(new_n557), .B2(KEYINPUT77), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n586), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n582), .B1(new_n592), .B2(G868), .ZN(G284));
  OAI21_X1  g168(.A(new_n582), .B1(new_n592), .B2(G868), .ZN(G321));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(G299), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n596), .B1(new_n595), .B2(G168), .ZN(G297));
  XNOR2_X1  g172(.A(G297), .B(KEYINPUT78), .ZN(G280));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n592), .B1(new_n599), .B2(G860), .ZN(G148));
  NAND2_X1  g175(.A1(new_n592), .A2(new_n599), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G868), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n602), .A2(KEYINPUT79), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(KEYINPUT79), .ZN(new_n604));
  OAI211_X1 g179(.A(new_n603), .B(new_n604), .C1(G868), .C2(new_n550), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g181(.A1(new_n483), .A2(G135), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n468), .A2(G111), .ZN(new_n608));
  OAI21_X1  g183(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n609));
  INV_X1    g184(.A(G123), .ZN(new_n610));
  OAI221_X1 g185(.A(new_n607), .B1(new_n608), .B2(new_n609), .C1(new_n610), .C2(new_n496), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(G2096), .Z(new_n612));
  NAND2_X1  g187(.A1(new_n488), .A2(new_n477), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT12), .Z(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n612), .B1(new_n615), .B2(G2100), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(G2100), .B2(new_n615), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT80), .Z(G156));
  XNOR2_X1  g193(.A(G2427), .B(G2438), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2430), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT15), .B(G2435), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n622), .A2(KEYINPUT14), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2451), .B(G2454), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT16), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n624), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2443), .B(G2446), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G1341), .B(G1348), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT81), .Z(new_n632));
  NAND2_X1  g207(.A1(new_n629), .A2(new_n630), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n632), .A2(G14), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT82), .ZN(G401));
  XNOR2_X1  g210(.A(G2084), .B(G2090), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT83), .Z(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2067), .B(G2678), .ZN(new_n639));
  NOR2_X1   g214(.A1(G2072), .A2(G2078), .ZN(new_n640));
  OAI211_X1 g215(.A(new_n638), .B(new_n639), .C1(new_n444), .C2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT18), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n639), .B(KEYINPUT84), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n444), .A2(new_n640), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(KEYINPUT17), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n645), .B(new_n637), .C1(new_n643), .C2(new_n646), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n638), .A2(new_n643), .A3(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n642), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2096), .B(G2100), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT85), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n649), .B(new_n651), .ZN(G227));
  XNOR2_X1  g227(.A(G1956), .B(G2474), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT87), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1961), .B(G1966), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT86), .B(KEYINPUT19), .Z(new_n657));
  XNOR2_X1  g232(.A(G1971), .B(G1976), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT20), .Z(new_n661));
  NAND2_X1  g236(.A1(new_n654), .A2(new_n655), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n662), .A2(new_n659), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT88), .Z(new_n664));
  NAND3_X1  g239(.A1(new_n656), .A2(new_n659), .A3(new_n662), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n661), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1991), .B(G1996), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1981), .B(G1986), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G229));
  INV_X1    g247(.A(G29), .ZN(new_n673));
  INV_X1    g248(.A(G34), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n674), .A2(KEYINPUT24), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(KEYINPUT24), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n673), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(G160), .B2(new_n673), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT96), .Z(new_n679));
  NOR2_X1   g254(.A1(new_n679), .A2(G2084), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT30), .B(G28), .ZN(new_n681));
  OR2_X1    g256(.A1(KEYINPUT31), .A2(G11), .ZN(new_n682));
  NAND2_X1  g257(.A1(KEYINPUT31), .A2(G11), .ZN(new_n683));
  AOI22_X1  g258(.A1(new_n681), .A2(new_n673), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(new_n611), .B2(new_n673), .ZN(new_n685));
  NAND2_X1  g260(.A1(G164), .A2(G29), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(G27), .B2(G29), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n685), .B1(new_n687), .B2(new_n443), .ZN(new_n688));
  NAND2_X1  g263(.A1(G168), .A2(G16), .ZN(new_n689));
  NOR2_X1   g264(.A1(G16), .A2(G21), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n689), .B1(KEYINPUT98), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(KEYINPUT98), .B2(new_n689), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT99), .B(G1966), .ZN(new_n693));
  OAI221_X1 g268(.A(new_n688), .B1(new_n443), .B2(new_n687), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  AOI211_X1 g269(.A(new_n680), .B(new_n694), .C1(new_n692), .C2(new_n693), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n679), .A2(G2084), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NOR2_X1   g273(.A1(G171), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G5), .B2(new_n698), .ZN(new_n700));
  INV_X1    g275(.A(G1961), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  NAND3_X1  g278(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT26), .Z(new_n705));
  INV_X1    g280(.A(G129), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n496), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G105), .B2(new_n488), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n483), .A2(G141), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT97), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n712), .A2(new_n673), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n673), .B2(G32), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT27), .B(G1996), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n673), .A2(G33), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT95), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT25), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n483), .A2(G139), .ZN(new_n720));
  AOI22_X1  g295(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n719), .B(new_n720), .C1(new_n468), .C2(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n716), .B1(new_n722), .B2(G29), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n714), .A2(new_n715), .B1(new_n442), .B2(new_n723), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n442), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n724), .B(new_n725), .C1(new_n714), .C2(new_n715), .ZN(new_n726));
  NOR4_X1   g301(.A1(new_n697), .A2(new_n702), .A3(new_n703), .A4(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT100), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  MUX2_X1   g304(.A(G6), .B(G305), .S(G16), .Z(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT89), .Z(new_n731));
  XOR2_X1   g306(.A(KEYINPUT32), .B(G1981), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT90), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(G16), .A2(G23), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT91), .Z(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G288), .B2(new_n698), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT33), .ZN(new_n738));
  INV_X1    g313(.A(G1976), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n698), .A2(G22), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G166), .B2(new_n698), .ZN(new_n742));
  INV_X1    g317(.A(G1971), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n731), .A2(new_n733), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n734), .A2(new_n740), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n746), .A2(KEYINPUT34), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(KEYINPUT34), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n483), .A2(G131), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n468), .A2(G107), .ZN(new_n750));
  OAI21_X1  g325(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n751));
  INV_X1    g326(.A(G119), .ZN(new_n752));
  OAI221_X1 g327(.A(new_n749), .B1(new_n750), .B2(new_n751), .C1(new_n752), .C2(new_n496), .ZN(new_n753));
  MUX2_X1   g328(.A(G25), .B(new_n753), .S(G29), .Z(new_n754));
  XOR2_X1   g329(.A(KEYINPUT35), .B(G1991), .Z(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n754), .B(new_n756), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n698), .A2(G24), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G290), .B2(G16), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n760), .A2(G1986), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n760), .A2(G1986), .ZN(new_n762));
  NOR3_X1   g337(.A1(new_n757), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n747), .A2(new_n748), .A3(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT36), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n727), .A2(new_n728), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n698), .A2(G4), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n592), .B2(new_n698), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1348), .ZN(new_n769));
  AOI21_X1  g344(.A(KEYINPUT23), .B1(new_n698), .B2(G20), .ZN(new_n770));
  AND3_X1   g345(.A1(new_n698), .A2(KEYINPUT23), .A3(G20), .ZN(new_n771));
  AOI211_X1 g346(.A(new_n770), .B(new_n771), .C1(G299), .C2(G16), .ZN(new_n772));
  INV_X1    g347(.A(G1956), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n698), .A2(G19), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n550), .B2(new_n698), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(G1341), .Z(new_n777));
  NAND2_X1  g352(.A1(new_n673), .A2(G35), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G162), .B2(new_n673), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT29), .B(G2090), .Z(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n772), .A2(new_n773), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n774), .A2(new_n777), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n673), .A2(G26), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT93), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT28), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n483), .A2(G140), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n468), .A2(G116), .ZN(new_n788));
  OAI21_X1  g363(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n789));
  INV_X1    g364(.A(G128), .ZN(new_n790));
  OAI221_X1 g365(.A(new_n787), .B1(new_n788), .B2(new_n789), .C1(new_n790), .C2(new_n496), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(G29), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n792), .A2(KEYINPUT92), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n792), .A2(KEYINPUT92), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n786), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT94), .B(G2067), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NOR3_X1   g372(.A1(new_n769), .A2(new_n783), .A3(new_n797), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n729), .A2(new_n765), .A3(new_n766), .A4(new_n798), .ZN(G150));
  INV_X1    g374(.A(G150), .ZN(G311));
  NAND2_X1  g375(.A1(new_n592), .A2(G559), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT38), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n535), .A2(G93), .B1(new_n523), .B2(G55), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n518), .B2(new_n804), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n550), .B(new_n805), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n802), .B(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT39), .ZN(new_n808));
  AOI21_X1  g383(.A(G860), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n808), .B2(new_n807), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n805), .A2(G860), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT37), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT101), .ZN(G145));
  NOR2_X1   g389(.A1(new_n722), .A2(KEYINPUT102), .ZN(new_n815));
  XNOR2_X1  g390(.A(G164), .B(new_n791), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n815), .B1(new_n711), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n711), .B2(new_n816), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n722), .A2(KEYINPUT102), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(G130), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n468), .A2(G118), .ZN(new_n822));
  OAI21_X1  g397(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n823));
  OAI22_X1  g398(.A1(new_n496), .A2(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G142), .B2(new_n483), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n614), .B(new_n825), .Z(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(new_n753), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n820), .B(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(G160), .B(new_n611), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(G162), .ZN(new_n830));
  AOI21_X1  g405(.A(G37), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(new_n830), .B2(new_n828), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g408(.A(G290), .B(G305), .Z(new_n834));
  XNOR2_X1  g409(.A(G166), .B(G288), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT42), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(KEYINPUT103), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n601), .B(new_n806), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n591), .B(G299), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(KEYINPUT41), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n842), .B2(new_n839), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n838), .B(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n837), .A2(KEYINPUT103), .ZN(new_n845));
  OAI21_X1  g420(.A(G868), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n805), .A2(new_n595), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(G295));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n847), .ZN(G331));
  XNOR2_X1  g424(.A(G286), .B(G301), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(new_n806), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(KEYINPUT105), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT105), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n850), .A2(new_n806), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n850), .A2(new_n806), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(new_n842), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n851), .B(KEYINPUT106), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n856), .A2(new_n840), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n859), .A2(new_n836), .A3(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(G37), .ZN(new_n864));
  AND2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT43), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n836), .B1(new_n859), .B2(new_n862), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n865), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n863), .A2(new_n864), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n860), .A2(new_n857), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n842), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n855), .A2(new_n861), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n836), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(KEYINPUT43), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n869), .A2(new_n875), .A3(KEYINPUT44), .ZN(new_n876));
  XNOR2_X1  g451(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n872), .A2(new_n873), .ZN(new_n879));
  INV_X1    g454(.A(new_n836), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n865), .A2(new_n866), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(KEYINPUT43), .B1(new_n870), .B2(new_n867), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n878), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(KEYINPUT107), .B1(new_n876), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n883), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n877), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT107), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n869), .A2(KEYINPUT44), .A3(new_n875), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n885), .A2(new_n890), .ZN(G397));
  INV_X1    g466(.A(G125), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n892), .B1(new_n481), .B2(new_n482), .ZN(new_n893));
  OAI22_X1  g468(.A1(new_n893), .A2(KEYINPUT70), .B1(new_n469), .B2(new_n470), .ZN(new_n894));
  INV_X1    g469(.A(new_n478), .ZN(new_n895));
  OAI21_X1  g470(.A(G2105), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n490), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(G40), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(G1384), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n502), .A2(new_n477), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n503), .A2(new_n505), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n507), .A2(new_n501), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n899), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT45), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n898), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(G1996), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n909), .A2(KEYINPUT46), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(KEYINPUT46), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n791), .B(G2067), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n912), .A2(new_n711), .ZN(new_n913));
  AOI22_X1  g488(.A1(new_n910), .A2(new_n911), .B1(new_n907), .B2(new_n913), .ZN(new_n914));
  XOR2_X1   g489(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n915));
  XNOR2_X1  g490(.A(new_n914), .B(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n909), .A2(new_n711), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT108), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n712), .A2(new_n908), .ZN(new_n919));
  OR2_X1    g494(.A1(new_n919), .A2(new_n912), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n918), .B1(new_n907), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n907), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n753), .B(new_n755), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n922), .A2(G1986), .A3(G290), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT48), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n916), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n753), .A2(new_n756), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n921), .A2(new_n928), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n791), .A2(G2067), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n922), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT126), .ZN(new_n933));
  XNOR2_X1  g508(.A(G290), .B(G1986), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n924), .B1(new_n907), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(G40), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n479), .A2(new_n936), .A3(new_n490), .ZN(new_n937));
  AOI21_X1  g512(.A(G1384), .B1(new_n506), .B2(new_n508), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(KEYINPUT45), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n906), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n743), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT50), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n898), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT115), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n945), .B1(new_n938), .B2(new_n942), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n938), .A2(new_n945), .A3(new_n942), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n941), .B1(new_n948), .B2(G2090), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(G8), .ZN(new_n950));
  NAND2_X1  g525(.A1(G303), .A2(G8), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(KEYINPUT55), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n952), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT110), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n509), .A2(new_n942), .A3(new_n899), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n904), .A2(KEYINPUT50), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n938), .A2(KEYINPUT109), .A3(new_n942), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n958), .A2(new_n937), .A3(new_n959), .A4(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n955), .B1(new_n961), .B2(G2090), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n938), .A2(KEYINPUT109), .A3(new_n942), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT109), .B1(new_n938), .B2(new_n942), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G2090), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n965), .A2(KEYINPUT110), .A3(new_n966), .A4(new_n944), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n962), .A2(new_n967), .A3(new_n941), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n954), .A2(new_n968), .A3(G8), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n953), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G288), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(G1976), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n896), .A2(new_n938), .A3(G40), .A4(new_n897), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT111), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n973), .A2(new_n974), .A3(G8), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n974), .B1(new_n973), .B2(G8), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n972), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT112), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT112), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n979), .B(new_n972), .C1(new_n975), .C2(new_n976), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n978), .A2(new_n980), .A3(KEYINPUT52), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n973), .A2(G8), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT111), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n973), .A2(new_n974), .A3(G8), .ZN(new_n984));
  AOI22_X1  g559(.A1(new_n983), .A2(new_n984), .B1(G1976), .B2(new_n971), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT52), .B1(G288), .B2(new_n739), .ZN(new_n986));
  INV_X1    g561(.A(G1981), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n535), .A2(G86), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n523), .A2(G48), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n577), .A2(new_n987), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT113), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n573), .A2(KEYINPUT113), .A3(new_n577), .A4(new_n987), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n987), .B1(new_n573), .B2(new_n577), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT49), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT49), .ZN(new_n998));
  AOI211_X1 g573(.A(new_n998), .B(new_n995), .C1(new_n992), .C2(new_n993), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n983), .A2(new_n984), .ZN(new_n1001));
  AOI22_X1  g576(.A1(new_n985), .A2(new_n986), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n981), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n937), .A2(new_n906), .A3(new_n443), .A4(new_n939), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n1004), .B(KEYINPUT53), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n961), .A2(KEYINPUT120), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT120), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n944), .A2(new_n1007), .A3(new_n958), .A4(new_n960), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n1008), .A3(new_n701), .ZN(new_n1009));
  AOI21_X1  g584(.A(G301), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n970), .A2(new_n1003), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n1012));
  XOR2_X1   g587(.A(KEYINPUT116), .B(G2084), .Z(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n961), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G1966), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n940), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(G8), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1012), .B1(new_n1018), .B2(KEYINPUT124), .ZN(new_n1019));
  OAI21_X1  g594(.A(G286), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n965), .A2(new_n944), .A3(new_n1013), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n940), .A2(new_n1016), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(G168), .A3(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1020), .A2(G8), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G8), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT124), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT51), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1023), .A2(G8), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1025), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT62), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT62), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1025), .A2(new_n1034), .A3(new_n1031), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1011), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n969), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n981), .A2(new_n1002), .A3(KEYINPUT114), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT114), .B1(new_n981), .B2(new_n1002), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1037), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AOI211_X1 g615(.A(G1976), .B(G288), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1041));
  INV_X1    g616(.A(new_n994), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1001), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G1348), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1006), .A2(new_n1008), .A3(new_n1046), .ZN(new_n1047));
  OR2_X1    g622(.A1(new_n973), .A2(G2067), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n592), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n947), .A2(new_n946), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n937), .A2(new_n959), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n773), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n937), .A2(new_n906), .A3(new_n939), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT56), .B(G2072), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT57), .ZN(new_n1058));
  XNOR2_X1  g633(.A(G299), .B(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1053), .A2(new_n1059), .A3(new_n1056), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT119), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1053), .A2(new_n1059), .A3(new_n1056), .A4(new_n1064), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n1050), .A2(new_n1061), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1061), .A2(KEYINPUT61), .A3(new_n1062), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1059), .B1(new_n1053), .B2(new_n1056), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1068), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1067), .B1(new_n1069), .B2(KEYINPUT61), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1047), .A2(KEYINPUT60), .A3(new_n1048), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n592), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1047), .A2(KEYINPUT60), .A3(new_n591), .A4(new_n1048), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT60), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1072), .A2(new_n1073), .B1(new_n1074), .B2(new_n1049), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1070), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT123), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1078), .B(G1341), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n973), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n973), .A2(KEYINPUT122), .A3(new_n1079), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(new_n940), .B2(G1996), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1077), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1054), .A2(new_n908), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1087), .A2(new_n1084), .A3(KEYINPUT123), .A4(new_n1082), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n550), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT59), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1089), .A2(new_n1092), .A3(new_n550), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1066), .B1(new_n1076), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n970), .A2(new_n1003), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT125), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1005), .A2(new_n1009), .A3(G301), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1098), .B1(new_n1099), .B2(new_n1010), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(KEYINPUT54), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT54), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1098), .B(new_n1102), .C1(new_n1099), .C2(new_n1010), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1097), .A2(new_n1101), .A3(new_n1032), .A4(new_n1103), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1036), .B(new_n1045), .C1(new_n1095), .C2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT63), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1018), .A2(G286), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1106), .B1(new_n1096), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n968), .A2(G8), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT117), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n968), .A2(KEYINPUT117), .A3(G8), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(new_n952), .A3(new_n1114), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1115), .B(KEYINPUT118), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n969), .A2(new_n1107), .A3(KEYINPUT63), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1115), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1117), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1110), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n933), .B(new_n935), .C1(new_n1105), .C2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1117), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1124), .A2(new_n1116), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n1109), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1075), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n948), .A2(new_n773), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1064), .B1(new_n1129), .B2(new_n1059), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1065), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1061), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT61), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1128), .A2(new_n1094), .A3(new_n1134), .A4(new_n1067), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1066), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1101), .A2(new_n1032), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1103), .A2(new_n970), .A3(new_n1003), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1044), .B1(new_n1142), .B2(new_n1011), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1127), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n933), .B1(new_n1144), .B2(new_n935), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n932), .B1(new_n1123), .B2(new_n1145), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g721(.A(G401), .ZN(new_n1148));
  NOR3_X1   g722(.A1(G229), .A2(new_n466), .A3(G227), .ZN(new_n1149));
  AND4_X1   g723(.A1(new_n1148), .A2(new_n832), .A3(new_n1149), .A4(new_n886), .ZN(G308));
  NAND4_X1  g724(.A1(new_n1148), .A2(new_n832), .A3(new_n1149), .A4(new_n886), .ZN(G225));
endmodule


