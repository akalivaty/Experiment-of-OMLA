

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XOR2_X1 U323 ( .A(G50GAT), .B(G162GAT), .Z(n430) );
  XOR2_X1 U324 ( .A(G43GAT), .B(G134GAT), .Z(n438) );
  NAND2_X1 U325 ( .A1(n471), .A2(n470), .ZN(n473) );
  XOR2_X1 U326 ( .A(n408), .B(n407), .Z(n291) );
  XOR2_X1 U327 ( .A(G92GAT), .B(G218GAT), .Z(n292) );
  AND2_X1 U328 ( .A1(G232GAT), .A2(G233GAT), .ZN(n293) );
  XOR2_X1 U329 ( .A(KEYINPUT37), .B(n488), .Z(n294) );
  INV_X1 U330 ( .A(n527), .ZN(n416) );
  NAND2_X1 U331 ( .A1(n416), .A2(n518), .ZN(n417) );
  XNOR2_X1 U332 ( .A(n364), .B(n293), .ZN(n304) );
  INV_X1 U333 ( .A(KEYINPUT98), .ZN(n472) );
  XNOR2_X1 U334 ( .A(n417), .B(KEYINPUT54), .ZN(n418) );
  XNOR2_X1 U335 ( .A(n305), .B(n304), .ZN(n309) );
  XNOR2_X1 U336 ( .A(n473), .B(n472), .ZN(n486) );
  XNOR2_X1 U337 ( .A(n437), .B(n436), .ZN(n452) );
  INV_X1 U338 ( .A(G190GAT), .ZN(n453) );
  XOR2_X1 U339 ( .A(KEYINPUT79), .B(n557), .Z(n541) );
  XNOR2_X1 U340 ( .A(n453), .B(KEYINPUT58), .ZN(n454) );
  XNOR2_X1 U341 ( .A(n455), .B(n454), .ZN(G1351GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT77), .B(KEYINPUT9), .Z(n296) );
  XNOR2_X1 U343 ( .A(KEYINPUT78), .B(KEYINPUT10), .ZN(n295) );
  XOR2_X1 U344 ( .A(n296), .B(n295), .Z(n300) );
  XOR2_X1 U345 ( .A(KEYINPUT11), .B(KEYINPUT64), .Z(n298) );
  XNOR2_X1 U346 ( .A(n438), .B(n430), .ZN(n297) );
  XNOR2_X1 U347 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U348 ( .A(n300), .B(n299), .ZN(n305) );
  XOR2_X1 U349 ( .A(KEYINPUT74), .B(KEYINPUT75), .Z(n302) );
  XNOR2_X1 U350 ( .A(G106GAT), .B(G85GAT), .ZN(n301) );
  XNOR2_X1 U351 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U352 ( .A(G99GAT), .B(n303), .Z(n364) );
  XNOR2_X1 U353 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n306), .B(KEYINPUT7), .ZN(n336) );
  XNOR2_X1 U355 ( .A(G36GAT), .B(G190GAT), .ZN(n307) );
  XNOR2_X1 U356 ( .A(n292), .B(n307), .ZN(n404) );
  XNOR2_X1 U357 ( .A(n336), .B(n404), .ZN(n308) );
  XNOR2_X1 U358 ( .A(n309), .B(n308), .ZN(n557) );
  XOR2_X1 U359 ( .A(KEYINPUT92), .B(KEYINPUT4), .Z(n311) );
  XNOR2_X1 U360 ( .A(G57GAT), .B(KEYINPUT94), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n311), .B(n310), .ZN(n317) );
  XOR2_X1 U362 ( .A(G127GAT), .B(KEYINPUT0), .Z(n313) );
  XNOR2_X1 U363 ( .A(G113GAT), .B(KEYINPUT83), .ZN(n312) );
  XNOR2_X1 U364 ( .A(n313), .B(n312), .ZN(n439) );
  XOR2_X1 U365 ( .A(n439), .B(KEYINPUT5), .Z(n315) );
  NAND2_X1 U366 ( .A1(G225GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U368 ( .A(n317), .B(n316), .ZN(n332) );
  XOR2_X1 U369 ( .A(KEYINPUT95), .B(G148GAT), .Z(n319) );
  XNOR2_X1 U370 ( .A(G141GAT), .B(G120GAT), .ZN(n318) );
  XNOR2_X1 U371 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U372 ( .A(KEYINPUT6), .B(KEYINPUT93), .Z(n321) );
  XNOR2_X1 U373 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U375 ( .A(n323), .B(n322), .Z(n330) );
  XOR2_X1 U376 ( .A(G85GAT), .B(G162GAT), .Z(n327) );
  XOR2_X1 U377 ( .A(G155GAT), .B(KEYINPUT2), .Z(n325) );
  XNOR2_X1 U378 ( .A(KEYINPUT89), .B(KEYINPUT3), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n325), .B(n324), .ZN(n423) );
  XNOR2_X1 U380 ( .A(G29GAT), .B(n423), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U382 ( .A(G134GAT), .B(n328), .ZN(n329) );
  XNOR2_X1 U383 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n332), .B(n331), .ZN(n516) );
  XNOR2_X1 U385 ( .A(KEYINPUT114), .B(KEYINPUT47), .ZN(n390) );
  XNOR2_X1 U386 ( .A(G15GAT), .B(G1GAT), .ZN(n333) );
  XNOR2_X1 U387 ( .A(n333), .B(G8GAT), .ZN(n381) );
  XOR2_X1 U388 ( .A(G141GAT), .B(G22GAT), .Z(n431) );
  XOR2_X1 U389 ( .A(n381), .B(n431), .Z(n335) );
  XNOR2_X1 U390 ( .A(G50GAT), .B(G43GAT), .ZN(n334) );
  XNOR2_X1 U391 ( .A(n335), .B(n334), .ZN(n340) );
  XOR2_X1 U392 ( .A(n336), .B(KEYINPUT69), .Z(n338) );
  NAND2_X1 U393 ( .A1(G229GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U395 ( .A(n340), .B(n339), .Z(n348) );
  XOR2_X1 U396 ( .A(G197GAT), .B(G113GAT), .Z(n342) );
  XNOR2_X1 U397 ( .A(G169GAT), .B(G36GAT), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U399 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n344) );
  XNOR2_X1 U400 ( .A(KEYINPUT68), .B(KEYINPUT29), .ZN(n343) );
  XNOR2_X1 U401 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U402 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U403 ( .A(n348), .B(n347), .ZN(n570) );
  INV_X1 U404 ( .A(n570), .ZN(n531) );
  XOR2_X1 U405 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n350) );
  NAND2_X1 U406 ( .A1(G230GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U407 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U408 ( .A(n351), .B(KEYINPUT71), .Z(n357) );
  XOR2_X1 U409 ( .A(G78GAT), .B(G148GAT), .Z(n353) );
  XNOR2_X1 U410 ( .A(KEYINPUT73), .B(KEYINPUT72), .ZN(n352) );
  XNOR2_X1 U411 ( .A(n353), .B(n352), .ZN(n422) );
  XOR2_X1 U412 ( .A(G57GAT), .B(KEYINPUT70), .Z(n354) );
  XNOR2_X1 U413 ( .A(KEYINPUT13), .B(n354), .ZN(n382) );
  INV_X1 U414 ( .A(n382), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n422), .B(n355), .ZN(n356) );
  XNOR2_X1 U416 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U417 ( .A(KEYINPUT76), .B(G64GAT), .Z(n407) );
  XOR2_X1 U418 ( .A(KEYINPUT33), .B(n407), .Z(n359) );
  XOR2_X1 U419 ( .A(G120GAT), .B(G71GAT), .Z(n442) );
  XNOR2_X1 U420 ( .A(n442), .B(G204GAT), .ZN(n358) );
  XNOR2_X1 U421 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U422 ( .A(n361), .B(n360), .Z(n363) );
  XNOR2_X1 U423 ( .A(G176GAT), .B(G92GAT), .ZN(n362) );
  XNOR2_X1 U424 ( .A(n363), .B(n362), .ZN(n366) );
  INV_X1 U425 ( .A(n364), .ZN(n365) );
  XNOR2_X1 U426 ( .A(n366), .B(n365), .ZN(n456) );
  XNOR2_X1 U427 ( .A(n456), .B(KEYINPUT41), .ZN(n501) );
  NAND2_X1 U428 ( .A1(n531), .A2(n501), .ZN(n367) );
  XNOR2_X1 U429 ( .A(KEYINPUT46), .B(n367), .ZN(n386) );
  XOR2_X1 U430 ( .A(KEYINPUT12), .B(KEYINPUT80), .Z(n369) );
  XNOR2_X1 U431 ( .A(KEYINPUT14), .B(KEYINPUT81), .ZN(n368) );
  XNOR2_X1 U432 ( .A(n369), .B(n368), .ZN(n377) );
  NAND2_X1 U433 ( .A1(G231GAT), .A2(G233GAT), .ZN(n375) );
  XOR2_X1 U434 ( .A(G155GAT), .B(G211GAT), .Z(n371) );
  XNOR2_X1 U435 ( .A(G22GAT), .B(G127GAT), .ZN(n370) );
  XNOR2_X1 U436 ( .A(n371), .B(n370), .ZN(n373) );
  XOR2_X1 U437 ( .A(G183GAT), .B(G71GAT), .Z(n372) );
  XNOR2_X1 U438 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U439 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U440 ( .A(n377), .B(n376), .ZN(n385) );
  XOR2_X1 U441 ( .A(KEYINPUT15), .B(KEYINPUT82), .Z(n379) );
  XNOR2_X1 U442 ( .A(G78GAT), .B(G64GAT), .ZN(n378) );
  XNOR2_X1 U443 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U444 ( .A(n381), .B(n380), .ZN(n383) );
  XNOR2_X1 U445 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U446 ( .A(n385), .B(n384), .ZN(n577) );
  NAND2_X1 U447 ( .A1(n386), .A2(n577), .ZN(n387) );
  XNOR2_X1 U448 ( .A(KEYINPUT113), .B(n387), .ZN(n388) );
  NAND2_X1 U449 ( .A1(n388), .A2(n557), .ZN(n389) );
  XNOR2_X1 U450 ( .A(n390), .B(n389), .ZN(n397) );
  INV_X1 U451 ( .A(n577), .ZN(n537) );
  XOR2_X1 U452 ( .A(KEYINPUT36), .B(KEYINPUT102), .Z(n391) );
  XNOR2_X1 U453 ( .A(n541), .B(n391), .ZN(n581) );
  NAND2_X1 U454 ( .A1(n537), .A2(n581), .ZN(n393) );
  XOR2_X1 U455 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n392) );
  XNOR2_X1 U456 ( .A(n393), .B(n392), .ZN(n395) );
  NAND2_X1 U457 ( .A1(n456), .A2(n570), .ZN(n394) );
  NOR2_X1 U458 ( .A1(n395), .A2(n394), .ZN(n396) );
  NOR2_X1 U459 ( .A1(n397), .A2(n396), .ZN(n398) );
  XNOR2_X1 U460 ( .A(KEYINPUT48), .B(n398), .ZN(n527) );
  XOR2_X1 U461 ( .A(KEYINPUT17), .B(KEYINPUT85), .Z(n400) );
  XNOR2_X1 U462 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n399) );
  XNOR2_X1 U463 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U464 ( .A(n401), .B(G183GAT), .Z(n403) );
  XNOR2_X1 U465 ( .A(G169GAT), .B(G176GAT), .ZN(n402) );
  XNOR2_X1 U466 ( .A(n403), .B(n402), .ZN(n449) );
  XOR2_X1 U467 ( .A(n404), .B(KEYINPUT96), .Z(n406) );
  NAND2_X1 U468 ( .A1(G226GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U469 ( .A(n406), .B(n405), .ZN(n408) );
  XNOR2_X1 U470 ( .A(G8GAT), .B(KEYINPUT97), .ZN(n409) );
  XNOR2_X1 U471 ( .A(n291), .B(n409), .ZN(n410) );
  XNOR2_X1 U472 ( .A(n449), .B(n410), .ZN(n415) );
  XOR2_X1 U473 ( .A(KEYINPUT88), .B(G211GAT), .Z(n412) );
  XNOR2_X1 U474 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n411) );
  XNOR2_X1 U475 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U476 ( .A(G197GAT), .B(n413), .Z(n435) );
  INV_X1 U477 ( .A(n435), .ZN(n414) );
  XOR2_X1 U478 ( .A(n415), .B(n414), .Z(n518) );
  INV_X1 U479 ( .A(n518), .ZN(n458) );
  NOR2_X1 U480 ( .A1(n516), .A2(n418), .ZN(n569) );
  XOR2_X1 U481 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n420) );
  NAND2_X1 U482 ( .A1(G228GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U483 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U484 ( .A(n421), .B(KEYINPUT22), .Z(n425) );
  XNOR2_X1 U485 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U486 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U487 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n427) );
  XNOR2_X1 U488 ( .A(G218GAT), .B(G106GAT), .ZN(n426) );
  XNOR2_X1 U489 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U490 ( .A(n429), .B(n428), .Z(n433) );
  XNOR2_X1 U491 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U492 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(n464) );
  NAND2_X1 U494 ( .A1(n569), .A2(n464), .ZN(n437) );
  XOR2_X1 U495 ( .A(KEYINPUT55), .B(KEYINPUT123), .Z(n436) );
  XOR2_X1 U496 ( .A(n439), .B(n438), .Z(n441) );
  NAND2_X1 U497 ( .A1(G227GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n441), .B(n440), .ZN(n443) );
  XOR2_X1 U499 ( .A(n443), .B(n442), .Z(n445) );
  XNOR2_X1 U500 ( .A(G99GAT), .B(G190GAT), .ZN(n444) );
  XNOR2_X1 U501 ( .A(n445), .B(n444), .ZN(n451) );
  XOR2_X1 U502 ( .A(KEYINPUT84), .B(KEYINPUT86), .Z(n447) );
  XNOR2_X1 U503 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n446) );
  XNOR2_X1 U504 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U505 ( .A(n449), .B(n448), .Z(n450) );
  XNOR2_X1 U506 ( .A(n451), .B(n450), .ZN(n528) );
  NAND2_X1 U507 ( .A1(n452), .A2(n528), .ZN(n566) );
  NOR2_X1 U508 ( .A1(n541), .A2(n566), .ZN(n455) );
  NAND2_X1 U509 ( .A1(n456), .A2(n531), .ZN(n489) );
  XNOR2_X1 U510 ( .A(n528), .B(KEYINPUT87), .ZN(n460) );
  XOR2_X1 U511 ( .A(KEYINPUT28), .B(KEYINPUT66), .Z(n457) );
  XNOR2_X1 U512 ( .A(n464), .B(n457), .ZN(n530) );
  XOR2_X1 U513 ( .A(KEYINPUT27), .B(n458), .Z(n462) );
  NAND2_X1 U514 ( .A1(n516), .A2(n462), .ZN(n526) );
  NOR2_X1 U515 ( .A1(n530), .A2(n526), .ZN(n459) );
  NAND2_X1 U516 ( .A1(n460), .A2(n459), .ZN(n471) );
  NOR2_X1 U517 ( .A1(n464), .A2(n528), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n461), .B(KEYINPUT26), .ZN(n568) );
  NAND2_X1 U519 ( .A1(n462), .A2(n568), .ZN(n467) );
  NAND2_X1 U520 ( .A1(n518), .A2(n528), .ZN(n463) );
  NAND2_X1 U521 ( .A1(n464), .A2(n463), .ZN(n465) );
  XOR2_X1 U522 ( .A(KEYINPUT25), .B(n465), .Z(n466) );
  NAND2_X1 U523 ( .A1(n467), .A2(n466), .ZN(n469) );
  INV_X1 U524 ( .A(n516), .ZN(n468) );
  NAND2_X1 U525 ( .A1(n469), .A2(n468), .ZN(n470) );
  NAND2_X1 U526 ( .A1(n541), .A2(n537), .ZN(n474) );
  XNOR2_X1 U527 ( .A(KEYINPUT16), .B(n474), .ZN(n475) );
  OR2_X1 U528 ( .A1(n486), .A2(n475), .ZN(n502) );
  NOR2_X1 U529 ( .A1(n489), .A2(n502), .ZN(n484) );
  NAND2_X1 U530 ( .A1(n484), .A2(n516), .ZN(n478) );
  XOR2_X1 U531 ( .A(G1GAT), .B(KEYINPUT34), .Z(n476) );
  XNOR2_X1 U532 ( .A(KEYINPUT99), .B(n476), .ZN(n477) );
  XNOR2_X1 U533 ( .A(n478), .B(n477), .ZN(G1324GAT) );
  NAND2_X1 U534 ( .A1(n484), .A2(n518), .ZN(n479) );
  XNOR2_X1 U535 ( .A(n479), .B(KEYINPUT100), .ZN(n480) );
  XNOR2_X1 U536 ( .A(G8GAT), .B(n480), .ZN(G1325GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n482) );
  NAND2_X1 U538 ( .A1(n484), .A2(n528), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U540 ( .A(G15GAT), .B(n483), .Z(G1326GAT) );
  NAND2_X1 U541 ( .A1(n484), .A2(n530), .ZN(n485) );
  XNOR2_X1 U542 ( .A(n485), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U543 ( .A(G29GAT), .B(KEYINPUT39), .Z(n493) );
  NOR2_X1 U544 ( .A1(n537), .A2(n486), .ZN(n487) );
  NAND2_X1 U545 ( .A1(n581), .A2(n487), .ZN(n488) );
  NOR2_X1 U546 ( .A1(n294), .A2(n489), .ZN(n491) );
  XOR2_X1 U547 ( .A(KEYINPUT38), .B(KEYINPUT103), .Z(n490) );
  XNOR2_X1 U548 ( .A(n491), .B(n490), .ZN(n499) );
  NAND2_X1 U549 ( .A1(n516), .A2(n499), .ZN(n492) );
  XNOR2_X1 U550 ( .A(n493), .B(n492), .ZN(G1328GAT) );
  NAND2_X1 U551 ( .A1(n499), .A2(n518), .ZN(n494) );
  XNOR2_X1 U552 ( .A(n494), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U553 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n498) );
  NAND2_X1 U554 ( .A1(n499), .A2(n528), .ZN(n496) );
  XOR2_X1 U555 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n495) );
  XNOR2_X1 U556 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n498), .B(n497), .ZN(G1330GAT) );
  NAND2_X1 U558 ( .A1(n499), .A2(n530), .ZN(n500) );
  XNOR2_X1 U559 ( .A(n500), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT42), .B(KEYINPUT106), .Z(n504) );
  INV_X1 U561 ( .A(n501), .ZN(n563) );
  NAND2_X1 U562 ( .A1(n570), .A2(n501), .ZN(n515) );
  NOR2_X1 U563 ( .A1(n515), .A2(n502), .ZN(n510) );
  NAND2_X1 U564 ( .A1(n510), .A2(n516), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U566 ( .A(G57GAT), .B(n505), .Z(G1332GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n507) );
  NAND2_X1 U568 ( .A1(n510), .A2(n518), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U570 ( .A(G64GAT), .B(n508), .ZN(G1333GAT) );
  NAND2_X1 U571 ( .A1(n528), .A2(n510), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n509), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n512) );
  NAND2_X1 U574 ( .A1(n510), .A2(n530), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n512), .B(n511), .ZN(n514) );
  XOR2_X1 U576 ( .A(G78GAT), .B(KEYINPUT110), .Z(n513) );
  XNOR2_X1 U577 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  NOR2_X1 U578 ( .A1(n294), .A2(n515), .ZN(n522) );
  NAND2_X1 U579 ( .A1(n516), .A2(n522), .ZN(n517) );
  XNOR2_X1 U580 ( .A(G85GAT), .B(n517), .ZN(G1336GAT) );
  NAND2_X1 U581 ( .A1(n522), .A2(n518), .ZN(n519) );
  XNOR2_X1 U582 ( .A(n519), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U583 ( .A(G99GAT), .B(KEYINPUT111), .Z(n521) );
  NAND2_X1 U584 ( .A1(n522), .A2(n528), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n521), .B(n520), .ZN(G1338GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT44), .B(KEYINPUT112), .Z(n524) );
  NAND2_X1 U587 ( .A1(n522), .A2(n530), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U589 ( .A(G106GAT), .B(n525), .Z(G1339GAT) );
  XOR2_X1 U590 ( .A(G113GAT), .B(KEYINPUT115), .Z(n533) );
  NOR2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n547) );
  NAND2_X1 U592 ( .A1(n547), .A2(n528), .ZN(n529) );
  NOR2_X1 U593 ( .A1(n530), .A2(n529), .ZN(n540) );
  NAND2_X1 U594 ( .A1(n540), .A2(n531), .ZN(n532) );
  XNOR2_X1 U595 ( .A(n533), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n535) );
  NAND2_X1 U597 ( .A1(n540), .A2(n501), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U599 ( .A(G120GAT), .B(n536), .ZN(G1341GAT) );
  NAND2_X1 U600 ( .A1(n537), .A2(n540), .ZN(n538) );
  XNOR2_X1 U601 ( .A(n538), .B(KEYINPUT50), .ZN(n539) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(n539), .ZN(G1342GAT) );
  INV_X1 U603 ( .A(n540), .ZN(n542) );
  NOR2_X1 U604 ( .A1(n542), .A2(n541), .ZN(n546) );
  XOR2_X1 U605 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n544) );
  XNOR2_X1 U606 ( .A(G134GAT), .B(KEYINPUT118), .ZN(n543) );
  XNOR2_X1 U607 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U608 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  NAND2_X1 U609 ( .A1(n547), .A2(n568), .ZN(n556) );
  NOR2_X1 U610 ( .A1(n570), .A2(n556), .ZN(n548) );
  XOR2_X1 U611 ( .A(G141GAT), .B(n548), .Z(G1344GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n550) );
  XNOR2_X1 U613 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(n554) );
  NOR2_X1 U615 ( .A1(n563), .A2(n556), .ZN(n552) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U618 ( .A(n554), .B(n553), .Z(G1345GAT) );
  NOR2_X1 U619 ( .A1(n577), .A2(n556), .ZN(n555) );
  XOR2_X1 U620 ( .A(G155GAT), .B(n555), .Z(G1346GAT) );
  NOR2_X1 U621 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U622 ( .A(KEYINPUT122), .B(n558), .Z(n559) );
  XNOR2_X1 U623 ( .A(G162GAT), .B(n559), .ZN(G1347GAT) );
  NOR2_X1 U624 ( .A1(n570), .A2(n566), .ZN(n560) );
  XOR2_X1 U625 ( .A(G169GAT), .B(n560), .Z(G1348GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n562) );
  XNOR2_X1 U627 ( .A(G176GAT), .B(KEYINPUT124), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n565) );
  NOR2_X1 U629 ( .A1(n563), .A2(n566), .ZN(n564) );
  XOR2_X1 U630 ( .A(n565), .B(n564), .Z(G1349GAT) );
  NOR2_X1 U631 ( .A1(n577), .A2(n566), .ZN(n567) );
  XOR2_X1 U632 ( .A(G183GAT), .B(n567), .Z(G1350GAT) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n580) );
  NOR2_X1 U634 ( .A1(n580), .A2(n570), .ZN(n574) );
  XOR2_X1 U635 ( .A(KEYINPUT59), .B(KEYINPUT60), .Z(n572) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  NOR2_X1 U639 ( .A1(n456), .A2(n580), .ZN(n576) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n580), .ZN(n578) );
  XOR2_X1 U643 ( .A(KEYINPUT126), .B(n578), .Z(n579) );
  XNOR2_X1 U644 ( .A(G211GAT), .B(n579), .ZN(G1354GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n584) );
  INV_X1 U646 ( .A(n580), .ZN(n582) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

