//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n561, new_n562, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n575, new_n576, new_n577, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1181, new_n1182;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT64), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n451), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(new_n452), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n465), .A2(G137), .B1(G101), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n464), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n466), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n470), .A2(new_n474), .ZN(G160));
  OAI21_X1  g050(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(G112), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n465), .A2(G136), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n464), .A2(new_n466), .ZN(new_n481));
  AOI211_X1 g056(.A(new_n478), .B(new_n480), .C1(G124), .C2(new_n481), .ZN(G162));
  NAND2_X1  g057(.A1(new_n465), .A2(G138), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT4), .ZN(new_n484));
  OR2_X1    g059(.A1(G102), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G114), .C2(new_n466), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n481), .A2(G126), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT65), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G164));
  OR2_X1    g066(.A1(KEYINPUT5), .A2(G543), .ZN(new_n492));
  NAND2_X1  g067(.A1(KEYINPUT5), .A2(G543), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n494), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n495));
  INV_X1    g070(.A(G651), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(KEYINPUT5), .A2(G543), .ZN(new_n498));
  AND2_X1   g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  AND2_X1   g074(.A1(KEYINPUT6), .A2(G651), .ZN(new_n500));
  NOR2_X1   g075(.A1(KEYINPUT6), .A2(G651), .ZN(new_n501));
  OAI22_X1  g076(.A1(new_n498), .A2(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G88), .ZN(new_n503));
  OAI21_X1  g078(.A(G543), .B1(new_n500), .B2(new_n501), .ZN(new_n504));
  INV_X1    g079(.A(G50), .ZN(new_n505));
  OAI22_X1  g080(.A1(new_n502), .A2(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n497), .A2(new_n506), .ZN(G166));
  XOR2_X1   g082(.A(KEYINPUT67), .B(G89), .Z(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(new_n496), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n508), .A2(new_n494), .A3(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT68), .ZN(new_n514));
  NAND3_X1  g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT66), .B(KEYINPUT7), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(new_n515), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n513), .A2(new_n514), .A3(new_n519), .A4(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G543), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n523), .B1(new_n510), .B2(new_n511), .ZN(new_n524));
  AND2_X1   g099(.A1(G63), .A2(G651), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n524), .A2(G51), .B1(new_n494), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n521), .A2(new_n519), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n514), .B1(new_n528), .B2(new_n513), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n527), .A2(new_n529), .ZN(G168));
  OAI211_X1 g105(.A(G52), .B(G543), .C1(new_n500), .C2(new_n501), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT69), .B(G90), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n502), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g108(.A(G64), .B1(new_n499), .B2(new_n498), .ZN(new_n534));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n496), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g111(.A(KEYINPUT70), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G64), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n538), .B1(new_n492), .B2(new_n493), .ZN(new_n539));
  INV_X1    g114(.A(new_n535), .ZN(new_n540));
  OAI21_X1  g115(.A(G651), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT70), .ZN(new_n542));
  XOR2_X1   g117(.A(KEYINPUT69), .B(G90), .Z(new_n543));
  NAND3_X1  g118(.A1(new_n543), .A2(new_n494), .A3(new_n512), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n541), .A2(new_n542), .A3(new_n544), .A4(new_n531), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n537), .A2(new_n545), .ZN(G171));
  NOR2_X1   g121(.A1(new_n499), .A2(new_n498), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  INV_X1    g123(.A(G68), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n547), .A2(new_n548), .B1(new_n549), .B2(new_n523), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT71), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI221_X1 g127(.A(KEYINPUT71), .B1(new_n549), .B2(new_n523), .C1(new_n547), .C2(new_n548), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n552), .A2(G651), .A3(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n492), .A2(new_n493), .B1(new_n510), .B2(new_n511), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n555), .A2(G81), .B1(new_n524), .B2(G43), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT72), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n566), .B1(new_n492), .B2(new_n493), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n555), .A2(G91), .ZN(new_n569));
  OAI211_X1 g144(.A(G53), .B(G543), .C1(new_n500), .C2(new_n501), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n570), .A2(KEYINPUT9), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n570), .A2(KEYINPUT9), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n568), .B(new_n569), .C1(new_n571), .C2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  INV_X1    g149(.A(new_n513), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n521), .A2(new_n519), .ZN(new_n576));
  OAI21_X1  g151(.A(KEYINPUT68), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n577), .A2(new_n522), .A3(new_n526), .ZN(G286));
  INV_X1    g153(.A(G166), .ZN(G303));
  NAND2_X1  g154(.A1(new_n524), .A2(G49), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT73), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n494), .A2(G74), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(G87), .B2(new_n555), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(G288));
  AOI22_X1  g159(.A1(new_n494), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n496), .ZN(new_n586));
  INV_X1    g161(.A(G86), .ZN(new_n587));
  INV_X1    g162(.A(G48), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n502), .A2(new_n587), .B1(new_n504), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n494), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n496), .ZN(new_n593));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n502), .A2(new_n594), .B1(new_n504), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G290));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  NOR2_X1   g174(.A1(G171), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT74), .ZN(new_n601));
  AOI21_X1  g176(.A(KEYINPUT10), .B1(new_n555), .B2(G92), .ZN(new_n602));
  AND4_X1   g177(.A1(KEYINPUT10), .A2(new_n494), .A3(new_n512), .A4(G92), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n504), .A2(KEYINPUT75), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT75), .ZN(new_n607));
  OAI211_X1 g182(.A(new_n607), .B(G543), .C1(new_n500), .C2(new_n501), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n606), .A2(G54), .A3(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(G66), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(new_n492), .B2(new_n493), .ZN(new_n611));
  AND2_X1   g186(.A1(G79), .A2(G543), .ZN(new_n612));
  OAI21_X1  g187(.A(G651), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AND3_X1   g188(.A1(new_n609), .A2(KEYINPUT76), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g189(.A(KEYINPUT76), .B1(new_n609), .B2(new_n613), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n605), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n601), .B1(G868), .B2(new_n617), .ZN(G284));
  OAI21_X1  g193(.A(new_n601), .B1(G868), .B2(new_n617), .ZN(G321));
  NAND2_X1  g194(.A1(G299), .A2(new_n599), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G168), .B2(new_n599), .ZN(G297));
  OAI21_X1  g196(.A(new_n620), .B1(G168), .B2(new_n599), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n617), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n617), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n558), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g203(.A1(new_n464), .A2(new_n467), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT77), .B(KEYINPUT12), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT78), .B(KEYINPUT13), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n633), .A2(G2100), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(G2100), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n465), .A2(G135), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n481), .A2(G123), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n638));
  INV_X1    g213(.A(G111), .ZN(new_n639));
  AOI22_X1  g214(.A1(new_n638), .A2(KEYINPUT79), .B1(new_n639), .B2(G2105), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(KEYINPUT79), .B2(new_n638), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n636), .A2(new_n637), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2096), .Z(new_n643));
  NAND3_X1  g218(.A1(new_n634), .A2(new_n635), .A3(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT80), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2427), .B(G2430), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(KEYINPUT14), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT81), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(G1341), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G1348), .ZN(new_n654));
  XOR2_X1   g229(.A(G2451), .B(G2454), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n656), .B(new_n657), .Z(new_n658));
  NAND2_X1  g233(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(G14), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n654), .A2(new_n658), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(G401));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT17), .Z(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n664), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT82), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n664), .A2(new_n665), .ZN(new_n670));
  INV_X1    g245(.A(new_n663), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n670), .B(new_n667), .C1(new_n671), .C2(new_n665), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n671), .A2(new_n665), .A3(new_n666), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT18), .Z(new_n674));
  NAND3_X1  g249(.A1(new_n669), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2096), .B(G2100), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G227));
  XOR2_X1   g252(.A(G1971), .B(G1976), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT20), .Z(new_n684));
  NOR2_X1   g259(.A1(new_n680), .A2(new_n681), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n679), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT83), .ZN(new_n687));
  NOR3_X1   g262(.A1(new_n679), .A2(new_n682), .A3(new_n685), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n684), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1981), .B(G1986), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT84), .B(KEYINPUT85), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(G229));
  NAND3_X1  g273(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT25), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n471), .A2(G127), .ZN(new_n701));
  NAND2_X1  g276(.A1(G115), .A2(G2104), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n466), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AOI211_X1 g278(.A(new_n700), .B(new_n703), .C1(G139), .C2(new_n465), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT90), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(new_n706), .B2(G33), .ZN(new_n708));
  INV_X1    g283(.A(G2072), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(G160), .A2(G29), .ZN(new_n711));
  INV_X1    g286(.A(G34), .ZN(new_n712));
  AOI21_X1  g287(.A(G29), .B1(new_n712), .B2(KEYINPUT24), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(KEYINPUT24), .B2(new_n712), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n711), .A2(G2084), .A3(new_n714), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n710), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT27), .B(G1996), .Z(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT91), .B(KEYINPUT26), .ZN(new_n718));
  NAND3_X1  g293(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G105), .B2(new_n468), .ZN(new_n721));
  AOI22_X1  g296(.A1(G129), .A2(new_n481), .B1(new_n465), .B2(G141), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT92), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G29), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT93), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n725), .B(new_n726), .C1(G29), .C2(G32), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n726), .B2(new_n725), .ZN(new_n728));
  OAI221_X1 g303(.A(new_n716), .B1(new_n709), .B2(new_n708), .C1(new_n717), .C2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT94), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(G164), .A2(new_n706), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G27), .B2(new_n706), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT96), .B(G2078), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(G5), .A2(G16), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G171), .B2(G16), .ZN(new_n737));
  INV_X1    g312(.A(G1961), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n642), .A2(new_n706), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT30), .B(G28), .ZN(new_n741));
  OR2_X1    g316(.A1(KEYINPUT31), .A2(G11), .ZN(new_n742));
  NAND2_X1  g317(.A1(KEYINPUT31), .A2(G11), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n741), .A2(new_n706), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n735), .A2(new_n739), .A3(new_n740), .A4(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(G2084), .B1(new_n711), .B2(new_n714), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT95), .Z(new_n747));
  INV_X1    g322(.A(G1966), .ZN(new_n748));
  INV_X1    g323(.A(G16), .ZN(new_n749));
  NOR2_X1   g324(.A1(G168), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n749), .B2(G21), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n747), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  OAI221_X1 g327(.A(new_n752), .B1(new_n748), .B2(new_n751), .C1(new_n733), .C2(new_n734), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n745), .B(new_n753), .C1(new_n717), .C2(new_n728), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n731), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n730), .B2(new_n729), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(KEYINPUT97), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(KEYINPUT97), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n749), .A2(KEYINPUT86), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n749), .A2(KEYINPUT86), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(G22), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G166), .B2(new_n761), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G1971), .ZN(new_n764));
  INV_X1    g339(.A(G288), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n765), .A2(new_n749), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n749), .B2(G23), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT33), .B(G1976), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G6), .A2(G16), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n590), .B2(G16), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT32), .B(G1981), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  AOI211_X1 g349(.A(new_n764), .B(new_n774), .C1(new_n767), .C2(new_n768), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT34), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n465), .A2(G131), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n481), .A2(G119), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n466), .A2(G107), .ZN(new_n781));
  OAI21_X1  g356(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n779), .B(new_n780), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  MUX2_X1   g358(.A(G25), .B(new_n783), .S(G29), .Z(new_n784));
  XOR2_X1   g359(.A(KEYINPUT35), .B(G1991), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n761), .A2(G24), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n597), .B(KEYINPUT87), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(new_n761), .ZN(new_n789));
  INV_X1    g364(.A(G1986), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n777), .A2(new_n778), .A3(new_n786), .A4(new_n791), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT36), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n761), .A2(G19), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n558), .B2(new_n761), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(G1341), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n706), .A2(G35), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G162), .B2(new_n706), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT29), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G2090), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n759), .A2(G20), .A3(new_n760), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT23), .ZN(new_n802));
  INV_X1    g377(.A(G299), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(new_n749), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1956), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n706), .A2(G26), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT89), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT28), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n465), .A2(G140), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n481), .A2(G128), .ZN(new_n810));
  OR2_X1    g385(.A1(G104), .A2(G2105), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n811), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n809), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n808), .B1(new_n814), .B2(new_n706), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G2067), .ZN(new_n816));
  NOR3_X1   g391(.A1(new_n800), .A2(new_n805), .A3(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(G4), .A2(G16), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(new_n617), .B2(G16), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT88), .B(G1348), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  AND4_X1   g396(.A1(new_n793), .A2(new_n796), .A3(new_n817), .A4(new_n821), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n757), .A2(new_n758), .A3(new_n822), .ZN(G150));
  INV_X1    g398(.A(G150), .ZN(G311));
  NOR2_X1   g399(.A1(new_n616), .A2(new_n623), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT38), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n494), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n827), .A2(new_n496), .ZN(new_n828));
  INV_X1    g403(.A(G93), .ZN(new_n829));
  INV_X1    g404(.A(G55), .ZN(new_n830));
  OAI22_X1  g405(.A1(new_n502), .A2(new_n829), .B1(new_n504), .B2(new_n830), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n557), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n828), .A2(new_n831), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n834), .A2(new_n554), .A3(new_n556), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n826), .B(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n838));
  INV_X1    g413(.A(G860), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n834), .A2(new_n839), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT37), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(G145));
  XNOR2_X1  g419(.A(new_n724), .B(new_n813), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(G164), .ZN(new_n846));
  INV_X1    g421(.A(new_n705), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(KEYINPUT98), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n847), .A2(KEYINPUT98), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n846), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n481), .A2(G130), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n466), .A2(G118), .ZN(new_n853));
  OAI21_X1  g428(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(G142), .B2(new_n465), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n783), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n631), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n851), .B(new_n860), .C1(new_n846), .C2(new_n849), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n858), .A2(new_n859), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(new_n863), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(G162), .B(G160), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n642), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(G37), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n864), .A2(new_n868), .A3(new_n865), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g449(.A(new_n836), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n625), .B(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n609), .A2(new_n613), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT76), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n609), .A2(KEYINPUT76), .A3(new_n613), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n803), .B1(new_n881), .B2(new_n605), .ZN(new_n882));
  AOI211_X1 g457(.A(new_n604), .B(G299), .C1(new_n879), .C2(new_n880), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n876), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT100), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n616), .A2(G299), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n803), .B(new_n605), .C1(new_n614), .C2(new_n615), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n886), .B1(new_n889), .B2(KEYINPUT41), .ZN(new_n890));
  OAI21_X1  g465(.A(KEYINPUT41), .B1(new_n882), .B2(new_n883), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n887), .A2(new_n892), .A3(new_n888), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n890), .B1(new_n894), .B2(new_n886), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n885), .B1(new_n876), .B2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT42), .ZN(new_n897));
  XNOR2_X1  g472(.A(G288), .B(new_n590), .ZN(new_n898));
  XOR2_X1   g473(.A(G166), .B(new_n597), .Z(new_n899));
  XNOR2_X1  g474(.A(new_n898), .B(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n599), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(new_n900), .B2(new_n897), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT101), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT101), .B1(new_n832), .B2(new_n599), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n904), .B1(new_n902), .B2(new_n905), .ZN(G295));
  AOI21_X1  g481(.A(new_n904), .B1(new_n902), .B2(new_n905), .ZN(G331));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n537), .A2(new_n909), .A3(new_n545), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n909), .B1(new_n537), .B2(new_n545), .ZN(new_n911));
  OAI21_X1  g486(.A(G286), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI22_X1  g487(.A1(new_n555), .A2(new_n543), .B1(new_n524), .B2(G52), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n542), .B1(new_n913), .B2(new_n541), .ZN(new_n914));
  NOR3_X1   g489(.A1(new_n533), .A2(new_n536), .A3(KEYINPUT70), .ZN(new_n915));
  OAI21_X1  g490(.A(KEYINPUT102), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n537), .A2(new_n545), .A3(new_n909), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(G168), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n912), .A2(new_n918), .A3(new_n836), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n836), .B1(new_n912), .B2(new_n918), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n894), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT103), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n919), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n912), .A2(new_n918), .A3(new_n836), .A4(KEYINPUT103), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n921), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n884), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n922), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n900), .ZN(new_n931));
  AOI21_X1  g506(.A(G37), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n921), .B1(new_n924), .B2(new_n925), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT104), .B1(new_n895), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n926), .A2(new_n928), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n887), .A2(new_n892), .A3(new_n888), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n892), .B1(new_n887), .B2(new_n888), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n886), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT100), .B1(new_n884), .B2(new_n892), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT104), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n935), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n934), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n929), .A2(new_n920), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  AND4_X1   g520(.A1(KEYINPUT105), .A2(new_n943), .A3(new_n900), .A4(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n944), .B1(new_n934), .B2(new_n942), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT105), .B1(new_n947), .B2(new_n900), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n932), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n908), .B1(new_n949), .B2(KEYINPUT43), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n895), .A2(new_n933), .A3(KEYINPUT104), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n941), .B1(new_n935), .B2(new_n940), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n945), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n951), .B1(new_n954), .B2(new_n931), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n947), .A2(KEYINPUT105), .A3(new_n900), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n958));
  AOI21_X1  g533(.A(G37), .B1(new_n954), .B2(new_n931), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n957), .A2(KEYINPUT106), .A3(new_n958), .A4(new_n959), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n959), .B(new_n958), .C1(new_n946), .C2(new_n948), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT106), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n950), .A2(new_n960), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT107), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n950), .A2(new_n963), .A3(new_n960), .A4(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n957), .A2(KEYINPUT43), .A3(new_n959), .ZN(new_n969));
  INV_X1    g544(.A(new_n949), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n969), .B1(new_n970), .B2(KEYINPUT43), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n908), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n968), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n968), .A2(new_n973), .A3(KEYINPUT108), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(G397));
  XNOR2_X1  g553(.A(KEYINPUT109), .B(G1384), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT45), .B1(new_n490), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G160), .ZN(new_n981));
  XOR2_X1   g556(.A(KEYINPUT110), .B(G40), .Z(new_n982));
  NOR2_X1   g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G1996), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(KEYINPUT111), .ZN(new_n987));
  OR2_X1    g562(.A1(new_n987), .A2(KEYINPUT46), .ZN(new_n988));
  XOR2_X1   g563(.A(new_n813), .B(G2067), .Z(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT112), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n724), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n984), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n987), .A2(KEYINPUT46), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n988), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT47), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT127), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n996), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n992), .B1(new_n985), .B2(new_n990), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n999), .B1(new_n987), .B2(new_n724), .ZN(new_n1000));
  INV_X1    g575(.A(new_n785), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n783), .B(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1002), .B(KEYINPUT113), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n984), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(G290), .A2(G1986), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n984), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1006), .B(KEYINPUT48), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1000), .A2(new_n1004), .A3(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n783), .A2(new_n1001), .ZN(new_n1009));
  XOR2_X1   g584(.A(new_n1009), .B(KEYINPUT126), .Z(new_n1010));
  NAND2_X1  g585(.A1(new_n1000), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1011), .B1(G2067), .B2(new_n813), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(new_n984), .ZN(new_n1013));
  AND4_X1   g588(.A1(new_n997), .A2(new_n998), .A3(new_n1008), .A4(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G8), .ZN(new_n1015));
  AOI21_X1  g590(.A(G1384), .B1(new_n487), .B2(new_n489), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1015), .B1(new_n1016), .B2(new_n983), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n765), .A2(G1976), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT52), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n590), .B(G1981), .ZN(new_n1021));
  NOR2_X1   g596(.A1(KEYINPUT116), .A2(KEYINPUT49), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1017), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(new_n765), .B2(G1976), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1020), .B(new_n1024), .C1(new_n1019), .C2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n983), .ZN(new_n1028));
  INV_X1    g603(.A(G1384), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n490), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1028), .B1(new_n1030), .B2(KEYINPUT50), .ZN(new_n1031));
  INV_X1    g606(.A(G2090), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT50), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1016), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1031), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1971), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n490), .A2(KEYINPUT45), .A3(new_n979), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n983), .B1(new_n1016), .B2(KEYINPUT45), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1036), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1015), .B1(new_n1035), .B2(new_n1040), .ZN(new_n1041));
  OAI211_X1 g616(.A(G303), .B(G8), .C1(KEYINPUT115), .C2(KEYINPUT55), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1043), .B1(G166), .B2(new_n1015), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1027), .B1(new_n1041), .B2(new_n1046), .ZN(new_n1047));
  OR2_X1    g622(.A1(new_n1041), .A2(new_n1046), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT45), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1030), .A2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1051), .A2(new_n1039), .ZN(new_n1052));
  INV_X1    g627(.A(G2078), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1052), .A2(KEYINPUT53), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n738), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1038), .A2(new_n1039), .A3(G2078), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1054), .B(new_n1056), .C1(new_n1057), .C2(KEYINPUT53), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1058), .A2(KEYINPUT121), .A3(G171), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(G171), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT121), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1049), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G2084), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1031), .A2(new_n1064), .A3(new_n1034), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n748), .B1(new_n1051), .B2(new_n1039), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(G8), .B1(new_n1067), .B2(G286), .ZN(new_n1068));
  OR2_X1    g643(.A1(new_n1068), .A2(KEYINPUT51), .ZN(new_n1069));
  AOI21_X1  g644(.A(G168), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT51), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1069), .A2(KEYINPUT62), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT62), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1063), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI211_X1 g649(.A(G1976), .B(G288), .C1(new_n1017), .C2(new_n1023), .ZN(new_n1075));
  NOR2_X1   g650(.A1(G305), .A2(G1981), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1017), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1041), .A2(new_n1046), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1077), .B1(new_n1078), .B2(new_n1027), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT63), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1067), .A2(G8), .A3(G168), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1080), .B1(new_n1049), .B2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1081), .A2(new_n1080), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1041), .A2(KEYINPUT117), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1045), .B1(new_n1041), .B2(KEYINPUT117), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1047), .B(new_n1083), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1079), .B1(new_n1082), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1074), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G1956), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1055), .A2(new_n1090), .ZN(new_n1091));
  XOR2_X1   g666(.A(G299), .B(KEYINPUT57), .Z(new_n1092));
  NAND2_X1  g667(.A1(new_n1030), .A2(new_n1050), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT56), .B(G2072), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1093), .A2(new_n983), .A3(new_n1037), .A4(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1091), .A2(new_n1092), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1092), .B1(new_n1091), .B2(new_n1095), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT61), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1091), .A2(new_n1095), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1092), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT61), .B1(new_n1103), .B2(new_n1096), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1100), .A2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1093), .A2(new_n985), .A3(new_n983), .A4(new_n1037), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1016), .A2(new_n983), .ZN(new_n1107));
  XOR2_X1   g682(.A(KEYINPUT58), .B(G1341), .Z(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT118), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n558), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT59), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1116), .B(new_n558), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G1348), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1034), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n983), .B1(new_n1016), .B2(new_n1033), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1119), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1107), .A2(G2067), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT60), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT119), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1125), .A2(new_n1126), .A3(new_n616), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1123), .B1(new_n1055), .B2(new_n1119), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1126), .B1(new_n1125), .B2(new_n616), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1128), .A2(KEYINPUT60), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(KEYINPUT60), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1130), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1132), .B1(new_n1133), .B2(new_n1127), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1105), .A2(new_n1118), .A3(new_n1131), .A4(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1129), .A2(new_n616), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1096), .B1(new_n1136), .B2(new_n1098), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1057), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT53), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1139), .A2(new_n1140), .B1(new_n1055), .B2(new_n738), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1141), .A2(G301), .A3(new_n1054), .ZN(new_n1142));
  NAND4_X1  g717(.A1(G160), .A2(KEYINPUT53), .A3(G40), .A4(new_n1053), .ZN(new_n1143));
  OR3_X1    g718(.A1(new_n1038), .A2(new_n980), .A3(new_n1143), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1056), .B(new_n1144), .C1(new_n1057), .C2(KEYINPUT53), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1145), .A2(new_n1146), .A3(G171), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1146), .B1(new_n1145), .B2(G171), .ZN(new_n1148));
  OAI211_X1 g723(.A(KEYINPUT54), .B(new_n1142), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1049), .B1(new_n1071), .B2(new_n1069), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1138), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1141), .A2(KEYINPUT122), .A3(G301), .A4(new_n1144), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT122), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1153), .B1(new_n1145), .B2(G171), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1062), .A2(new_n1152), .A3(new_n1059), .A4(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT123), .ZN(new_n1156));
  XNOR2_X1  g731(.A(KEYINPUT120), .B(KEYINPUT54), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1156), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1089), .B1(new_n1151), .B2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n597), .A2(new_n790), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n984), .B1(new_n1005), .B2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1000), .A2(new_n1004), .A3(new_n1164), .ZN(new_n1165));
  XOR2_X1   g740(.A(new_n1165), .B(KEYINPUT114), .Z(new_n1166));
  INV_X1    g741(.A(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(KEYINPUT125), .B1(new_n1162), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(KEYINPUT123), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n1158), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1049), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1149), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1174), .B1(new_n1137), .B2(new_n1135), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1088), .B1(new_n1171), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT125), .ZN(new_n1177));
  NOR3_X1   g752(.A1(new_n1176), .A2(new_n1177), .A3(new_n1166), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1014), .B1(new_n1168), .B2(new_n1178), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g754(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1181));
  AND3_X1   g755(.A1(new_n873), .A2(new_n697), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g756(.A1(new_n1182), .A2(new_n972), .ZN(G225));
  INV_X1    g757(.A(G225), .ZN(G308));
endmodule


