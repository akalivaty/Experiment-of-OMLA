//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 0 1 1 0 1 1 1 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G116), .ZN(new_n188));
  INV_X1    g002(.A(G116), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT2), .B(G113), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(new_n192), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(KEYINPUT67), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT67), .ZN(new_n197));
  INV_X1    g011(.A(new_n195), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(new_n193), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n196), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  AND2_X1   g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT64), .ZN(new_n208));
  XNOR2_X1  g022(.A(G143), .B(G146), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(new_n206), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n203), .A2(new_n205), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT0), .A2(G128), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n206), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g028(.A1(new_n208), .A2(new_n211), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G131), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT11), .ZN(new_n217));
  INV_X1    g031(.A(G134), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n217), .B1(new_n218), .B2(G137), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(G137), .ZN(new_n220));
  INV_X1    g034(.A(G137), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(KEYINPUT11), .A3(G134), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT66), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n219), .A2(new_n222), .A3(new_n225), .A4(new_n220), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n216), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  XOR2_X1   g041(.A(KEYINPUT65), .B(G131), .Z(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(new_n223), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n215), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT30), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n221), .A2(G134), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n216), .B1(new_n220), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n223), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n234), .B1(new_n235), .B2(new_n228), .ZN(new_n236));
  INV_X1    g050(.A(G128), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n202), .A2(G143), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n212), .A2(new_n237), .B1(KEYINPUT1), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT1), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n203), .A2(new_n205), .A3(new_n240), .A4(G128), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n236), .A2(new_n242), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n231), .A2(new_n232), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n238), .A2(KEYINPUT1), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n245), .B1(new_n209), .B2(G128), .ZN(new_n246));
  AND4_X1   g060(.A1(new_n240), .A2(new_n203), .A3(new_n205), .A4(G128), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT68), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n212), .A2(new_n237), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n249), .A2(new_n250), .A3(new_n241), .A4(new_n245), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n248), .A2(new_n236), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n232), .B1(new_n231), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n201), .B1(new_n244), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n231), .A2(new_n200), .A3(new_n252), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G237), .ZN(new_n257));
  INV_X1    g071(.A(G953), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n258), .A3(G210), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n259), .B(KEYINPUT27), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT26), .B(G101), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n260), .B(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n256), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT29), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT28), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n231), .A2(new_n243), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n201), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n266), .B1(new_n268), .B2(new_n255), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n255), .A2(new_n266), .ZN(new_n270));
  OR2_X1    g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n264), .B(new_n265), .C1(new_n271), .C2(new_n263), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n208), .A2(new_n211), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n212), .A2(new_n214), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT11), .B1(new_n221), .B2(G134), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n221), .A2(G134), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n225), .B1(new_n278), .B2(new_n222), .ZN(new_n279));
  INV_X1    g093(.A(new_n226), .ZN(new_n280));
  OAI21_X1  g094(.A(G131), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n230), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n275), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n248), .A2(new_n236), .A3(new_n251), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n201), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n255), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n270), .B1(new_n286), .B2(KEYINPUT28), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n263), .A2(new_n265), .ZN(new_n288));
  AOI21_X1  g102(.A(G902), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n272), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G472), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT32), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n263), .B1(new_n269), .B2(new_n270), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT30), .B1(new_n283), .B2(new_n284), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n231), .A2(new_n232), .A3(new_n243), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n200), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT31), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n255), .A2(new_n262), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n298), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT31), .B1(new_n254), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n293), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT69), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n297), .B1(new_n296), .B2(new_n298), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n254), .A2(KEYINPUT31), .A3(new_n300), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(KEYINPUT69), .A3(new_n293), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(G472), .A2(G902), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n292), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n310), .ZN(new_n312));
  AOI211_X1 g126(.A(KEYINPUT32), .B(new_n312), .C1(new_n304), .C2(new_n308), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n291), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT70), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(G234), .A2(G237), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(G952), .A3(new_n258), .ZN(new_n318));
  XOR2_X1   g132(.A(KEYINPUT21), .B(G898), .Z(new_n319));
  NAND3_X1  g133(.A1(new_n317), .A2(G902), .A3(G953), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(G214), .B1(G237), .B2(G902), .ZN(new_n322));
  XNOR2_X1  g136(.A(G110), .B(G122), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n323), .B(KEYINPUT82), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n325));
  XNOR2_X1  g139(.A(G104), .B(G107), .ZN(new_n326));
  INV_X1    g140(.A(G101), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G107), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G104), .ZN(new_n330));
  INV_X1    g144(.A(G104), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G107), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(KEYINPUT77), .A3(G101), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n328), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT3), .B1(new_n331), .B2(G107), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT3), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(new_n329), .A3(G104), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n336), .A2(new_n338), .A3(new_n327), .A4(new_n332), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT76), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n339), .A2(new_n340), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n335), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n336), .A2(new_n332), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n346), .A2(KEYINPUT76), .A3(new_n327), .A4(new_n338), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n339), .A2(new_n340), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(KEYINPUT79), .A3(new_n335), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT5), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n188), .A2(KEYINPUT5), .ZN(new_n352));
  INV_X1    g166(.A(G113), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n193), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n345), .A2(new_n350), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT81), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n345), .A2(new_n350), .A3(KEYINPUT81), .A4(new_n355), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n336), .A2(new_n338), .A3(new_n332), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT4), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n361), .A3(G101), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n361), .B1(new_n360), .B2(G101), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n363), .B1(new_n349), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n201), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n359), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n324), .B1(new_n358), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n356), .A2(new_n357), .ZN(new_n369));
  INV_X1    g183(.A(new_n324), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n369), .A2(new_n370), .A3(new_n359), .A4(new_n366), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(KEYINPUT6), .A3(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n246), .A2(new_n247), .ZN(new_n373));
  INV_X1    g187(.A(G125), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n376), .B1(G125), .B2(new_n275), .ZN(new_n377));
  INV_X1    g191(.A(G224), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n378), .A2(G953), .ZN(new_n379));
  XOR2_X1   g193(.A(new_n377), .B(new_n379), .Z(new_n380));
  INV_X1    g194(.A(KEYINPUT6), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n381), .B(new_n324), .C1(new_n358), .C2(new_n367), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n372), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n375), .A2(KEYINPUT84), .B1(new_n275), .B2(G125), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n384), .B1(KEYINPUT84), .B2(new_n375), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT7), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n385), .B1(new_n386), .B2(new_n379), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n377), .B(KEYINPUT7), .C1(new_n378), .C2(G953), .ZN(new_n388));
  AOI22_X1  g202(.A1(new_n347), .A2(new_n348), .B1(new_n328), .B2(new_n334), .ZN(new_n389));
  OR2_X1    g203(.A1(new_n354), .A2(KEYINPUT83), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n354), .A2(KEYINPUT83), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n390), .A2(new_n351), .A3(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n389), .B1(new_n392), .B2(new_n193), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n343), .A2(new_n355), .ZN(new_n394));
  XOR2_X1   g208(.A(new_n324), .B(KEYINPUT8), .Z(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n387), .A2(new_n388), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(G902), .B1(new_n397), .B2(new_n371), .ZN(new_n398));
  OAI21_X1  g212(.A(G210), .B1(G237), .B2(G902), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n383), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n399), .B1(new_n383), .B2(new_n398), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n321), .B(new_n322), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT9), .B(G234), .ZN(new_n403));
  OAI21_X1  g217(.A(G221), .B1(new_n403), .B2(G902), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n227), .A2(new_n230), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n248), .A2(KEYINPUT10), .A3(new_n251), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n345), .A2(new_n350), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n241), .A2(KEYINPUT78), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT78), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n209), .A2(new_n411), .A3(new_n240), .A4(G128), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n239), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n349), .A2(new_n335), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT10), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n349), .A2(new_n364), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(new_n215), .A3(new_n362), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n406), .B1(new_n409), .B2(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(G110), .B(G140), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n258), .A2(G227), .ZN(new_n422));
  XOR2_X1   g236(.A(new_n421), .B(new_n422), .Z(new_n423));
  AOI22_X1  g237(.A1(new_n365), .A2(new_n215), .B1(new_n414), .B2(new_n415), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(new_n405), .A3(new_n408), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n420), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n424), .A2(new_n405), .A3(new_n408), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT80), .B1(new_n389), .B2(new_n242), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT80), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n343), .A2(new_n429), .A3(new_n373), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(new_n430), .A3(new_n414), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n406), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT12), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n431), .A2(KEYINPUT12), .A3(new_n406), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n427), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI211_X1 g250(.A(G469), .B(new_n426), .C1(new_n436), .C2(new_n423), .ZN(new_n437));
  NAND2_X1  g251(.A1(G469), .A2(G902), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n431), .A2(KEYINPUT12), .A3(new_n406), .ZN(new_n440));
  AOI21_X1  g254(.A(KEYINPUT12), .B1(new_n431), .B2(new_n406), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n423), .B(new_n425), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n423), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n405), .B1(new_n424), .B2(new_n408), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n443), .B1(new_n427), .B2(new_n444), .ZN(new_n445));
  AOI211_X1 g259(.A(G469), .B(G902), .C1(new_n442), .C2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n404), .B1(new_n439), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n257), .A2(new_n258), .A3(G214), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n448), .B(new_n204), .ZN(new_n449));
  NAND2_X1  g263(.A1(KEYINPUT18), .A2(G131), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n449), .B(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G125), .B(G140), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT71), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G140), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(KEYINPUT71), .A3(G125), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(KEYINPUT85), .B1(new_n458), .B2(G146), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n454), .A2(KEYINPUT85), .A3(G146), .A4(new_n456), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n452), .B(KEYINPUT73), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n460), .B1(new_n461), .B2(G146), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n451), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n449), .B(new_n229), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n454), .A2(KEYINPUT16), .A3(new_n456), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT16), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(new_n374), .B2(G140), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(G146), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT19), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n461), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n457), .A2(KEYINPUT19), .ZN(new_n473));
  AOI21_X1  g287(.A(G146), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n463), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(G113), .B(G122), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT86), .B(G104), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n476), .B(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n478), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n449), .A2(KEYINPUT17), .A3(new_n229), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n481), .B1(new_n464), .B2(KEYINPUT17), .ZN(new_n482));
  OAI21_X1  g296(.A(KEYINPUT72), .B1(new_n468), .B2(G146), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT72), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n465), .A2(new_n484), .A3(new_n202), .A4(new_n467), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(new_n485), .A3(new_n469), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n463), .B(new_n480), .C1(new_n482), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n479), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT20), .ZN(new_n489));
  INV_X1    g303(.A(G475), .ZN(new_n490));
  INV_X1    g304(.A(G902), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(KEYINPUT87), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n488), .A2(new_n489), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n489), .B1(new_n488), .B2(new_n493), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n463), .B1(new_n482), .B2(new_n486), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n478), .ZN(new_n498));
  AOI21_X1  g312(.A(G902), .B1(new_n498), .B2(new_n487), .ZN(new_n499));
  OAI22_X1  g313(.A1(new_n495), .A2(new_n496), .B1(new_n490), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n189), .A2(G122), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n189), .A2(G122), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(new_n504), .A3(new_n329), .ZN(new_n505));
  OR2_X1    g319(.A1(new_n505), .A2(KEYINPUT89), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(KEYINPUT89), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n204), .A2(G128), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n237), .A2(G143), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n218), .ZN(new_n511));
  INV_X1    g325(.A(new_n510), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G134), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n506), .A2(new_n507), .A3(new_n511), .A4(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n504), .ZN(new_n515));
  INV_X1    g329(.A(G122), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT14), .B1(new_n516), .B2(G116), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT90), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n504), .A2(KEYINPUT14), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT90), .ZN(new_n521));
  NOR3_X1   g335(.A1(new_n504), .A2(new_n521), .A3(KEYINPUT14), .ZN(new_n522));
  OAI211_X1 g336(.A(KEYINPUT91), .B(G107), .C1(new_n520), .C2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT91), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n522), .B1(new_n518), .B2(new_n519), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n524), .B1(new_n525), .B2(new_n329), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n514), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT13), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n218), .B1(new_n509), .B2(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n512), .B(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n515), .A2(new_n502), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(new_n329), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT88), .ZN(new_n535));
  INV_X1    g349(.A(new_n505), .ZN(new_n536));
  OR3_X1    g350(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n535), .B1(new_n534), .B2(new_n536), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n532), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(G217), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n403), .A2(new_n541), .A3(G953), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n528), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n542), .B1(new_n527), .B2(new_n539), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n544), .A2(KEYINPUT92), .A3(new_n545), .A4(new_n491), .ZN(new_n546));
  INV_X1    g360(.A(G478), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n547), .A2(KEYINPUT15), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n546), .B(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n501), .A2(new_n550), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n402), .A2(new_n447), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n541), .B1(G234), .B2(new_n491), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT22), .B(G137), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n258), .A2(G221), .A3(G234), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n555), .B(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n237), .A2(G119), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n187), .A2(G128), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT24), .B(G110), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT23), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n237), .A2(KEYINPUT23), .A3(G119), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n566), .A3(new_n560), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n563), .B1(G110), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n486), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n561), .A2(new_n562), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n570), .B1(new_n567), .B2(G110), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n469), .B(new_n571), .C1(G146), .C2(new_n461), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n558), .B1(new_n569), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n569), .A2(new_n572), .A3(new_n558), .ZN(new_n575));
  AOI21_X1  g389(.A(G902), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT25), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n554), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n575), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n491), .B1(new_n579), .B2(new_n573), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT25), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n553), .A2(G902), .ZN(new_n582));
  XOR2_X1   g396(.A(new_n582), .B(KEYINPUT74), .Z(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n584), .B1(new_n579), .B2(new_n573), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT75), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g401(.A(KEYINPUT75), .B(new_n584), .C1(new_n579), .C2(new_n573), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n578), .A2(new_n581), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI211_X1 g403(.A(KEYINPUT70), .B(new_n291), .C1(new_n311), .C2(new_n313), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n316), .A2(new_n552), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(KEYINPUT93), .B(G101), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n591), .B(new_n592), .ZN(G3));
  INV_X1    g407(.A(new_n308), .ZN(new_n594));
  AOI21_X1  g408(.A(KEYINPUT69), .B1(new_n307), .B2(new_n293), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n491), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT94), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n597), .A3(G472), .ZN(new_n598));
  AOI21_X1  g412(.A(G902), .B1(new_n304), .B2(new_n308), .ZN(new_n599));
  INV_X1    g413(.A(G472), .ZN(new_n600));
  OAI21_X1  g414(.A(KEYINPUT94), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n309), .A2(new_n310), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n598), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT95), .ZN(new_n604));
  INV_X1    g418(.A(new_n589), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n447), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n606), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n598), .A2(new_n601), .A3(new_n602), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT95), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT96), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n528), .B(new_n540), .C1(KEYINPUT98), .C2(new_n542), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n542), .A2(KEYINPUT98), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n614), .B1(new_n527), .B2(new_n539), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n613), .A2(KEYINPUT33), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT97), .B(KEYINPUT33), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n544), .A2(new_n545), .A3(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n616), .A2(G478), .A3(new_n618), .A4(new_n491), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n544), .A2(new_n491), .A3(new_n545), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n547), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n500), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(new_n623), .B(KEYINPUT99), .Z(new_n624));
  INV_X1    g438(.A(new_n402), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n612), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT100), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT34), .B(G104), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  NAND2_X1  g445(.A1(new_n501), .A2(new_n549), .ZN(new_n632));
  OR2_X1    g446(.A1(new_n402), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n612), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT35), .B(G107), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G9));
  AND2_X1   g451(.A1(new_n569), .A2(new_n572), .ZN(new_n638));
  OR2_X1    g452(.A1(new_n558), .A2(KEYINPUT36), .ZN(new_n639));
  XOR2_X1   g453(.A(new_n639), .B(KEYINPUT101), .Z(new_n640));
  OR2_X1    g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n640), .A2(new_n569), .A3(new_n572), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI22_X1  g457(.A1(new_n578), .A2(new_n581), .B1(new_n584), .B2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n603), .A2(new_n552), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT37), .B(G110), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT102), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT103), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n646), .B(new_n649), .ZN(G12));
  INV_X1    g464(.A(new_n322), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n383), .A2(new_n398), .ZN(new_n652));
  INV_X1    g466(.A(new_n399), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n383), .A2(new_n398), .A3(new_n399), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n651), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n496), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n494), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n499), .A2(new_n490), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n318), .B1(new_n320), .B2(G900), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n658), .A2(new_n549), .A3(new_n659), .A4(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(new_n644), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n447), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n316), .A2(new_n664), .A3(new_n590), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G128), .ZN(G30));
  XNOR2_X1  g481(.A(new_n660), .B(KEYINPUT39), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(new_n669), .B(KEYINPUT40), .Z(new_n670));
  NAND2_X1  g484(.A1(new_n654), .A2(new_n655), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT38), .ZN(new_n672));
  AOI22_X1  g486(.A1(new_n254), .A2(new_n300), .B1(new_n286), .B2(new_n263), .ZN(new_n673));
  OAI21_X1  g487(.A(G472), .B1(new_n673), .B2(G902), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n674), .B1(new_n311), .B2(new_n313), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n501), .A2(new_n550), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n676), .A2(new_n322), .A3(new_n644), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT104), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n670), .A2(new_n672), .A3(new_n675), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G143), .ZN(G45));
  NAND3_X1  g494(.A1(new_n500), .A2(new_n622), .A3(new_n660), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n671), .A2(new_n322), .A3(new_n645), .A4(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n684), .A2(new_n316), .A3(new_n590), .A4(new_n665), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G146), .ZN(G48));
  NAND2_X1  g500(.A1(new_n434), .A2(new_n435), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n425), .A2(new_n423), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n420), .A2(new_n425), .ZN(new_n690));
  AOI22_X1  g504(.A1(new_n687), .A2(new_n689), .B1(new_n690), .B2(new_n443), .ZN(new_n691));
  OAI21_X1  g505(.A(G469), .B1(new_n691), .B2(G902), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n442), .A2(new_n445), .ZN(new_n693));
  INV_X1    g507(.A(G469), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n693), .A2(new_n694), .A3(new_n491), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n692), .A2(new_n404), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(KEYINPUT105), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT105), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n692), .A2(new_n695), .A3(new_n698), .A4(new_n404), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n316), .A2(new_n589), .A3(new_n590), .A4(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n627), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT41), .B(G113), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G15));
  NAND2_X1  g519(.A1(new_n702), .A2(new_n634), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G116), .ZN(G18));
  AND2_X1   g521(.A1(new_n316), .A2(new_n590), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n402), .A2(new_n551), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n697), .A2(new_n699), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n711), .A2(new_n644), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n708), .A2(new_n709), .A3(new_n710), .A4(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n712), .A2(new_n316), .A3(new_n590), .A4(new_n710), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(KEYINPUT106), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  NAND3_X1  g531(.A1(new_n697), .A2(new_n676), .A3(new_n699), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n402), .ZN(new_n719));
  XOR2_X1   g533(.A(KEYINPUT107), .B(G472), .Z(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n596), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT108), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n307), .B1(new_n287), .B2(new_n262), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n310), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n722), .A2(new_n723), .A3(new_n589), .A4(new_n725), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n589), .B(new_n725), .C1(new_n599), .C2(new_n720), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(KEYINPUT108), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n719), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G122), .ZN(G24));
  OAI211_X1 g545(.A(new_n645), .B(new_n725), .C1(new_n599), .C2(new_n720), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n681), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(new_n700), .A3(new_n656), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G125), .ZN(G27));
  NAND3_X1  g549(.A1(new_n314), .A2(new_n589), .A3(new_n682), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n654), .A2(new_n322), .A3(new_n655), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n447), .A2(KEYINPUT109), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n695), .A2(new_n437), .A3(new_n438), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n740), .B1(new_n741), .B2(new_n404), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n738), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(KEYINPUT42), .B1(new_n736), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n447), .A2(KEYINPUT109), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n741), .A2(new_n740), .A3(new_n404), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n737), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n316), .A2(new_n747), .A3(new_n589), .A4(new_n590), .ZN(new_n748));
  OR2_X1    g562(.A1(new_n681), .A2(KEYINPUT42), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n744), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(new_n216), .ZN(G33));
  NOR2_X1   g565(.A1(new_n748), .A2(new_n661), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n218), .ZN(G36));
  OAI21_X1  g567(.A(new_n426), .B1(new_n436), .B2(new_n423), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(KEYINPUT45), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(G469), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n756), .A2(KEYINPUT46), .A3(new_n438), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT46), .B1(new_n756), .B2(new_n438), .ZN(new_n758));
  OR3_X1    g572(.A1(new_n757), .A2(new_n758), .A3(new_n446), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n404), .A3(new_n668), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT110), .ZN(new_n761));
  INV_X1    g575(.A(new_n622), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n500), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(KEYINPUT43), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n609), .A3(new_n645), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n738), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n767), .B1(new_n766), .B2(new_n765), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n761), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G137), .ZN(G39));
  INV_X1    g584(.A(new_n708), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n771), .A2(new_n605), .A3(new_n682), .A4(new_n738), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n759), .A2(new_n404), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT47), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n759), .A2(KEYINPUT47), .A3(new_n404), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n772), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(new_n455), .ZN(G42));
  NAND2_X1  g592(.A1(new_n692), .A2(new_n695), .ZN(new_n779));
  XOR2_X1   g593(.A(new_n779), .B(KEYINPUT111), .Z(new_n780));
  XOR2_X1   g594(.A(new_n780), .B(KEYINPUT49), .Z(new_n781));
  NAND4_X1  g595(.A1(new_n763), .A2(new_n589), .A3(new_n404), .A4(new_n322), .ZN(new_n782));
  OR4_X1    g596(.A1(new_n672), .A2(new_n781), .A3(new_n675), .A4(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n730), .A2(new_n591), .A3(new_n646), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n785), .B1(new_n713), .B2(new_n715), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n733), .A2(new_n747), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n501), .A2(new_n550), .A3(new_n660), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n737), .A2(new_n788), .A3(new_n644), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n316), .A2(new_n590), .A3(new_n665), .A4(new_n789), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n787), .B(new_n790), .C1(new_n748), .C2(new_n661), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n750), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n701), .B1(new_n626), .B2(new_n633), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n632), .A2(new_n623), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(new_n402), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n607), .A2(new_n610), .A3(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n665), .A2(new_n644), .A3(new_n660), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n798), .A2(new_n656), .A3(new_n675), .A4(new_n676), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n685), .A2(new_n666), .A3(new_n734), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(KEYINPUT52), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n786), .A2(new_n792), .A3(new_n797), .A4(new_n801), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n666), .A2(new_n734), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT112), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n803), .A2(new_n804), .A3(new_n685), .A4(new_n799), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n800), .A2(KEYINPUT112), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT52), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n784), .B1(new_n802), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n786), .A2(new_n792), .A3(new_n797), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n805), .A2(KEYINPUT52), .A3(new_n806), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n808), .B1(new_n812), .B2(new_n784), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(KEYINPUT54), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n814), .A2(KEYINPUT113), .ZN(new_n815));
  INV_X1    g629(.A(new_n404), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n780), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n775), .A2(new_n776), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n764), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n318), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n820), .A2(new_n729), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n821), .A2(new_n738), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n700), .A2(new_n738), .ZN(new_n824));
  NOR4_X1   g638(.A1(new_n824), .A2(new_n675), .A3(new_n605), .A4(new_n318), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(new_n501), .A3(new_n762), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n820), .A2(new_n700), .A3(new_n738), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n826), .B1(new_n732), .B2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n828), .B(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n672), .A2(new_n322), .A3(new_n711), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n832), .A2(new_n833), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n821), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT50), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n830), .A2(new_n831), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n831), .B1(new_n830), .B2(new_n840), .ZN(new_n842));
  OAI211_X1 g656(.A(KEYINPUT51), .B(new_n823), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n314), .A2(new_n589), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n827), .A2(new_n844), .ZN(new_n845));
  XOR2_X1   g659(.A(new_n845), .B(KEYINPUT48), .Z(new_n846));
  NAND3_X1  g660(.A1(new_n821), .A2(new_n656), .A3(new_n700), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n258), .A2(G952), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n848), .B1(new_n825), .B2(new_n624), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n828), .B1(new_n838), .B2(new_n839), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n775), .A2(KEYINPUT115), .A3(new_n776), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n817), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT115), .B1(new_n775), .B2(new_n776), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n822), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  XOR2_X1   g670(.A(KEYINPUT114), .B(KEYINPUT51), .Z(new_n857));
  AOI21_X1  g671(.A(new_n850), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n843), .A2(new_n858), .ZN(new_n859));
  OR3_X1    g673(.A1(new_n802), .A2(new_n807), .A3(new_n784), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n861));
  INV_X1    g675(.A(new_n811), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n862), .A2(new_n807), .A3(new_n809), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n860), .B(new_n861), .C1(new_n863), .C2(KEYINPUT53), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n864), .B1(new_n814), .B2(KEYINPUT113), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n815), .A2(new_n859), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(G952), .A2(G953), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n783), .B1(new_n866), .B2(new_n867), .ZN(G75));
  OAI21_X1  g682(.A(new_n860), .B1(new_n863), .B2(KEYINPUT53), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n869), .A2(G210), .A3(G902), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT56), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n372), .A2(new_n382), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(new_n380), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT55), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n870), .A2(new_n871), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n874), .B1(new_n870), .B2(new_n871), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n258), .A2(G952), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(G51));
  INV_X1    g692(.A(new_n877), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT53), .B1(new_n810), .B2(new_n811), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n802), .A2(new_n807), .A3(new_n784), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT54), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n864), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n438), .B(KEYINPUT57), .Z(new_n884));
  AOI21_X1  g698(.A(new_n691), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n756), .ZN(new_n886));
  OAI211_X1 g700(.A(G902), .B(new_n886), .C1(new_n880), .C2(new_n881), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT119), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n869), .A2(KEYINPUT119), .A3(G902), .A4(new_n886), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n879), .B1(new_n885), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT120), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT120), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n894), .B(new_n879), .C1(new_n885), .C2(new_n891), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n893), .A2(new_n895), .ZN(G54));
  AND2_X1   g710(.A1(KEYINPUT58), .A2(G475), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n869), .A2(G902), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n898), .A2(new_n479), .A3(new_n487), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n869), .A2(G902), .A3(new_n488), .A4(new_n897), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n899), .A2(new_n879), .A3(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n901), .B(new_n902), .ZN(G60));
  NAND2_X1  g717(.A1(G478), .A2(G902), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT59), .Z(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n883), .A2(new_n616), .A3(new_n618), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n879), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n906), .B1(new_n815), .B2(new_n865), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n616), .A2(new_n618), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(G63));
  NOR2_X1   g725(.A1(new_n880), .A2(new_n881), .ZN(new_n912));
  NAND2_X1  g726(.A1(G217), .A2(G902), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT60), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n643), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n575), .B(new_n574), .C1(new_n912), .C2(new_n914), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n916), .A2(new_n879), .A3(new_n917), .ZN(new_n918));
  XOR2_X1   g732(.A(KEYINPUT122), .B(KEYINPUT61), .Z(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n918), .B(new_n920), .ZN(G66));
  NAND2_X1  g735(.A1(new_n786), .A2(new_n797), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT123), .Z(new_n923));
  NOR2_X1   g737(.A1(new_n378), .A2(new_n258), .ZN(new_n924));
  AOI22_X1  g738(.A1(new_n923), .A2(new_n258), .B1(new_n319), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n872), .B1(G898), .B2(new_n258), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(G69));
  NAND2_X1  g741(.A1(G227), .A2(G900), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n803), .A2(new_n685), .ZN(new_n929));
  NOR4_X1   g743(.A1(new_n777), .A2(new_n750), .A3(new_n752), .A4(new_n929), .ZN(new_n930));
  AND4_X1   g744(.A1(new_n589), .A2(new_n314), .A3(new_n656), .A4(new_n676), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n761), .B1(new_n768), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(G953), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n258), .A2(G900), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT124), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n933), .A2(KEYINPUT124), .A3(new_n934), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n244), .A2(new_n253), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n472), .A2(new_n473), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(new_n942));
  OAI211_X1 g756(.A(G953), .B(new_n928), .C1(new_n939), .C2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n928), .A2(G953), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n771), .A2(new_n605), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n669), .A2(new_n794), .A3(new_n737), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n777), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n769), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n679), .A2(new_n685), .A3(new_n803), .ZN(new_n949));
  OR2_X1    g763(.A1(new_n949), .A2(KEYINPUT62), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(KEYINPUT62), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n942), .B1(new_n952), .B2(G953), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n937), .A2(new_n938), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n944), .B(new_n953), .C1(new_n954), .C2(new_n942), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n943), .A2(new_n955), .ZN(G72));
  XNOR2_X1  g770(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n600), .A2(new_n491), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT126), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n952), .B2(new_n923), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT127), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n262), .B(new_n256), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n963), .B1(new_n962), .B2(new_n961), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n256), .A2(new_n262), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n923), .A2(new_n930), .A3(new_n932), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n965), .B1(new_n966), .B2(new_n960), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n254), .A2(new_n300), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n959), .B1(new_n264), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n813), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n967), .A2(new_n879), .A3(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n964), .A2(new_n971), .ZN(G57));
endmodule


