//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 1 1 1 0 0 0 0 1 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(KEYINPUT64), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n190), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n190), .A2(G146), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n193), .A2(KEYINPUT64), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n191), .A2(G146), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G143), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT68), .A3(KEYINPUT1), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G128), .ZN(new_n203));
  AOI21_X1  g017(.A(KEYINPUT68), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n198), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G125), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n193), .A2(G143), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(KEYINPUT1), .ZN(new_n210));
  AND3_X1   g024(.A1(new_n201), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n205), .A2(new_n206), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT84), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT84), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n205), .A2(new_n215), .A3(new_n206), .A4(new_n212), .ZN(new_n216));
  AND2_X1   g030(.A1(KEYINPUT0), .A2(G128), .ZN(new_n217));
  NOR2_X1   g031(.A1(KEYINPUT0), .A2(G128), .ZN(new_n218));
  OR2_X1    g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n198), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT64), .B(G146), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n207), .B1(new_n222), .B2(G143), .ZN(new_n223));
  AOI21_X1  g037(.A(KEYINPUT65), .B1(new_n223), .B2(new_n217), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n201), .A2(KEYINPUT65), .A3(new_n208), .A4(new_n217), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n221), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G125), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n214), .A2(new_n216), .A3(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT83), .B(G224), .ZN(new_n230));
  OR2_X1    g044(.A1(new_n230), .A2(G953), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT7), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT85), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n205), .A2(new_n206), .A3(new_n212), .ZN(new_n235));
  INV_X1    g049(.A(new_n232), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n219), .B1(new_n195), .B2(new_n197), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n201), .A2(new_n208), .A3(new_n217), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n237), .B1(new_n240), .B2(new_n225), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n236), .B1(new_n241), .B2(new_n206), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n234), .B1(new_n235), .B2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n232), .B1(new_n227), .B2(G125), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(KEYINPUT85), .A3(new_n213), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT86), .ZN(new_n247));
  INV_X1    g061(.A(G113), .ZN(new_n248));
  XOR2_X1   g062(.A(KEYINPUT81), .B(KEYINPUT5), .Z(new_n249));
  INV_X1    g063(.A(G116), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(G119), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n248), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT5), .ZN(new_n253));
  XOR2_X1   g067(.A(G116), .B(G119), .Z(new_n254));
  OAI21_X1  g068(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT2), .B(G113), .ZN(new_n256));
  OR2_X1    g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT77), .B(G101), .ZN(new_n259));
  INV_X1    g073(.A(G107), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G104), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n262));
  INV_X1    g076(.A(G104), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G107), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT3), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(new_n260), .A3(G104), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n259), .A2(new_n262), .A3(new_n264), .A4(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(G104), .B(G107), .ZN(new_n268));
  INV_X1    g082(.A(G101), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT78), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n261), .A2(new_n264), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT78), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(G101), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n267), .A2(new_n270), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n258), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n252), .B1(new_n254), .B2(new_n249), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(new_n257), .A3(new_n274), .ZN(new_n278));
  XNOR2_X1  g092(.A(G110), .B(G122), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n279), .B(KEYINPUT8), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n276), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n233), .A2(new_n246), .A3(new_n247), .A4(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n262), .A2(new_n266), .A3(new_n264), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n267), .A2(KEYINPUT4), .B1(new_n283), .B2(G101), .ZN(new_n284));
  AND3_X1   g098(.A1(new_n283), .A2(KEYINPUT4), .A3(G101), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  XOR2_X1   g100(.A(new_n254), .B(new_n256), .Z(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n275), .A2(new_n277), .A3(new_n257), .ZN(new_n289));
  INV_X1    g103(.A(new_n279), .ZN(new_n290));
  OR3_X1    g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n282), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n281), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n293), .B1(new_n243), .B2(new_n245), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n247), .B1(new_n294), .B2(new_n233), .ZN(new_n295));
  OAI211_X1 g109(.A(KEYINPUT87), .B(new_n189), .C1(new_n292), .C2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n290), .B1(new_n288), .B2(new_n289), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n291), .A2(KEYINPUT82), .A3(KEYINPUT6), .A4(new_n297), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n291), .A2(KEYINPUT6), .A3(new_n297), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT82), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n300), .B1(new_n297), .B2(KEYINPUT6), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n298), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n228), .A2(new_n213), .ZN(new_n303));
  XOR2_X1   g117(.A(new_n303), .B(new_n231), .Z(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n296), .A2(new_n305), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n235), .A2(new_n242), .A3(new_n234), .ZN(new_n307));
  AOI21_X1  g121(.A(KEYINPUT85), .B1(new_n244), .B2(new_n213), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n281), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n213), .A2(KEYINPUT84), .B1(G125), .B2(new_n227), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n236), .B1(new_n310), .B2(new_n216), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT86), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(new_n291), .A3(new_n282), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT87), .B1(new_n313), .B2(new_n189), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n188), .B1(new_n306), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n189), .B1(new_n292), .B2(new_n295), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT87), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n318), .A2(new_n187), .A3(new_n305), .A4(new_n296), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT91), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n322));
  INV_X1    g136(.A(G140), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(new_n323), .A3(G125), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(G125), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n206), .A2(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g141(.A(KEYINPUT16), .B(new_n324), .C1(new_n327), .C2(new_n322), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT16), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G146), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n328), .A2(new_n193), .A3(new_n330), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT17), .ZN(new_n335));
  NOR2_X1   g149(.A1(G237), .A2(G953), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(G143), .A3(G214), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(G143), .B1(new_n336), .B2(G214), .ZN(new_n339));
  OAI21_X1  g153(.A(G131), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT88), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G237), .ZN(new_n343));
  INV_X1    g157(.A(G953), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n344), .A3(G214), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n190), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n337), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(KEYINPUT88), .A3(G131), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n335), .B1(new_n342), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n321), .B1(new_n334), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT88), .B1(new_n347), .B2(G131), .ZN(new_n351));
  INV_X1    g165(.A(G131), .ZN(new_n352));
  AOI211_X1 g166(.A(new_n341), .B(new_n352), .C1(new_n346), .C2(new_n337), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT17), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n354), .A2(KEYINPUT91), .A3(new_n333), .A4(new_n332), .ZN(new_n355));
  INV_X1    g169(.A(new_n347), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n352), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n342), .A2(new_n357), .A3(new_n348), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n335), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n350), .A2(new_n355), .A3(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(G113), .B(G122), .ZN(new_n361));
  XNOR2_X1  g175(.A(KEYINPUT89), .B(G104), .ZN(new_n362));
  XOR2_X1   g176(.A(new_n361), .B(new_n362), .Z(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT18), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n356), .B1(new_n365), .B2(new_n352), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n222), .A2(new_n325), .A3(new_n326), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n324), .B1(new_n327), .B2(new_n322), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n367), .B1(new_n368), .B2(new_n193), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n347), .A2(KEYINPUT18), .A3(G131), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n366), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n360), .A2(new_n364), .A3(new_n371), .ZN(new_n372));
  MUX2_X1   g186(.A(new_n327), .B(new_n368), .S(KEYINPUT19), .Z(new_n373));
  AOI22_X1  g187(.A1(new_n373), .A2(new_n222), .B1(G146), .B2(new_n331), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n342), .A2(new_n357), .A3(new_n348), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n371), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT90), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(new_n363), .ZN(new_n379));
  INV_X1    g193(.A(new_n371), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n380), .B1(new_n374), .B2(new_n375), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT90), .B1(new_n381), .B2(new_n364), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n372), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(G475), .A2(G902), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT20), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT20), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n383), .A2(new_n387), .A3(new_n384), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT96), .B(G952), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n390), .A2(G953), .ZN(new_n391));
  NAND2_X1  g205(.A1(G234), .A2(G237), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT21), .B(G898), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n392), .A2(G902), .A3(G953), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n394), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n372), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n364), .B1(new_n360), .B2(new_n371), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n189), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n398), .B1(new_n401), .B2(G475), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT15), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G478), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT9), .B(G234), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(G217), .A3(new_n344), .ZN(new_n407));
  INV_X1    g221(.A(G122), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT92), .B1(new_n408), .B2(G116), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT92), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n410), .A2(new_n250), .A3(G122), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n408), .A2(G116), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n260), .A3(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(G128), .B(G143), .ZN(new_n415));
  OR2_X1    g229(.A1(new_n415), .A2(G134), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(G134), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n414), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT14), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n409), .A2(new_n411), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT93), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n421), .B1(new_n412), .B2(KEYINPUT14), .ZN(new_n422));
  AOI211_X1 g236(.A(KEYINPUT93), .B(new_n419), .C1(new_n409), .C2(new_n411), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n413), .B(new_n420), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n418), .B1(new_n424), .B2(G107), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n209), .A2(G143), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT13), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n427), .A3(G134), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n416), .A2(new_n417), .A3(new_n428), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n415), .A2(new_n427), .A3(G134), .A4(new_n426), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n414), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n260), .B1(new_n412), .B2(new_n413), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n407), .B1(new_n425), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n418), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n420), .A2(new_n413), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n412), .A2(KEYINPUT14), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT93), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n412), .A2(new_n421), .A3(KEYINPUT14), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n438), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n437), .B1(new_n442), .B2(new_n260), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n429), .B(new_n430), .C1(new_n433), .C2(new_n432), .ZN(new_n444));
  INV_X1    g258(.A(new_n407), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(G902), .B1(new_n436), .B2(new_n446), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(KEYINPUT94), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT94), .ZN(new_n449));
  AOI211_X1 g263(.A(new_n449), .B(G902), .C1(new_n436), .C2(new_n446), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n404), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT95), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n447), .A2(KEYINPUT94), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(new_n403), .A3(G478), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n452), .B1(new_n451), .B2(new_n454), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n389), .B(new_n402), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G221), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n459), .B1(new_n406), .B2(new_n189), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(G110), .B(G140), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n344), .A2(G227), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n462), .B(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT11), .ZN(new_n466));
  INV_X1    g280(.A(G134), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n466), .B1(new_n467), .B2(G137), .ZN(new_n468));
  INV_X1    g282(.A(G137), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(KEYINPUT11), .A3(G134), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n467), .A2(G137), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n468), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G131), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n468), .A2(new_n470), .A3(new_n352), .A4(new_n471), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT10), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT1), .B1(new_n190), .B2(G146), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n201), .A2(new_n208), .B1(G128), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n211), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n476), .B1(new_n479), .B2(new_n274), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n480), .B1(new_n227), .B2(new_n286), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n267), .A2(new_n270), .A3(new_n273), .A4(KEYINPUT10), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n482), .B1(new_n205), .B2(new_n212), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n475), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n205), .A2(new_n212), .ZN(new_n485));
  INV_X1    g299(.A(new_n482), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n475), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n241), .B1(new_n284), .B2(new_n285), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n487), .A2(new_n488), .A3(new_n489), .A4(new_n480), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n465), .B1(new_n484), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n479), .A2(new_n274), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT68), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(G128), .A3(new_n202), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n211), .B1(new_n496), .B2(new_n198), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n492), .B1(new_n497), .B2(new_n274), .ZN(new_n498));
  OAI21_X1  g312(.A(KEYINPUT12), .B1(new_n498), .B2(new_n488), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n205), .A2(new_n212), .A3(new_n274), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n275), .B1(new_n211), .B2(new_n478), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT12), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n503), .A3(new_n475), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n499), .A2(new_n465), .A3(new_n504), .A4(new_n490), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT80), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n491), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n481), .A2(new_n475), .A3(new_n483), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n503), .B1(new_n502), .B2(new_n475), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n510), .A2(KEYINPUT80), .A3(new_n465), .A4(new_n504), .ZN(new_n511));
  AOI211_X1 g325(.A(G469), .B(G902), .C1(new_n507), .C2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n499), .A2(new_n504), .A3(new_n490), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n464), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT79), .B1(new_n490), .B2(new_n465), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n490), .A2(KEYINPUT79), .A3(new_n465), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n484), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n514), .B(G469), .C1(new_n515), .C2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(G469), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n519), .A2(new_n189), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n461), .B1(new_n512), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n458), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(G214), .B1(G237), .B2(G902), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n320), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n469), .A2(G134), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n471), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G131), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT67), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT67), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n529), .A2(new_n532), .A3(G131), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n531), .A2(new_n474), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n198), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT1), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n537), .B1(new_n222), .B2(G143), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n209), .B1(new_n538), .B2(KEYINPUT68), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n536), .B1(new_n539), .B2(new_n495), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n535), .B1(new_n540), .B2(new_n211), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n475), .B(new_n221), .C1(new_n224), .C2(new_n226), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT66), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT66), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n241), .A2(new_n544), .A3(new_n475), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n541), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT30), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n287), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT69), .B1(new_n497), .B2(new_n534), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT69), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n485), .A2(new_n551), .A3(new_n535), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n547), .B1(new_n241), .B2(new_n475), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n548), .A2(new_n549), .A3(new_n554), .ZN(new_n555));
  XOR2_X1   g369(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n556));
  NAND2_X1  g370(.A1(new_n336), .A2(G210), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT26), .B(G101), .ZN(new_n559));
  XOR2_X1   g373(.A(new_n558), .B(new_n559), .Z(new_n560));
  AOI21_X1  g374(.A(new_n551), .B1(new_n485), .B2(new_n535), .ZN(new_n561));
  AOI211_X1 g375(.A(KEYINPUT69), .B(new_n534), .C1(new_n205), .C2(new_n212), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n549), .B1(new_n241), .B2(new_n475), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n560), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT31), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n555), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT71), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT71), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n555), .A2(new_n565), .A3(new_n569), .A4(new_n566), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n550), .A2(new_n552), .A3(new_n564), .ZN(new_n572));
  AOI22_X1  g386(.A1(new_n485), .A2(new_n535), .B1(new_n542), .B2(KEYINPUT66), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n287), .B1(new_n573), .B2(new_n545), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT28), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT28), .B1(new_n564), .B2(new_n541), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n555), .A2(new_n565), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n578), .A2(new_n560), .B1(new_n579), .B2(KEYINPUT31), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n571), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(G472), .A2(G902), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT32), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT28), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n546), .A2(new_n549), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n550), .A2(new_n552), .A3(new_n564), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n590), .A2(new_n560), .A3(new_n576), .ZN(new_n591));
  INV_X1    g405(.A(new_n560), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n592), .B1(new_n555), .B2(new_n589), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n591), .A2(new_n593), .A3(KEYINPUT29), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT29), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n560), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n550), .A2(new_n552), .A3(new_n542), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n572), .B1(new_n549), .B2(new_n597), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n577), .B(new_n596), .C1(new_n598), .C2(new_n587), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n189), .ZN(new_n600));
  OAI21_X1  g414(.A(G472), .B1(new_n594), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n583), .B1(new_n571), .B2(new_n580), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n586), .B(new_n601), .C1(KEYINPUT32), .C2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(G234), .ZN(new_n604));
  OAI21_X1  g418(.A(G217), .B1(new_n604), .B2(G902), .ZN(new_n605));
  XOR2_X1   g419(.A(new_n605), .B(KEYINPUT72), .Z(new_n606));
  OR2_X1    g420(.A1(new_n209), .A2(G119), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n209), .A2(G119), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT24), .B(G110), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n610), .A2(KEYINPUT73), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n610), .A2(KEYINPUT73), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n609), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT23), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n608), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n209), .A2(KEYINPUT23), .A3(G119), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n615), .A2(new_n607), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(G110), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n617), .A2(KEYINPUT75), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n613), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(KEYINPUT75), .B1(new_n617), .B2(new_n618), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n332), .B(new_n367), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n611), .A2(new_n612), .A3(new_n609), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n617), .A2(new_n618), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n334), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT22), .B(G137), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n459), .A2(new_n604), .A3(G953), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n628), .B(new_n629), .Z(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n622), .A2(new_n626), .A3(new_n630), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(new_n189), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT25), .ZN(new_n635));
  OR2_X1    g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n606), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n632), .A2(new_n633), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n605), .A2(new_n189), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n603), .A2(KEYINPUT76), .A3(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT76), .B1(new_n603), .B2(new_n642), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n527), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT97), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(new_n259), .ZN(G3));
  INV_X1    g462(.A(new_n642), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n523), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n581), .A2(new_n189), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n651), .A2(KEYINPUT98), .A3(G472), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT98), .ZN(new_n653));
  INV_X1    g467(.A(G472), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n581), .B(new_n189), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n650), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n401), .A2(G475), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n383), .A2(new_n387), .A3(new_n384), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n387), .B1(new_n383), .B2(new_n384), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT99), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n425), .A2(new_n435), .A3(new_n407), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n445), .B1(new_n443), .B2(new_n444), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT33), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n189), .A2(G478), .ZN(new_n666));
  OAI22_X1  g480(.A1(new_n665), .A2(new_n666), .B1(G478), .B2(new_n447), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n660), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n525), .ZN(new_n670));
  AOI211_X1 g484(.A(new_n670), .B(new_n398), .C1(new_n315), .C2(new_n319), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n656), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n672), .B(KEYINPUT100), .Z(new_n673));
  XOR2_X1   g487(.A(KEYINPUT34), .B(G104), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G6));
  INV_X1    g489(.A(KEYINPUT101), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n676), .B1(new_n658), .B2(new_n659), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n386), .A2(KEYINPUT101), .A3(new_n388), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n189), .B1(new_n662), .B2(new_n663), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n449), .ZN(new_n681));
  AOI22_X1  g495(.A1(new_n681), .A2(new_n453), .B1(new_n403), .B2(G478), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n450), .A2(new_n404), .ZN(new_n683));
  OAI21_X1  g497(.A(KEYINPUT95), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n684), .A2(new_n455), .A3(new_n657), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n679), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n656), .A2(new_n671), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT35), .B(G107), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G9));
  NOR2_X1   g503(.A1(new_n631), .A2(KEYINPUT36), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n627), .B(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n640), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n638), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n652), .A2(new_n655), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n526), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT37), .B(G110), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G12));
  NOR2_X1   g514(.A1(new_n523), .A2(new_n695), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n320), .A2(new_n525), .A3(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(G900), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n394), .B1(new_n703), .B2(new_n397), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n679), .A2(new_n685), .A3(new_n704), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n603), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G128), .ZN(G30));
  NAND3_X1  g522(.A1(new_n660), .A2(new_n684), .A3(new_n455), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n710), .A2(new_n525), .A3(new_n695), .ZN(new_n711));
  AOI21_X1  g525(.A(G902), .B1(new_n598), .B2(new_n560), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n555), .A2(new_n589), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n592), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n654), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n715), .B1(new_n581), .B2(new_n585), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n716), .B1(KEYINPUT32), .B2(new_n602), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n522), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n507), .A2(new_n511), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n519), .A3(new_n189), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n460), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  XOR2_X1   g536(.A(new_n704), .B(KEYINPUT39), .Z(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI211_X1 g538(.A(new_n711), .B(new_n718), .C1(KEYINPUT40), .C2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n320), .B(new_n726), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n725), .B(new_n727), .C1(KEYINPUT40), .C2(new_n724), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G143), .ZN(G45));
  AOI21_X1  g543(.A(new_n670), .B1(new_n315), .B2(new_n319), .ZN(new_n730));
  INV_X1    g544(.A(new_n704), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n660), .A2(new_n667), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n730), .A2(new_n603), .A3(new_n701), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G146), .ZN(G48));
  AOI21_X1  g549(.A(new_n519), .B1(new_n720), .B2(new_n189), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(new_n512), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT103), .B1(new_n737), .B2(new_n461), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT103), .ZN(new_n739));
  NOR4_X1   g553(.A1(new_n736), .A2(new_n512), .A3(new_n739), .A4(new_n460), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n581), .A2(new_n582), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n584), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n597), .A2(new_n549), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n589), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n576), .B1(new_n745), .B2(KEYINPUT28), .ZN(new_n746));
  AOI21_X1  g560(.A(G902), .B1(new_n746), .B2(new_n596), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n713), .A2(new_n560), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n575), .A2(new_n592), .A3(new_n577), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n749), .A3(new_n595), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n654), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n585), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n752), .B1(new_n571), .B2(new_n580), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n649), .B1(new_n743), .B2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n671), .A2(new_n741), .A3(new_n755), .A4(new_n669), .ZN(new_n756));
  XNOR2_X1  g570(.A(KEYINPUT41), .B(G113), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n756), .B(new_n757), .ZN(G15));
  NAND4_X1  g572(.A1(new_n671), .A2(new_n741), .A3(new_n755), .A4(new_n686), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G116), .ZN(G18));
  NOR2_X1   g574(.A1(new_n458), .A2(new_n695), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n741), .A2(new_n603), .A3(new_n730), .A4(new_n761), .ZN(new_n762));
  XOR2_X1   g576(.A(KEYINPUT104), .B(G119), .Z(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(G21));
  AOI211_X1 g578(.A(new_n670), .B(new_n709), .C1(new_n315), .C2(new_n319), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n654), .B1(new_n581), .B2(new_n189), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n577), .B1(new_n598), .B2(new_n587), .ZN(new_n767));
  AOI22_X1  g581(.A1(new_n767), .A2(new_n560), .B1(KEYINPUT31), .B2(new_n579), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n583), .B1(new_n768), .B2(new_n571), .ZN(new_n769));
  NOR4_X1   g583(.A1(new_n766), .A2(new_n769), .A3(new_n649), .A4(new_n398), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n765), .A2(new_n741), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G122), .ZN(G24));
  NOR4_X1   g586(.A1(new_n766), .A2(new_n732), .A3(new_n769), .A4(new_n695), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n773), .A2(new_n741), .A3(new_n730), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G125), .ZN(G27));
  AND4_X1   g589(.A1(new_n525), .A2(new_n315), .A3(new_n722), .A4(new_n319), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n776), .A2(new_n755), .A3(new_n733), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT42), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n776), .A2(new_n755), .A3(KEYINPUT42), .A4(new_n733), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G131), .ZN(G33));
  NAND3_X1  g596(.A1(new_n776), .A2(new_n755), .A3(new_n705), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G134), .ZN(G36));
  AOI22_X1  g598(.A1(new_n386), .A2(new_n388), .B1(G475), .B2(new_n401), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n667), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT43), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(new_n695), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n652), .A2(new_n655), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(KEYINPUT44), .A3(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n315), .A2(new_n525), .A3(new_n319), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT106), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n514), .B1(new_n515), .B2(new_n517), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n519), .B1(new_n795), .B2(new_n796), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n521), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT46), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n800), .A2(KEYINPUT105), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n799), .A2(KEYINPUT46), .A3(new_n521), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n721), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT105), .B1(new_n800), .B2(new_n801), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n461), .A3(new_n723), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT44), .B1(new_n788), .B2(new_n789), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n794), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(KEYINPUT107), .B(G137), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n810), .B(new_n811), .ZN(G39));
  NAND2_X1  g626(.A1(new_n806), .A2(new_n461), .ZN(new_n813));
  XOR2_X1   g627(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n816), .B1(new_n806), .B2(new_n461), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n603), .A2(new_n642), .A3(new_n732), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(new_n792), .A3(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G140), .ZN(G42));
  NOR2_X1   g635(.A1(new_n787), .A2(new_n393), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n791), .A2(new_n738), .A3(new_n740), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR4_X1   g638(.A1(new_n824), .A2(new_n695), .A3(new_n766), .A4(new_n769), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n823), .A2(new_n642), .A3(new_n394), .A4(new_n718), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n826), .A2(new_n660), .A3(new_n667), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n766), .A2(new_n769), .A3(new_n649), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n822), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n741), .A2(new_n670), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n829), .A2(new_n727), .A3(new_n830), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n831), .A2(KEYINPUT50), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(KEYINPUT50), .ZN(new_n833));
  AOI211_X1 g647(.A(new_n825), .B(new_n827), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n829), .A2(new_n791), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n736), .A2(new_n512), .A3(new_n461), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n835), .B1(new_n818), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n834), .A2(KEYINPUT51), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n586), .A2(new_n601), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n602), .A2(KEYINPUT32), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n642), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n824), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT48), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n720), .A2(new_n189), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(G469), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n461), .A3(new_n721), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n739), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n737), .A2(KEYINPUT103), .A3(new_n461), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n320), .A2(new_n847), .A3(new_n525), .A4(new_n848), .ZN(new_n849));
  OAI221_X1 g663(.A(new_n391), .B1(new_n829), .B2(new_n849), .C1(new_n826), .C2(new_n668), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n843), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n838), .A2(new_n851), .ZN(new_n852));
  XOR2_X1   g666(.A(new_n836), .B(KEYINPUT114), .Z(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n817), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT113), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n855), .B(new_n856), .C1(new_n813), .C2(new_n814), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT113), .B1(new_n815), .B2(new_n817), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n854), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT115), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n860), .A2(new_n861), .A3(new_n835), .ZN(new_n862));
  INV_X1    g676(.A(new_n835), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT115), .B1(new_n859), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n862), .A2(new_n834), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT51), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n852), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n732), .B1(new_n743), .B2(new_n754), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n638), .A2(new_n694), .A3(new_n704), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n869), .B(new_n461), .C1(new_n512), .C2(new_n522), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n870), .B1(new_n743), .B2(new_n716), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n702), .A2(new_n868), .B1(new_n765), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT52), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n872), .A2(new_n873), .A3(new_n707), .A4(new_n774), .ZN(new_n874));
  INV_X1    g688(.A(new_n766), .ZN(new_n875));
  INV_X1    g689(.A(new_n769), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n875), .A2(new_n733), .A3(new_n696), .A4(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n320), .A2(new_n701), .A3(new_n525), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n603), .A2(new_n705), .ZN(new_n879));
  OAI22_X1  g693(.A1(new_n849), .A2(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n869), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n523), .A2(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n730), .A2(new_n717), .A3(new_n710), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n734), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(KEYINPUT52), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT111), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n874), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n886), .B1(new_n874), .B2(new_n885), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n756), .A2(new_n759), .A3(new_n762), .A4(new_n771), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n773), .A2(new_n776), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n657), .A2(new_n451), .A3(new_n454), .A4(new_n731), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n679), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n603), .A2(new_n701), .A3(new_n894), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n783), .B(new_n892), .C1(new_n791), .C2(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n896), .B1(new_n779), .B2(new_n780), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT76), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n841), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n643), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n698), .B1(new_n900), .B2(new_n527), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n447), .A2(G478), .ZN(new_n902));
  INV_X1    g716(.A(new_n665), .ZN(new_n903));
  INV_X1    g717(.A(new_n666), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT109), .B1(new_n785), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n785), .B1(new_n682), .B2(new_n683), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT109), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n660), .A2(new_n667), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n906), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n656), .A2(new_n671), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT110), .B1(new_n901), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n526), .B1(new_n899), .B2(new_n643), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n910), .A2(new_n650), .A3(new_n652), .A4(new_n655), .ZN(new_n914));
  INV_X1    g728(.A(new_n398), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n730), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT110), .ZN(new_n918));
  NOR4_X1   g732(.A1(new_n913), .A2(new_n917), .A3(new_n698), .A4(new_n918), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n891), .B(new_n897), .C1(new_n912), .C2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT53), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n889), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n756), .A2(new_n762), .A3(new_n771), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n315), .A2(new_n722), .A3(new_n319), .A4(new_n525), .ZN(new_n924));
  OAI22_X1  g738(.A1(new_n895), .A2(new_n791), .B1(new_n877), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n705), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n841), .A2(new_n926), .A3(new_n924), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n923), .A2(new_n781), .A3(new_n759), .A4(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n698), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n646), .A2(new_n911), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n918), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n901), .A2(KEYINPUT110), .A3(new_n911), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AND4_X1   g748(.A1(new_n525), .A2(new_n320), .A3(new_n847), .A4(new_n848), .ZN(new_n935));
  AOI22_X1  g749(.A1(new_n935), .A2(new_n773), .B1(new_n702), .B2(new_n706), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n873), .B1(new_n936), .B2(new_n872), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n880), .A2(new_n884), .A3(KEYINPUT52), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT53), .B1(new_n934), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(KEYINPUT54), .B1(new_n922), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT112), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n921), .B1(new_n889), .B2(new_n920), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT54), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n934), .A2(KEYINPUT53), .A3(new_n939), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n941), .A2(new_n942), .A3(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(KEYINPUT111), .B1(new_n937), .B2(new_n938), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n874), .A2(new_n885), .A3(new_n886), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(KEYINPUT53), .B1(new_n934), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n932), .A2(new_n933), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n781), .A2(new_n928), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n953), .A2(new_n890), .ZN(new_n954));
  AND4_X1   g768(.A1(KEYINPUT53), .A2(new_n952), .A3(new_n954), .A4(new_n939), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n951), .A2(new_n955), .A3(KEYINPUT54), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n934), .A2(new_n950), .A3(KEYINPUT53), .ZN(new_n957));
  INV_X1    g771(.A(new_n939), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n921), .B1(new_n920), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n944), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(KEYINPUT112), .B1(new_n956), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n867), .A2(new_n947), .A3(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(G952), .B2(G953), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n642), .A2(new_n525), .A3(new_n461), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n964), .A2(new_n786), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n737), .B(KEYINPUT49), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n965), .A2(new_n966), .A3(new_n718), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n963), .B1(new_n727), .B2(new_n967), .ZN(G75));
  OAI21_X1  g782(.A(G902), .B1(new_n951), .B2(new_n955), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT116), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n943), .A2(new_n945), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n972), .A2(KEYINPUT116), .A3(G902), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n971), .A2(new_n188), .A3(new_n973), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n302), .B(new_n304), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT55), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n976), .A2(KEYINPUT56), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n344), .A2(G952), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT56), .ZN(new_n980));
  INV_X1    g794(.A(G210), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n980), .B1(new_n969), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n979), .B1(new_n982), .B2(new_n976), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n978), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(KEYINPUT117), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT117), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n978), .A2(new_n986), .A3(new_n983), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n985), .A2(new_n987), .ZN(G51));
  NAND2_X1  g802(.A1(new_n972), .A2(KEYINPUT54), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n946), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n520), .B(KEYINPUT57), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(KEYINPUT118), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT118), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n990), .A2(new_n994), .A3(new_n991), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n720), .B(KEYINPUT119), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n993), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n799), .B(KEYINPUT120), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n971), .A2(new_n973), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n979), .B1(new_n997), .B2(new_n999), .ZN(G54));
  INV_X1    g814(.A(new_n979), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n971), .A2(new_n973), .A3(KEYINPUT58), .A4(G475), .ZN(new_n1002));
  INV_X1    g816(.A(new_n383), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT121), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1002), .A2(KEYINPUT121), .A3(new_n1003), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1004), .B1(new_n1007), .B2(new_n1008), .ZN(G60));
  NAND2_X1  g823(.A1(G478), .A2(G902), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1010), .B(KEYINPUT59), .Z(new_n1011));
  AOI21_X1  g825(.A(new_n1011), .B1(new_n961), .B2(new_n947), .ZN(new_n1012));
  OAI21_X1  g826(.A(KEYINPUT122), .B1(new_n1012), .B2(new_n903), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1011), .ZN(new_n1014));
  NOR3_X1   g828(.A1(new_n956), .A2(new_n960), .A3(KEYINPUT112), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n942), .B1(new_n941), .B2(new_n946), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT122), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1017), .A2(new_n1018), .A3(new_n665), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n665), .A2(new_n1011), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n979), .B1(new_n990), .B2(new_n1020), .ZN(new_n1021));
  AND3_X1   g835(.A1(new_n1013), .A2(new_n1019), .A3(new_n1021), .ZN(G63));
  NAND2_X1  g836(.A1(G217), .A2(G902), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(KEYINPUT60), .Z(new_n1024));
  NAND2_X1  g838(.A1(new_n972), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1025), .A2(new_n639), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n972), .A2(new_n691), .A3(new_n1024), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1026), .A2(new_n1001), .A3(new_n1027), .ZN(new_n1028));
  XOR2_X1   g842(.A(new_n1028), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g843(.A(G953), .B1(new_n230), .B2(new_n395), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n890), .B1(new_n932), .B2(new_n933), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1030), .B1(new_n1031), .B2(G953), .ZN(new_n1032));
  INV_X1    g846(.A(new_n302), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1033), .B1(G898), .B2(new_n344), .ZN(new_n1034));
  XNOR2_X1  g848(.A(new_n1032), .B(new_n1034), .ZN(G69));
  AND2_X1   g849(.A1(new_n548), .A2(new_n554), .ZN(new_n1036));
  XOR2_X1   g850(.A(new_n1036), .B(new_n373), .Z(new_n1037));
  AOI21_X1  g851(.A(new_n880), .B1(new_n702), .B2(new_n868), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n728), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g853(.A1(new_n1039), .A2(KEYINPUT62), .ZN(new_n1040));
  XNOR2_X1  g854(.A(new_n1040), .B(KEYINPUT124), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1039), .A2(KEYINPUT62), .ZN(new_n1042));
  OR2_X1    g856(.A1(new_n910), .A2(KEYINPUT125), .ZN(new_n1043));
  AOI21_X1  g857(.A(new_n724), .B1(new_n910), .B2(KEYINPUT125), .ZN(new_n1044));
  NAND4_X1  g858(.A1(new_n900), .A2(new_n792), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  AND4_X1   g859(.A1(new_n810), .A2(new_n820), .A3(new_n1042), .A4(new_n1045), .ZN(new_n1046));
  AOI21_X1  g860(.A(G953), .B1(new_n1041), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g861(.A(KEYINPUT123), .ZN(new_n1048));
  OAI21_X1  g862(.A(new_n1037), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AND2_X1   g863(.A1(new_n810), .A2(new_n820), .ZN(new_n1050));
  INV_X1    g864(.A(KEYINPUT127), .ZN(new_n1051));
  NAND3_X1  g865(.A1(new_n1038), .A2(new_n781), .A3(new_n783), .ZN(new_n1052));
  INV_X1    g866(.A(new_n1052), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n765), .A2(new_n755), .ZN(new_n1054));
  OR3_X1    g868(.A1(new_n807), .A2(KEYINPUT126), .A3(new_n1054), .ZN(new_n1055));
  OAI21_X1  g869(.A(KEYINPUT126), .B1(new_n807), .B2(new_n1054), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g871(.A1(new_n1050), .A2(new_n1051), .A3(new_n1053), .A4(new_n1057), .ZN(new_n1058));
  NAND3_X1  g872(.A1(new_n810), .A2(new_n820), .A3(new_n1057), .ZN(new_n1059));
  OAI21_X1  g873(.A(KEYINPUT127), .B1(new_n1059), .B2(new_n1052), .ZN(new_n1060));
  NAND3_X1  g874(.A1(new_n1058), .A2(new_n344), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g875(.A1(G900), .A2(G953), .ZN(new_n1062));
  AND2_X1   g876(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g877(.A(new_n1037), .ZN(new_n1064));
  OAI21_X1  g878(.A(new_n1064), .B1(new_n1047), .B2(KEYINPUT123), .ZN(new_n1065));
  OAI21_X1  g879(.A(new_n1049), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g880(.A(new_n344), .B1(G227), .B2(G900), .ZN(new_n1067));
  INV_X1    g881(.A(new_n1067), .ZN(new_n1068));
  NAND2_X1  g882(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  OAI211_X1 g883(.A(new_n1067), .B(new_n1049), .C1(new_n1063), .C2(new_n1065), .ZN(new_n1070));
  NAND2_X1  g884(.A1(new_n1069), .A2(new_n1070), .ZN(G72));
  NAND3_X1  g885(.A1(new_n1058), .A2(new_n1031), .A3(new_n1060), .ZN(new_n1072));
  NAND2_X1  g886(.A1(G472), .A2(G902), .ZN(new_n1073));
  XOR2_X1   g887(.A(new_n1073), .B(KEYINPUT63), .Z(new_n1074));
  AOI211_X1 g888(.A(new_n592), .B(new_n713), .C1(new_n1072), .C2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g889(.A1(new_n1041), .A2(new_n1046), .A3(new_n1031), .ZN(new_n1076));
  AOI21_X1  g890(.A(new_n714), .B1(new_n1076), .B2(new_n1074), .ZN(new_n1077));
  NAND2_X1  g891(.A1(new_n748), .A2(new_n579), .ZN(new_n1078));
  NAND2_X1  g892(.A1(new_n1078), .A2(new_n1074), .ZN(new_n1079));
  AOI21_X1  g893(.A(new_n1079), .B1(new_n957), .B2(new_n959), .ZN(new_n1080));
  NOR4_X1   g894(.A1(new_n1075), .A2(new_n1077), .A3(new_n979), .A4(new_n1080), .ZN(G57));
endmodule


