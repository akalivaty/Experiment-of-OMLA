

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734;

  AND2_X1 U368 ( .A1(n710), .A2(KEYINPUT76), .ZN(n361) );
  NOR2_X1 U369 ( .A1(n688), .A2(G902), .ZN(n349) );
  XNOR2_X1 U370 ( .A(n718), .B(G146), .ZN(n518) );
  XNOR2_X1 U371 ( .A(n348), .B(n716), .ZN(n516) );
  XNOR2_X1 U372 ( .A(G137), .B(G140), .ZN(n433) );
  BUF_X1 U373 ( .A(G128), .Z(n384) );
  XNOR2_X2 U374 ( .A(n346), .B(n409), .ZN(n548) );
  AND2_X2 U375 ( .A1(n532), .A2(n531), .ZN(n346) );
  XNOR2_X1 U376 ( .A(n347), .B(KEYINPUT77), .ZN(n547) );
  NAND2_X1 U377 ( .A1(n536), .A2(n537), .ZN(n347) );
  INV_X1 U378 ( .A(n514), .ZN(n348) );
  INV_X2 U379 ( .A(G128), .ZN(n423) );
  XNOR2_X1 U380 ( .A(G113), .B(G140), .ZN(n453) );
  NAND2_X2 U381 ( .A1(n429), .A2(n603), .ZN(n426) );
  XNOR2_X2 U382 ( .A(n452), .B(n352), .ZN(n422) );
  XNOR2_X2 U383 ( .A(n579), .B(KEYINPUT32), .ZN(n730) );
  NOR2_X1 U384 ( .A1(n692), .A2(n703), .ZN(n693) );
  NOR2_X1 U385 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U386 ( .A1(n578), .A2(n650), .ZN(n580) );
  NOR2_X1 U387 ( .A1(n617), .A2(n703), .ZN(n620) );
  AND2_X1 U388 ( .A1(n612), .A2(n428), .ZN(n427) );
  NOR2_X1 U389 ( .A1(n594), .A2(n624), .ZN(n419) );
  XNOR2_X1 U390 ( .A(n559), .B(KEYINPUT33), .ZN(n681) );
  INV_X1 U391 ( .A(n654), .ZN(n582) );
  XNOR2_X1 U392 ( .A(n474), .B(n473), .ZN(n552) );
  AND2_X1 U393 ( .A1(n547), .A2(n545), .ZN(n360) );
  XNOR2_X2 U394 ( .A(n349), .B(n350), .ZN(n529) );
  XOR2_X1 U395 ( .A(KEYINPUT68), .B(G469), .Z(n350) );
  NOR2_X2 U396 ( .A1(n551), .A2(n526), .ZN(n635) );
  NOR2_X2 U397 ( .A1(n728), .A2(n733), .ZN(n424) );
  XNOR2_X2 U398 ( .A(n550), .B(n549), .ZN(n728) );
  INV_X1 U399 ( .A(KEYINPUT107), .ZN(n393) );
  AND2_X1 U400 ( .A1(n400), .A2(n399), .ZN(n398) );
  XNOR2_X1 U401 ( .A(n413), .B(G125), .ZN(n459) );
  INV_X1 U402 ( .A(G146), .ZN(n413) );
  XOR2_X1 U403 ( .A(G104), .B(G122), .Z(n460) );
  XNOR2_X1 U404 ( .A(n459), .B(n412), .ZN(n715) );
  INV_X1 U405 ( .A(KEYINPUT10), .ZN(n412) );
  XNOR2_X1 U406 ( .A(n387), .B(KEYINPUT74), .ZN(n573) );
  INV_X1 U407 ( .A(G472), .ZN(n431) );
  XNOR2_X1 U408 ( .A(n463), .B(n353), .ZN(n533) );
  AND2_X1 U409 ( .A1(n730), .A2(n402), .ZN(n397) );
  NOR2_X1 U410 ( .A1(n730), .A2(n402), .ZN(n401) );
  NOR2_X1 U411 ( .A1(n669), .A2(n593), .ZN(n594) );
  NOR2_X1 U412 ( .A1(n626), .A2(n643), .ZN(n593) );
  NOR2_X1 U413 ( .A1(G953), .A2(G237), .ZN(n504) );
  XNOR2_X1 U414 ( .A(n447), .B(n380), .ZN(n379) );
  INV_X1 U415 ( .A(KEYINPUT86), .ZN(n380) );
  XOR2_X1 U416 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n447) );
  INV_X1 U417 ( .A(n732), .ZN(n373) );
  INV_X1 U418 ( .A(KEYINPUT48), .ZN(n375) );
  XNOR2_X1 U419 ( .A(n479), .B(KEYINPUT23), .ZN(n416) );
  INV_X1 U420 ( .A(KEYINPUT91), .ZN(n479) );
  XNOR2_X1 U421 ( .A(n464), .B(n418), .ZN(n477) );
  INV_X1 U422 ( .A(KEYINPUT8), .ZN(n418) );
  NAND2_X1 U423 ( .A1(n720), .A2(G234), .ZN(n464) );
  XNOR2_X1 U424 ( .A(G134), .B(G122), .ZN(n465) );
  AND2_X2 U425 ( .A1(n427), .A2(n426), .ZN(n695) );
  XNOR2_X1 U426 ( .A(n382), .B(n381), .ZN(n519) );
  INV_X1 U427 ( .A(KEYINPUT108), .ZN(n381) );
  NAND2_X1 U428 ( .A1(n422), .A2(n665), .ZN(n541) );
  XNOR2_X1 U429 ( .A(n439), .B(KEYINPUT1), .ZN(n438) );
  INV_X1 U430 ( .A(KEYINPUT65), .ZN(n439) );
  XNOR2_X1 U431 ( .A(n566), .B(KEYINPUT34), .ZN(n436) );
  NOR2_X1 U432 ( .A1(n681), .A2(n590), .ZN(n566) );
  XNOR2_X1 U433 ( .A(n386), .B(n385), .ZN(n578) );
  INV_X1 U434 ( .A(KEYINPUT22), .ZN(n385) );
  NOR2_X1 U435 ( .A1(n590), .A2(n420), .ZN(n386) );
  NAND2_X1 U436 ( .A1(n571), .A2(n421), .ZN(n420) );
  XNOR2_X1 U437 ( .A(n485), .B(n484), .ZN(n486) );
  NOR2_X1 U438 ( .A1(n699), .A2(G902), .ZN(n487) );
  XNOR2_X1 U439 ( .A(KEYINPUT103), .B(G478), .ZN(n473) );
  INV_X1 U440 ( .A(KEYINPUT6), .ZN(n430) );
  XNOR2_X1 U441 ( .A(n715), .B(n388), .ZN(n461) );
  INV_X1 U442 ( .A(KEYINPUT85), .ZN(n402) );
  XNOR2_X1 U443 ( .A(G137), .B(KEYINPUT70), .ZN(n500) );
  XOR2_X1 U444 ( .A(G119), .B(G116), .Z(n506) );
  XOR2_X1 U445 ( .A(KEYINPUT9), .B(KEYINPUT101), .Z(n466) );
  XNOR2_X1 U446 ( .A(n498), .B(n499), .ZN(n718) );
  XNOR2_X1 U447 ( .A(G131), .B(G134), .ZN(n499) );
  NAND2_X1 U448 ( .A1(G234), .A2(G237), .ZN(n488) );
  INV_X1 U449 ( .A(n719), .ZN(n362) );
  OR2_X1 U450 ( .A1(G237), .A2(G902), .ZN(n511) );
  XNOR2_X1 U451 ( .A(G902), .B(KEYINPUT15), .ZN(n613) );
  INV_X1 U452 ( .A(n570), .ZN(n421) );
  XNOR2_X1 U453 ( .A(n449), .B(G113), .ZN(n503) );
  XNOR2_X1 U454 ( .A(G101), .B(KEYINPUT3), .ZN(n449) );
  XOR2_X1 U455 ( .A(KEYINPUT16), .B(KEYINPUT69), .Z(n443) );
  INV_X1 U456 ( .A(G953), .ZN(n709) );
  XNOR2_X1 U457 ( .A(KEYINPUT45), .B(KEYINPUT79), .ZN(n601) );
  XOR2_X1 U458 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n454) );
  XNOR2_X1 U459 ( .A(n460), .B(n354), .ZN(n388) );
  XOR2_X1 U460 ( .A(KEYINPUT99), .B(KEYINPUT11), .Z(n456) );
  XNOR2_X1 U461 ( .A(G101), .B(G107), .ZN(n512) );
  XNOR2_X1 U462 ( .A(n433), .B(KEYINPUT88), .ZN(n716) );
  XNOR2_X1 U463 ( .A(n372), .B(n705), .ZN(n614) );
  XNOR2_X1 U464 ( .A(n366), .B(n448), .ZN(n372) );
  XNOR2_X1 U465 ( .A(n446), .B(n379), .ZN(n448) );
  AND2_X1 U466 ( .A1(n437), .A2(n558), .ZN(n559) );
  AND2_X1 U467 ( .A1(n649), .A2(n650), .ZN(n437) );
  INV_X1 U468 ( .A(KEYINPUT71), .ZN(n409) );
  XNOR2_X1 U469 ( .A(n541), .B(n355), .ZN(n564) );
  AND2_X1 U470 ( .A1(n357), .A2(n529), .ZN(n525) );
  XNOR2_X1 U471 ( .A(n524), .B(KEYINPUT28), .ZN(n357) );
  XNOR2_X1 U472 ( .A(n417), .B(n480), .ZN(n389) );
  XNOR2_X1 U473 ( .A(n468), .B(n472), .ZN(n376) );
  XNOR2_X1 U474 ( .A(n520), .B(n383), .ZN(n521) );
  XNOR2_X1 U475 ( .A(KEYINPUT109), .B(KEYINPUT43), .ZN(n383) );
  NOR2_X1 U476 ( .A1(n540), .A2(n541), .ZN(n363) );
  XNOR2_X1 U477 ( .A(n539), .B(KEYINPUT113), .ZN(n540) );
  XNOR2_X1 U478 ( .A(n569), .B(KEYINPUT80), .ZN(n434) );
  NOR2_X1 U479 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X2 U480 ( .A1(n572), .A2(n654), .ZN(n630) );
  INV_X1 U481 ( .A(KEYINPUT104), .ZN(n358) );
  NAND2_X1 U482 ( .A1(n552), .A2(n533), .ZN(n359) );
  XNOR2_X1 U483 ( .A(n586), .B(KEYINPUT96), .ZN(n626) );
  NOR2_X1 U484 ( .A1(n585), .A2(n653), .ZN(n586) );
  INV_X1 U485 ( .A(KEYINPUT94), .ZN(n377) );
  NOR2_X1 U486 ( .A1(n370), .A2(n582), .ZN(n624) );
  XNOR2_X1 U487 ( .A(n581), .B(n371), .ZN(n370) );
  INV_X1 U488 ( .A(KEYINPUT83), .ZN(n371) );
  XNOR2_X1 U489 ( .A(n690), .B(n691), .ZN(n692) );
  XOR2_X1 U490 ( .A(n689), .B(KEYINPUT59), .Z(n691) );
  NOR2_X1 U491 ( .A1(n521), .A2(n422), .ZN(n351) );
  AND2_X1 U492 ( .A1(G210), .A2(n511), .ZN(n352) );
  XOR2_X1 U493 ( .A(KEYINPUT13), .B(G475), .Z(n353) );
  XOR2_X1 U494 ( .A(G143), .B(G131), .Z(n354) );
  XNOR2_X1 U495 ( .A(KEYINPUT19), .B(KEYINPUT66), .ZN(n355) );
  XNOR2_X1 U496 ( .A(n411), .B(n389), .ZN(n699) );
  NOR2_X1 U497 ( .A1(n720), .A2(G952), .ZN(n703) );
  INV_X1 U498 ( .A(n703), .ZN(n367) );
  XNOR2_X1 U499 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n356) );
  XNOR2_X1 U500 ( .A(n498), .B(n451), .ZN(n366) );
  XNOR2_X2 U501 ( .A(n471), .B(KEYINPUT4), .ZN(n498) );
  XNOR2_X1 U502 ( .A(n414), .B(n715), .ZN(n411) );
  XNOR2_X2 U503 ( .A(n359), .B(n358), .ZN(n642) );
  XNOR2_X1 U504 ( .A(n376), .B(n469), .ZN(n694) );
  XNOR2_X1 U505 ( .A(n467), .B(n444), .ZN(n468) );
  NOR2_X1 U506 ( .A1(n397), .A2(n404), .ZN(n396) );
  XNOR2_X2 U507 ( .A(n587), .B(n430), .ZN(n387) );
  NAND2_X1 U508 ( .A1(n360), .A2(n546), .ZN(n425) );
  NAND2_X1 U509 ( .A1(n362), .A2(n361), .ZN(n429) );
  XNOR2_X1 U510 ( .A(n363), .B(KEYINPUT36), .ZN(n390) );
  NAND2_X1 U511 ( .A1(n364), .A2(KEYINPUT44), .ZN(n595) );
  NAND2_X1 U512 ( .A1(n597), .A2(n731), .ZN(n364) );
  XNOR2_X1 U513 ( .A(n365), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U514 ( .A1(n368), .A2(n367), .ZN(n365) );
  XNOR2_X1 U515 ( .A(n622), .B(n369), .ZN(n368) );
  INV_X1 U516 ( .A(n623), .ZN(n369) );
  NAND2_X1 U517 ( .A1(n477), .A2(G221), .ZN(n417) );
  NOR2_X1 U518 ( .A1(n387), .A2(n523), .ZN(n510) );
  NAND2_X1 U519 ( .A1(n436), .A2(n568), .ZN(n435) );
  INV_X1 U520 ( .A(n731), .ZN(n404) );
  XNOR2_X1 U521 ( .A(n425), .B(KEYINPUT67), .ZN(n406) );
  AND2_X2 U522 ( .A1(n374), .A2(n373), .ZN(n604) );
  XNOR2_X1 U523 ( .A(n391), .B(n375), .ZN(n374) );
  XNOR2_X1 U524 ( .A(n394), .B(n450), .ZN(n705) );
  XNOR2_X1 U525 ( .A(n378), .B(n377), .ZN(n585) );
  NOR2_X1 U526 ( .A1(n590), .A2(n584), .ZN(n378) );
  OR2_X2 U527 ( .A1(n621), .A2(G902), .ZN(n432) );
  NAND2_X1 U528 ( .A1(n539), .A2(n665), .ZN(n382) );
  XOR2_X2 U529 ( .A(G116), .B(G107), .Z(n470) );
  NAND2_X1 U530 ( .A1(n583), .A2(n635), .ZN(n542) );
  XNOR2_X1 U531 ( .A(n522), .B(KEYINPUT106), .ZN(n583) );
  XNOR2_X1 U532 ( .A(n470), .B(n443), .ZN(n395) );
  XNOR2_X1 U533 ( .A(n395), .B(n503), .ZN(n394) );
  NAND2_X1 U534 ( .A1(n542), .A2(KEYINPUT47), .ZN(n537) );
  XNOR2_X1 U535 ( .A(n433), .B(n416), .ZN(n415) );
  XNOR2_X1 U536 ( .A(n415), .B(n478), .ZN(n414) );
  NAND2_X1 U537 ( .A1(n390), .A2(n650), .ZN(n646) );
  NAND2_X1 U538 ( .A1(n406), .A2(n407), .ZN(n391) );
  XNOR2_X1 U539 ( .A(n518), .B(n509), .ZN(n621) );
  AND2_X2 U540 ( .A1(n392), .A2(n639), .ZN(n539) );
  XNOR2_X1 U541 ( .A(n510), .B(n393), .ZN(n392) );
  NOR2_X1 U542 ( .A1(n730), .A2(n630), .ZN(n597) );
  NAND2_X1 U543 ( .A1(n398), .A2(n396), .ZN(n598) );
  NAND2_X1 U544 ( .A1(n630), .A2(n402), .ZN(n399) );
  NAND2_X1 U545 ( .A1(n403), .A2(n401), .ZN(n400) );
  INV_X1 U546 ( .A(n630), .ZN(n403) );
  XNOR2_X2 U547 ( .A(n405), .B(KEYINPUT0), .ZN(n590) );
  NAND2_X1 U548 ( .A1(n564), .A2(n565), .ZN(n405) );
  INV_X2 U549 ( .A(n491), .ZN(n720) );
  XNOR2_X2 U550 ( .A(G953), .B(KEYINPUT64), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n424), .B(KEYINPUT46), .ZN(n407) );
  XNOR2_X2 U552 ( .A(n408), .B(KEYINPUT39), .ZN(n557) );
  NAND2_X1 U553 ( .A1(n548), .A2(n666), .ZN(n408) );
  NAND2_X1 U554 ( .A1(n419), .A2(n595), .ZN(n596) );
  INV_X1 U555 ( .A(n422), .ZN(n534) );
  XNOR2_X1 U556 ( .A(n534), .B(KEYINPUT38), .ZN(n666) );
  XNOR2_X2 U557 ( .A(n423), .B(G143), .ZN(n471) );
  NAND2_X1 U558 ( .A1(n426), .A2(n612), .ZN(n684) );
  INV_X1 U559 ( .A(n613), .ZN(n428) );
  XNOR2_X2 U560 ( .A(n432), .B(n431), .ZN(n587) );
  XNOR2_X2 U561 ( .A(n435), .B(n434), .ZN(n731) );
  XNOR2_X2 U562 ( .A(n529), .B(n438), .ZN(n650) );
  AND2_X1 U563 ( .A1(n440), .A2(n367), .ZN(G54) );
  XNOR2_X1 U564 ( .A(n442), .B(n441), .ZN(n440) );
  XNOR2_X1 U565 ( .A(n688), .B(n356), .ZN(n441) );
  NAND2_X1 U566 ( .A1(n700), .A2(G469), .ZN(n442) );
  XNOR2_X2 U567 ( .A(n602), .B(n601), .ZN(n710) );
  BUF_X1 U568 ( .A(n695), .Z(n700) );
  INV_X1 U569 ( .A(n459), .ZN(n451) );
  NOR2_X2 U570 ( .A1(n600), .A2(n599), .ZN(n602) );
  XNOR2_X1 U571 ( .A(KEYINPUT102), .B(KEYINPUT7), .ZN(n444) );
  XNOR2_X1 U572 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n445) );
  INV_X1 U573 ( .A(KEYINPUT25), .ZN(n484) );
  NAND2_X1 U574 ( .A1(n695), .A2(G472), .ZN(n622) );
  XNOR2_X1 U575 ( .A(n614), .B(n445), .ZN(n615) );
  XNOR2_X1 U576 ( .A(n616), .B(n615), .ZN(n617) );
  NAND2_X1 U577 ( .A1(G224), .A2(n720), .ZN(n446) );
  XOR2_X1 U578 ( .A(G119), .B(G110), .Z(n478) );
  XOR2_X1 U579 ( .A(n460), .B(n478), .Z(n450) );
  NAND2_X1 U580 ( .A1(n614), .A2(n613), .ZN(n452) );
  XNOR2_X1 U581 ( .A(n454), .B(n453), .ZN(n458) );
  NAND2_X1 U582 ( .A1(G214), .A2(n504), .ZN(n455) );
  XNOR2_X1 U583 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U584 ( .A(n458), .B(n457), .ZN(n462) );
  XNOR2_X1 U585 ( .A(n462), .B(n461), .ZN(n689) );
  NOR2_X1 U586 ( .A1(G902), .A2(n689), .ZN(n463) );
  NAND2_X1 U587 ( .A1(G217), .A2(n477), .ZN(n469) );
  XNOR2_X1 U588 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U589 ( .A(n471), .B(n470), .ZN(n472) );
  NOR2_X1 U590 ( .A1(G902), .A2(n694), .ZN(n474) );
  NOR2_X1 U591 ( .A1(n533), .A2(n552), .ZN(n639) );
  XOR2_X1 U592 ( .A(KEYINPUT90), .B(KEYINPUT24), .Z(n476) );
  XNOR2_X1 U593 ( .A(n384), .B(KEYINPUT89), .ZN(n475) );
  XOR2_X1 U594 ( .A(n476), .B(n475), .Z(n480) );
  XOR2_X1 U595 ( .A(KEYINPUT72), .B(KEYINPUT92), .Z(n483) );
  NAND2_X1 U596 ( .A1(G234), .A2(n613), .ZN(n481) );
  XNOR2_X1 U597 ( .A(KEYINPUT20), .B(n481), .ZN(n495) );
  NAND2_X1 U598 ( .A1(n495), .A2(G217), .ZN(n482) );
  XNOR2_X1 U599 ( .A(n483), .B(n482), .ZN(n485) );
  XNOR2_X2 U600 ( .A(n487), .B(n486), .ZN(n654) );
  XNOR2_X1 U601 ( .A(n488), .B(KEYINPUT14), .ZN(n490) );
  NAND2_X1 U602 ( .A1(G952), .A2(n490), .ZN(n489) );
  XOR2_X1 U603 ( .A(KEYINPUT87), .B(n489), .Z(n679) );
  NOR2_X1 U604 ( .A1(G953), .A2(n679), .ZN(n561) );
  AND2_X1 U605 ( .A1(G902), .A2(n490), .ZN(n560) );
  NAND2_X1 U606 ( .A1(n491), .A2(n560), .ZN(n492) );
  NOR2_X1 U607 ( .A1(G900), .A2(n492), .ZN(n493) );
  NOR2_X1 U608 ( .A1(n561), .A2(n493), .ZN(n494) );
  XOR2_X1 U609 ( .A(KEYINPUT75), .B(n494), .Z(n530) );
  NAND2_X1 U610 ( .A1(n495), .A2(G221), .ZN(n496) );
  XOR2_X1 U611 ( .A(n496), .B(KEYINPUT21), .Z(n655) );
  INV_X1 U612 ( .A(n655), .ZN(n528) );
  NOR2_X1 U613 ( .A1(n530), .A2(n528), .ZN(n497) );
  NAND2_X1 U614 ( .A1(n582), .A2(n497), .ZN(n523) );
  XOR2_X1 U615 ( .A(KEYINPUT95), .B(KEYINPUT5), .Z(n501) );
  XNOR2_X1 U616 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U617 ( .A(n503), .B(n502), .ZN(n508) );
  NAND2_X1 U618 ( .A1(n504), .A2(G210), .ZN(n505) );
  XNOR2_X1 U619 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U620 ( .A(n508), .B(n507), .ZN(n509) );
  NAND2_X1 U621 ( .A1(G214), .A2(n511), .ZN(n665) );
  XOR2_X1 U622 ( .A(G104), .B(G110), .Z(n513) );
  XNOR2_X1 U623 ( .A(n513), .B(n512), .ZN(n514) );
  NAND2_X1 U624 ( .A1(G227), .A2(n720), .ZN(n515) );
  XNOR2_X1 U625 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U626 ( .A(n518), .B(n517), .ZN(n688) );
  INV_X1 U627 ( .A(n650), .ZN(n575) );
  NAND2_X1 U628 ( .A1(n519), .A2(n575), .ZN(n520) );
  XNOR2_X1 U629 ( .A(KEYINPUT110), .B(n351), .ZN(n732) );
  XOR2_X1 U630 ( .A(KEYINPUT105), .B(n642), .Z(n556) );
  OR2_X1 U631 ( .A1(n556), .A2(n639), .ZN(n522) );
  NOR2_X1 U632 ( .A1(n523), .A2(n587), .ZN(n524) );
  XNOR2_X1 U633 ( .A(KEYINPUT111), .B(n525), .ZN(n551) );
  INV_X1 U634 ( .A(n564), .ZN(n526) );
  INV_X1 U635 ( .A(n587), .ZN(n653) );
  NAND2_X1 U636 ( .A1(n653), .A2(n665), .ZN(n527) );
  XOR2_X1 U637 ( .A(KEYINPUT30), .B(n527), .Z(n532) );
  XOR2_X1 U638 ( .A(KEYINPUT93), .B(n528), .Z(n570) );
  NOR2_X2 U639 ( .A1(n582), .A2(n570), .ZN(n649) );
  NAND2_X1 U640 ( .A1(n649), .A2(n529), .ZN(n584) );
  NOR2_X1 U641 ( .A1(n584), .A2(n530), .ZN(n531) );
  INV_X1 U642 ( .A(n533), .ZN(n553) );
  NAND2_X1 U643 ( .A1(n553), .A2(n552), .ZN(n567) );
  NOR2_X1 U644 ( .A1(n534), .A2(n567), .ZN(n535) );
  NAND2_X1 U645 ( .A1(n548), .A2(n535), .ZN(n633) );
  XNOR2_X1 U646 ( .A(n633), .B(KEYINPUT78), .ZN(n536) );
  XNOR2_X1 U647 ( .A(n646), .B(KEYINPUT82), .ZN(n546) );
  INV_X1 U648 ( .A(KEYINPUT47), .ZN(n544) );
  INV_X1 U649 ( .A(n542), .ZN(n543) );
  NAND2_X1 U650 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U651 ( .A(KEYINPUT112), .B(KEYINPUT40), .Z(n550) );
  NAND2_X1 U652 ( .A1(n557), .A2(n639), .ZN(n549) );
  NAND2_X1 U653 ( .A1(n666), .A2(n665), .ZN(n670) );
  NOR2_X1 U654 ( .A1(n553), .A2(n552), .ZN(n571) );
  INV_X1 U655 ( .A(n571), .ZN(n668) );
  NOR2_X1 U656 ( .A1(n670), .A2(n668), .ZN(n554) );
  XNOR2_X1 U657 ( .A(n554), .B(KEYINPUT41), .ZN(n680) );
  NOR2_X1 U658 ( .A1(n551), .A2(n680), .ZN(n555) );
  XNOR2_X1 U659 ( .A(KEYINPUT42), .B(n555), .ZN(n733) );
  NAND2_X1 U660 ( .A1(n557), .A2(n556), .ZN(n648) );
  NAND2_X1 U661 ( .A1(n604), .A2(n648), .ZN(n719) );
  INV_X1 U662 ( .A(KEYINPUT76), .ZN(n605) );
  INV_X1 U663 ( .A(n387), .ZN(n558) );
  NOR2_X1 U664 ( .A1(G898), .A2(n709), .ZN(n704) );
  NAND2_X1 U665 ( .A1(n704), .A2(n560), .ZN(n563) );
  INV_X1 U666 ( .A(n561), .ZN(n562) );
  NAND2_X1 U667 ( .A1(n563), .A2(n562), .ZN(n565) );
  INV_X1 U668 ( .A(n567), .ZN(n568) );
  INV_X1 U669 ( .A(KEYINPUT35), .ZN(n569) );
  NAND2_X1 U670 ( .A1(n580), .A2(n587), .ZN(n572) );
  NAND2_X1 U671 ( .A1(n573), .A2(n582), .ZN(n574) );
  XNOR2_X1 U672 ( .A(n576), .B(KEYINPUT73), .ZN(n577) );
  NOR2_X1 U673 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U674 ( .A1(n580), .A2(n387), .ZN(n581) );
  INV_X1 U675 ( .A(n583), .ZN(n669) );
  NAND2_X1 U676 ( .A1(n650), .A2(n649), .ZN(n588) );
  NOR2_X1 U677 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U678 ( .A(n589), .B(KEYINPUT97), .ZN(n659) );
  NOR2_X1 U679 ( .A1(n590), .A2(n659), .ZN(n592) );
  XOR2_X1 U680 ( .A(KEYINPUT98), .B(KEYINPUT31), .Z(n591) );
  XNOR2_X1 U681 ( .A(n592), .B(n591), .ZN(n643) );
  XNOR2_X1 U682 ( .A(n596), .B(KEYINPUT84), .ZN(n600) );
  NOR2_X1 U683 ( .A1(n598), .A2(KEYINPUT44), .ZN(n599) );
  INV_X1 U684 ( .A(KEYINPUT2), .ZN(n603) );
  INV_X1 U685 ( .A(n604), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n605), .A2(n648), .ZN(n608) );
  NAND2_X1 U687 ( .A1(n648), .A2(KEYINPUT2), .ZN(n606) );
  NAND2_X1 U688 ( .A1(n606), .A2(KEYINPUT76), .ZN(n607) );
  NAND2_X1 U689 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U690 ( .A1(n611), .A2(n710), .ZN(n612) );
  NAND2_X1 U691 ( .A1(n695), .A2(G210), .ZN(n616) );
  XOR2_X1 U692 ( .A(KEYINPUT122), .B(KEYINPUT56), .Z(n618) );
  XNOR2_X1 U693 ( .A(KEYINPUT81), .B(n618), .ZN(n619) );
  XNOR2_X1 U694 ( .A(n620), .B(n619), .ZN(G51) );
  XNOR2_X1 U695 ( .A(n621), .B(KEYINPUT62), .ZN(n623) );
  XOR2_X1 U696 ( .A(n624), .B(G101), .Z(G3) );
  NAND2_X1 U697 ( .A1(n626), .A2(n639), .ZN(n625) );
  XNOR2_X1 U698 ( .A(n625), .B(G104), .ZN(G6) );
  XOR2_X1 U699 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n628) );
  NAND2_X1 U700 ( .A1(n626), .A2(n642), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U702 ( .A(G107), .B(n629), .ZN(G9) );
  XOR2_X1 U703 ( .A(G110), .B(n630), .Z(G12) );
  XOR2_X1 U704 ( .A(n384), .B(KEYINPUT29), .Z(n632) );
  NAND2_X1 U705 ( .A1(n635), .A2(n642), .ZN(n631) );
  XNOR2_X1 U706 ( .A(n632), .B(n631), .ZN(G30) );
  XNOR2_X1 U707 ( .A(G143), .B(KEYINPUT114), .ZN(n634) );
  XNOR2_X1 U708 ( .A(n634), .B(n633), .ZN(G45) );
  XOR2_X1 U709 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n637) );
  NAND2_X1 U710 ( .A1(n635), .A2(n639), .ZN(n636) );
  XNOR2_X1 U711 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U712 ( .A(G146), .B(n638), .ZN(G48) );
  XOR2_X1 U713 ( .A(G113), .B(KEYINPUT117), .Z(n641) );
  NAND2_X1 U714 ( .A1(n639), .A2(n643), .ZN(n640) );
  XNOR2_X1 U715 ( .A(n641), .B(n640), .ZN(G15) );
  NAND2_X1 U716 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U717 ( .A(n644), .B(KEYINPUT118), .ZN(n645) );
  XNOR2_X1 U718 ( .A(G116), .B(n645), .ZN(G18) );
  XOR2_X1 U719 ( .A(G125), .B(KEYINPUT37), .Z(n647) );
  XNOR2_X1 U720 ( .A(n646), .B(n647), .ZN(G27) );
  XNOR2_X1 U721 ( .A(G134), .B(n648), .ZN(G36) );
  XOR2_X1 U722 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n662) );
  NOR2_X1 U723 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U724 ( .A(n651), .B(KEYINPUT50), .ZN(n652) );
  NOR2_X1 U725 ( .A1(n653), .A2(n652), .ZN(n658) );
  NOR2_X1 U726 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U727 ( .A(n656), .B(KEYINPUT49), .ZN(n657) );
  NAND2_X1 U728 ( .A1(n658), .A2(n657), .ZN(n660) );
  NAND2_X1 U729 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U730 ( .A(n662), .B(n661), .ZN(n663) );
  NOR2_X1 U731 ( .A1(n663), .A2(n680), .ZN(n664) );
  XNOR2_X1 U732 ( .A(n664), .B(KEYINPUT120), .ZN(n676) );
  NOR2_X1 U733 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U734 ( .A1(n668), .A2(n667), .ZN(n673) );
  NOR2_X1 U735 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U736 ( .A(KEYINPUT121), .B(n671), .Z(n672) );
  NOR2_X1 U737 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U738 ( .A1(n681), .A2(n674), .ZN(n675) );
  NOR2_X1 U739 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U740 ( .A(n677), .B(KEYINPUT52), .ZN(n678) );
  NOR2_X1 U741 ( .A1(n679), .A2(n678), .ZN(n683) );
  NOR2_X1 U742 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U743 ( .A1(n683), .A2(n682), .ZN(n685) );
  NAND2_X1 U744 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U745 ( .A1(n686), .A2(G953), .ZN(n687) );
  XNOR2_X1 U746 ( .A(n687), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U747 ( .A1(n695), .A2(G475), .ZN(n690) );
  XNOR2_X1 U748 ( .A(n693), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U749 ( .A(n694), .B(KEYINPUT123), .Z(n697) );
  NAND2_X1 U750 ( .A1(n700), .A2(G478), .ZN(n696) );
  XNOR2_X1 U751 ( .A(n697), .B(n696), .ZN(n698) );
  NOR2_X1 U752 ( .A1(n703), .A2(n698), .ZN(G63) );
  NAND2_X1 U753 ( .A1(G217), .A2(n700), .ZN(n701) );
  XNOR2_X1 U754 ( .A(n699), .B(n701), .ZN(n702) );
  NOR2_X1 U755 ( .A1(n703), .A2(n702), .ZN(G66) );
  NOR2_X1 U756 ( .A1(n705), .A2(n704), .ZN(n714) );
  NAND2_X1 U757 ( .A1(G953), .A2(G224), .ZN(n706) );
  XNOR2_X1 U758 ( .A(KEYINPUT61), .B(n706), .ZN(n707) );
  NAND2_X1 U759 ( .A1(n707), .A2(G898), .ZN(n708) );
  XNOR2_X1 U760 ( .A(n708), .B(KEYINPUT124), .ZN(n712) );
  NAND2_X1 U761 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U762 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U763 ( .A(n714), .B(n713), .ZN(G69) );
  XNOR2_X1 U764 ( .A(n716), .B(n715), .ZN(n717) );
  XNOR2_X1 U765 ( .A(n718), .B(n717), .ZN(n722) );
  XNOR2_X1 U766 ( .A(n722), .B(n719), .ZN(n721) );
  NAND2_X1 U767 ( .A1(n721), .A2(n720), .ZN(n727) );
  XNOR2_X1 U768 ( .A(G227), .B(n722), .ZN(n723) );
  NAND2_X1 U769 ( .A1(n723), .A2(G900), .ZN(n724) );
  XOR2_X1 U770 ( .A(KEYINPUT125), .B(n724), .Z(n725) );
  NAND2_X1 U771 ( .A1(G953), .A2(n725), .ZN(n726) );
  NAND2_X1 U772 ( .A1(n727), .A2(n726), .ZN(G72) );
  XOR2_X1 U773 ( .A(G131), .B(n728), .Z(G33) );
  XOR2_X1 U774 ( .A(G119), .B(KEYINPUT126), .Z(n729) );
  XNOR2_X1 U775 ( .A(n730), .B(n729), .ZN(G21) );
  XNOR2_X1 U776 ( .A(n731), .B(G122), .ZN(G24) );
  XOR2_X1 U777 ( .A(G140), .B(n732), .Z(G42) );
  XNOR2_X1 U778 ( .A(G137), .B(KEYINPUT127), .ZN(n734) );
  XNOR2_X1 U779 ( .A(n734), .B(n733), .ZN(G39) );
endmodule

