//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT64), .ZN(new_n209));
  XOR2_X1   g0009(.A(KEYINPUT67), .B(G68), .Z(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G107), .A2(G264), .ZN(new_n217));
  NAND4_X1  g0017(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n209), .B1(new_n213), .B2(new_n218), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT68), .Z(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT69), .Z(new_n222));
  NOR2_X1   g0022(.A1(new_n209), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT0), .Z(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(new_n201), .ZN(new_n229));
  INV_X1    g0029(.A(KEYINPUT65), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n202), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n231), .B1(new_n230), .B2(new_n229), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT66), .Z(new_n233));
  AOI21_X1  g0033(.A(new_n225), .B1(new_n228), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n220), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n222), .A2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  INV_X1    g0045(.A(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT70), .B(G50), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XOR2_X1   g0050(.A(G107), .B(G116), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(G41), .ZN(new_n254));
  INV_X1    g0054(.A(G45), .ZN(new_n255));
  AOI21_X1  g0055(.A(G1), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G274), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n256), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G244), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n257), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT73), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI211_X1 g0065(.A(KEYINPUT73), .B(new_n257), .C1(new_n261), .C2(new_n262), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT3), .B(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(G107), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n212), .A2(G1698), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n269), .B1(G232), .B2(G1698), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n268), .B1(new_n267), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n258), .A2(KEYINPUT71), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT71), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(new_n254), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n273), .B1(new_n275), .B2(new_n226), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n271), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n265), .A2(new_n266), .A3(new_n279), .ZN(new_n280));
  OR3_X1    g0080(.A1(new_n280), .A2(KEYINPUT76), .A3(G179), .ZN(new_n281));
  OAI21_X1  g0081(.A(KEYINPUT76), .B1(new_n280), .B2(G179), .ZN(new_n282));
  INV_X1    g0082(.A(G169), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT75), .ZN(new_n284));
  NAND3_X1  g0084(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n226), .ZN(new_n286));
  INV_X1    g0086(.A(G1), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n286), .B1(new_n287), .B2(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G77), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n284), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n288), .A2(KEYINPUT75), .A3(G77), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n287), .A2(G13), .A3(G20), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n291), .A2(new_n292), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(KEYINPUT8), .B(G58), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT74), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT72), .B1(G20), .B2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NOR3_X1   g0099(.A1(KEYINPUT72), .A2(G20), .A3(G33), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g0102(.A(KEYINPUT15), .B(G87), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n227), .A2(G33), .ZN(new_n304));
  OAI22_X1  g0104(.A1(new_n303), .A2(new_n304), .B1(new_n227), .B2(new_n290), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n286), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n283), .A2(new_n280), .B1(new_n295), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n281), .A2(new_n282), .A3(new_n307), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n295), .A2(new_n306), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n280), .A2(G200), .ZN(new_n310));
  INV_X1    g0110(.A(G190), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n309), .B(new_n310), .C1(new_n311), .C2(new_n280), .ZN(new_n312));
  AND2_X1   g0112(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n203), .A2(G20), .ZN(new_n314));
  INV_X1    g0114(.A(G150), .ZN(new_n315));
  OAI221_X1 g0115(.A(new_n314), .B1(new_n296), .B2(new_n304), .C1(new_n301), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n286), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n293), .A2(G50), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n318), .B1(new_n288), .B2(G50), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n267), .A2(G223), .A3(G1698), .ZN(new_n321));
  INV_X1    g0121(.A(G1698), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n267), .A2(G222), .A3(new_n322), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n321), .B(new_n323), .C1(new_n290), .C2(new_n267), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n278), .ZN(new_n325));
  INV_X1    g0125(.A(new_n257), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n258), .A2(new_n256), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n326), .B1(new_n327), .B2(G226), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n320), .B1(new_n330), .B2(G169), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n329), .A2(G179), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT9), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n317), .A2(new_n334), .A3(new_n319), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n334), .B1(new_n317), .B2(new_n319), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n329), .A2(G200), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n325), .A2(G190), .A3(new_n328), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT10), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n337), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n335), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT10), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n344), .A2(new_n339), .A3(new_n345), .A4(new_n340), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n333), .B1(new_n342), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n211), .A2(G20), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(new_n290), .B2(new_n304), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n301), .A2(new_n202), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n286), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  XNOR2_X1  g0151(.A(new_n351), .B(KEYINPUT11), .ZN(new_n352));
  INV_X1    g0152(.A(G13), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(G1), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT12), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n348), .A2(new_n355), .B1(KEYINPUT12), .B2(new_n294), .ZN(new_n356));
  INV_X1    g0156(.A(G68), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n357), .B1(new_n289), .B2(KEYINPUT12), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n352), .A2(new_n359), .ZN(new_n360));
  OR2_X1    g0160(.A1(new_n283), .A2(KEYINPUT78), .ZN(new_n361));
  INV_X1    g0161(.A(G97), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT77), .B1(new_n274), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT77), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n364), .A2(G33), .A3(G97), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G226), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n322), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n267), .B(new_n368), .C1(G232), .C2(new_n322), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n277), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n257), .B1(new_n261), .B2(new_n212), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT13), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT13), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n326), .B1(new_n327), .B2(G238), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n369), .A2(new_n366), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n373), .B(new_n374), .C1(new_n375), .C2(new_n277), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n361), .B1(new_n372), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT14), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n372), .A2(new_n376), .ZN(new_n379));
  INV_X1    g0179(.A(G179), .ZN(new_n380));
  OAI22_X1  g0180(.A1(new_n377), .A2(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AOI211_X1 g0181(.A(KEYINPUT14), .B(new_n361), .C1(new_n372), .C2(new_n376), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n360), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n379), .A2(G200), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n372), .A2(G190), .A3(new_n376), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n352), .A2(new_n359), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n313), .A2(new_n347), .A3(new_n383), .A4(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n296), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n388), .A2(new_n294), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n389), .B1(new_n289), .B2(new_n388), .ZN(new_n390));
  INV_X1    g0190(.A(new_n286), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT79), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT3), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(G33), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT80), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n397), .B1(KEYINPUT3), .B2(new_n274), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT7), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n394), .A2(new_n397), .A3(G33), .A4(new_n395), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n399), .A2(new_n400), .A3(new_n227), .A4(new_n401), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n402), .A2(G68), .ZN(new_n403));
  AND2_X1   g0203(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n404));
  NOR2_X1   g0204(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n405));
  NOR3_X1   g0205(.A1(new_n404), .A2(new_n405), .A3(new_n274), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n274), .A2(KEYINPUT3), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT80), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n401), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT7), .B1(new_n409), .B2(G20), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT81), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT67), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n412), .A2(G68), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n357), .A2(KEYINPUT67), .ZN(new_n414));
  OAI21_X1  g0214(.A(G58), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n227), .B1(new_n415), .B2(new_n229), .ZN(new_n416));
  INV_X1    g0216(.A(G159), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n301), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n411), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  OR3_X1    g0219(.A1(KEYINPUT72), .A2(G20), .A3(G33), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n298), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(G159), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n201), .B1(new_n210), .B2(G58), .ZN(new_n423));
  OAI211_X1 g0223(.A(KEYINPUT81), .B(new_n422), .C1(new_n423), .C2(new_n227), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n403), .A2(new_n410), .B1(new_n419), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n391), .B1(new_n425), .B2(KEYINPUT16), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT16), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n393), .A2(G33), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n407), .ZN(new_n429));
  AOI21_X1  g0229(.A(KEYINPUT7), .B1(new_n429), .B2(new_n227), .ZN(new_n430));
  INV_X1    g0230(.A(new_n428), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n274), .B1(new_n404), .B2(new_n405), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n431), .B1(new_n432), .B2(KEYINPUT82), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT82), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n434), .B(new_n274), .C1(new_n404), .C2(new_n405), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n400), .A2(G20), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n430), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n438), .A2(new_n211), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n416), .A2(new_n418), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n427), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n390), .B1(new_n426), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n367), .A2(G1698), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(G223), .B2(G1698), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n445), .B1(new_n399), .B2(new_n401), .ZN(new_n446));
  INV_X1    g0246(.A(G87), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n274), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n278), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n326), .B1(new_n327), .B2(G232), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(G169), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n380), .B2(new_n451), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT18), .B1(new_n443), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n390), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n410), .A2(G68), .A3(new_n402), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n419), .A2(new_n424), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n457), .A2(new_n458), .A3(KEYINPUT16), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n286), .ZN(new_n460));
  AOI211_X1 g0260(.A(new_n400), .B(G20), .C1(new_n433), .C2(new_n435), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n210), .B1(new_n461), .B2(new_n430), .ZN(new_n462));
  AOI21_X1  g0262(.A(KEYINPUT16), .B1(new_n462), .B2(new_n440), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n456), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT18), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(new_n465), .A3(new_n453), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n449), .A2(G190), .A3(new_n450), .ZN(new_n467));
  INV_X1    g0267(.A(G200), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n468), .B1(new_n449), .B2(new_n450), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n456), .B(new_n470), .C1(new_n460), .C2(new_n463), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT17), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n426), .A2(new_n442), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n474), .A2(KEYINPUT17), .A3(new_n456), .A4(new_n470), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n455), .A2(new_n466), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT83), .ZN(new_n477));
  OR3_X1    g0277(.A1(new_n387), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n477), .B1(new_n387), .B2(new_n476), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n294), .A2(new_n362), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n287), .A2(G33), .ZN(new_n482));
  AND4_X1   g0282(.A1(new_n226), .A2(new_n293), .A3(new_n285), .A4(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n481), .B1(new_n484), .B2(new_n362), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  XNOR2_X1  g0286(.A(G97), .B(G107), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT6), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NOR3_X1   g0289(.A1(new_n488), .A2(new_n362), .A3(G107), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI22_X1  g0291(.A1(new_n491), .A2(new_n227), .B1(new_n290), .B2(new_n301), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n436), .A2(new_n437), .ZN(new_n493));
  INV_X1    g0293(.A(new_n430), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n492), .B1(new_n495), .B2(G107), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n486), .B1(new_n496), .B2(new_n391), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n255), .A2(G1), .ZN(new_n498));
  XNOR2_X1  g0298(.A(KEYINPUT5), .B(G41), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n258), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G257), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n259), .A2(G274), .A3(new_n498), .A4(new_n499), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n262), .A2(G1698), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n506));
  OAI21_X1  g0306(.A(KEYINPUT85), .B1(new_n506), .B2(new_n429), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n267), .A2(G250), .A3(G1698), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT85), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n267), .A2(new_n509), .A3(KEYINPUT4), .A4(new_n505), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G283), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n507), .A2(new_n508), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n505), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n513), .B1(new_n399), .B2(new_n401), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT84), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT4), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n409), .A2(new_n505), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT84), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n512), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n380), .B(new_n504), .C1(new_n519), .C2(new_n277), .ZN(new_n520));
  INV_X1    g0320(.A(new_n512), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT4), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(new_n517), .B2(KEYINPUT84), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n514), .A2(new_n515), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n503), .B1(new_n525), .B2(new_n278), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n497), .B(new_n520), .C1(new_n526), .C2(G169), .ZN(new_n527));
  OR2_X1    g0327(.A1(new_n489), .A2(new_n490), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n528), .A2(G20), .B1(G77), .B2(new_n421), .ZN(new_n529));
  INV_X1    g0329(.A(G107), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n529), .B1(new_n438), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n485), .B1(new_n531), .B2(new_n286), .ZN(new_n532));
  OAI211_X1 g0332(.A(G190), .B(new_n504), .C1(new_n519), .C2(new_n277), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n532), .B(new_n533), .C1(new_n526), .C2(new_n468), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n527), .A2(new_n534), .ZN(new_n535));
  AND2_X1   g0335(.A1(KEYINPUT22), .A2(G87), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n409), .A2(new_n227), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT24), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n447), .A2(G20), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT22), .B1(new_n267), .B2(new_n539), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n530), .A2(KEYINPUT23), .A3(G20), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT23), .B1(new_n530), .B2(G20), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G116), .ZN(new_n543));
  OAI22_X1  g0343(.A1(new_n541), .A2(new_n542), .B1(G20), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n537), .A2(new_n538), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n538), .B1(new_n537), .B2(new_n545), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n286), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n500), .A2(G264), .ZN(new_n549));
  INV_X1    g0349(.A(G294), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n274), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(G257), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G1698), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(G250), .B2(G1698), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n551), .B1(new_n409), .B2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n502), .B(new_n549), .C1(new_n556), .C2(new_n277), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G200), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT87), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT25), .ZN(new_n560));
  AOI211_X1 g0360(.A(G107), .B(new_n293), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n559), .A2(new_n560), .ZN(new_n562));
  OR2_X1    g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n562), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n563), .A2(new_n564), .B1(G107), .B2(new_n483), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n554), .B1(new_n399), .B2(new_n401), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n278), .B1(new_n566), .B2(new_n551), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n567), .A2(G190), .A3(new_n502), .A4(new_n549), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n548), .A2(new_n558), .A3(new_n565), .A4(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT19), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n570), .B1(new_n363), .B2(new_n365), .ZN(new_n571));
  OAI22_X1  g0371(.A1(new_n571), .A2(G20), .B1(G87), .B2(new_n206), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n570), .B1(new_n304), .B2(new_n362), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI211_X1 g0374(.A(G20), .B(new_n357), .C1(new_n399), .C2(new_n401), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n286), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n303), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n577), .A2(new_n293), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n483), .A2(new_n577), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n576), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n262), .A2(G1698), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(G238), .B2(G1698), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n583), .B1(new_n399), .B2(new_n401), .ZN(new_n584));
  INV_X1    g0384(.A(new_n543), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n278), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(G250), .ZN(new_n587));
  NOR3_X1   g0387(.A1(new_n258), .A2(new_n587), .A3(new_n498), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(G274), .B2(new_n498), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n283), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n586), .A2(new_n380), .A3(new_n589), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n581), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n590), .A2(G200), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n409), .A2(new_n227), .A3(G68), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n595), .A2(new_n573), .A3(new_n572), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n578), .B1(new_n596), .B2(new_n286), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n483), .A2(G87), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n586), .A2(G190), .A3(new_n589), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n594), .A2(new_n597), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n569), .A2(new_n593), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n537), .A2(new_n545), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT24), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n537), .A2(new_n538), .A3(new_n545), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n391), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n565), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n557), .A2(new_n283), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n567), .A2(new_n380), .A3(new_n502), .A4(new_n549), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n500), .A2(G270), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n502), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(G257), .A2(G1698), .ZN(new_n615));
  INV_X1    g0415(.A(G264), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n615), .B1(new_n616), .B2(G1698), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n618), .B1(new_n399), .B2(new_n401), .ZN(new_n619));
  INV_X1    g0419(.A(G303), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n267), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n278), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n614), .A2(new_n622), .A3(G190), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n511), .B(new_n227), .C1(G33), .C2(new_n362), .ZN(new_n624));
  INV_X1    g0424(.A(G116), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(G20), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n286), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT20), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n624), .A2(KEYINPUT20), .A3(new_n286), .A4(new_n626), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT86), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n293), .B2(G116), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n354), .A2(KEYINPUT86), .A3(G20), .A4(new_n625), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n483), .A2(G116), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n409), .A2(new_n617), .ZN(new_n638));
  INV_X1    g0438(.A(new_n621), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n277), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(new_n613), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n623), .B(new_n637), .C1(new_n641), .C2(new_n468), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT21), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n283), .B1(new_n631), .B2(new_n635), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n643), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n644), .B(KEYINPUT21), .C1(new_n640), .C2(new_n613), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n614), .A2(new_n622), .A3(new_n636), .A4(G179), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n642), .A2(new_n646), .A3(new_n647), .A4(new_n648), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n601), .A2(new_n611), .A3(new_n649), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n480), .A2(new_n535), .A3(new_n650), .ZN(G372));
  NAND2_X1  g0451(.A1(new_n593), .A2(new_n600), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n504), .B1(new_n519), .B2(new_n277), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n532), .B1(new_n654), .B2(new_n283), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n653), .A2(new_n655), .A3(KEYINPUT26), .A4(new_n520), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n527), .B2(new_n652), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n569), .A2(new_n593), .A3(new_n600), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n609), .B(new_n608), .C1(new_n605), .C2(new_n606), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n647), .A2(new_n648), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n614), .A2(new_n622), .ZN(new_n663));
  AOI21_X1  g0463(.A(KEYINPUT21), .B1(new_n663), .B2(new_n644), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n660), .A2(new_n666), .A3(new_n527), .A4(new_n534), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n593), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n480), .B1(new_n659), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n383), .A2(new_n308), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n670), .A2(new_n473), .A3(new_n475), .A4(new_n386), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n455), .A2(new_n466), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n342), .A2(new_n346), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n333), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n669), .A2(new_n675), .ZN(G369));
  NAND2_X1  g0476(.A1(new_n354), .A2(new_n227), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n665), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n682), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n569), .B1(new_n607), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n661), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n661), .B2(new_n682), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT88), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT88), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n684), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n661), .A2(new_n682), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n689), .A2(new_n690), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n685), .A2(new_n637), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n662), .B2(new_n664), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n649), .B2(new_n695), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n693), .A2(new_n700), .ZN(G399));
  INV_X1    g0501(.A(new_n223), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(G41), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(G1), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n232), .B2(new_n704), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT28), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT29), .ZN(new_n709));
  INV_X1    g0509(.A(new_n593), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n601), .B1(new_n665), .B2(new_n661), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n710), .B1(new_n711), .B2(new_n535), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT89), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n656), .A2(new_n658), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n527), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n715), .A2(KEYINPUT89), .A3(KEYINPUT26), .A4(new_n653), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n712), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n709), .B1(new_n717), .B2(new_n685), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n656), .A2(new_n658), .ZN(new_n719));
  AOI211_X1 g0519(.A(KEYINPUT29), .B(new_n682), .C1(new_n712), .C2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n650), .A2(new_n535), .A3(new_n685), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n586), .A2(new_n567), .A3(new_n589), .A4(new_n549), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n614), .A2(new_n622), .A3(G179), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n723), .B1(new_n726), .B2(new_n654), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n724), .A2(new_n725), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n526), .A2(new_n728), .A3(KEYINPUT30), .ZN(new_n729));
  AND3_X1   g0529(.A1(new_n663), .A2(new_n590), .A3(new_n380), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(new_n654), .A3(new_n557), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n727), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n682), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT31), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n732), .A2(KEYINPUT31), .A3(new_n682), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n722), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G330), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n721), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n708), .B1(new_n740), .B2(G1), .ZN(G364));
  NOR2_X1   g0541(.A1(new_n353), .A2(G20), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G45), .ZN(new_n743));
  OR2_X1    g0543(.A1(new_n743), .A2(KEYINPUT90), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n287), .B1(new_n743), .B2(KEYINPUT90), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OR3_X1    g0546(.A1(new_n703), .A2(KEYINPUT91), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(KEYINPUT91), .B1(new_n703), .B2(new_n746), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n699), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(G330), .B2(new_n697), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G13), .A2(G33), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n226), .B1(G20), .B2(new_n283), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n702), .A2(new_n429), .ZN(new_n759));
  XOR2_X1   g0559(.A(new_n759), .B(KEYINPUT92), .Z(new_n760));
  XOR2_X1   g0560(.A(G355), .B(KEYINPUT93), .Z(new_n761));
  AOI22_X1  g0561(.A1(new_n760), .A2(new_n761), .B1(new_n625), .B2(new_n702), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n702), .A2(new_n409), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n764), .B1(new_n233), .B2(new_n255), .ZN(new_n765));
  INV_X1    g0565(.A(new_n249), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n765), .B1(new_n766), .B2(new_n255), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n758), .B1(new_n762), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n756), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n227), .A2(G190), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G179), .A2(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n417), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT95), .ZN(new_n774));
  XNOR2_X1  g0574(.A(KEYINPUT94), .B(KEYINPUT32), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n227), .A2(new_n311), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n380), .A2(G200), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n380), .A2(new_n468), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(new_n770), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n246), .A2(new_n779), .B1(new_n781), .B2(new_n357), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n227), .B1(new_n771), .B2(G190), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n777), .A2(new_n780), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n267), .B1(new_n783), .B2(new_n362), .C1(new_n784), .C2(new_n202), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n778), .A2(new_n770), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n782), .B(new_n785), .C1(G77), .C2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n468), .A2(G179), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT96), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n777), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G87), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n790), .A2(new_n770), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G107), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n776), .A2(new_n788), .A3(new_n793), .A4(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G326), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n429), .B1(new_n783), .B2(new_n550), .C1(new_n784), .C2(new_n798), .ZN(new_n799));
  XOR2_X1   g0599(.A(KEYINPUT33), .B(G317), .Z(new_n800));
  INV_X1    g0600(.A(G322), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n800), .A2(new_n781), .B1(new_n779), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G311), .ZN(new_n803));
  INV_X1    g0603(.A(G329), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n786), .A2(new_n803), .B1(new_n772), .B2(new_n804), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n799), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G283), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n806), .B1(new_n807), .B2(new_n794), .C1(new_n620), .C2(new_n791), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n769), .B1(new_n797), .B2(new_n808), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n768), .A2(new_n809), .A3(new_n749), .ZN(new_n810));
  INV_X1    g0610(.A(new_n755), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n810), .B1(new_n697), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n752), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(G396));
  OAI22_X1  g0614(.A1(new_n781), .A2(new_n807), .B1(new_n786), .B2(new_n625), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT97), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n816), .B1(new_n447), .B2(new_n794), .C1(new_n530), .C2(new_n791), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n783), .A2(new_n362), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n429), .B1(new_n784), .B2(new_n620), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n779), .A2(new_n550), .B1(new_n772), .B2(new_n803), .ZN(new_n820));
  NOR4_X1   g0620(.A1(new_n817), .A2(new_n818), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(KEYINPUT98), .ZN(new_n823));
  INV_X1    g0623(.A(new_n779), .ZN(new_n824));
  AOI22_X1  g0624(.A1(G143), .A2(new_n824), .B1(new_n787), .B2(G159), .ZN(new_n825));
  INV_X1    g0625(.A(G137), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n825), .B1(new_n826), .B2(new_n784), .C1(new_n315), .C2(new_n781), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT34), .ZN(new_n828));
  INV_X1    g0628(.A(new_n772), .ZN(new_n829));
  INV_X1    g0629(.A(new_n783), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G132), .A2(new_n829), .B1(new_n830), .B2(G58), .ZN(new_n831));
  AOI22_X1  g0631(.A1(G50), .A2(new_n792), .B1(new_n795), .B2(G68), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n828), .A2(new_n409), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT98), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n833), .B1(new_n821), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n756), .B1(new_n823), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n756), .A2(new_n753), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n749), .B1(new_n290), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n308), .A2(new_n682), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n312), .B1(new_n309), .B2(new_n685), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n839), .B1(new_n308), .B2(new_n840), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n836), .B(new_n838), .C1(new_n754), .C2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n682), .B1(new_n712), .B2(new_n719), .ZN(new_n843));
  AOI21_X1  g0643(.A(KEYINPUT99), .B1(new_n843), .B2(new_n841), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n843), .A2(new_n841), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n738), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n749), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n846), .A2(new_n738), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n842), .B1(new_n848), .B2(new_n849), .ZN(G384));
  NOR2_X1   g0650(.A1(new_n742), .A2(new_n287), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT102), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n464), .A2(new_n453), .ZN(new_n853));
  INV_X1    g0653(.A(new_n680), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n464), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n853), .A2(new_n855), .A3(new_n471), .ZN(new_n856));
  XNOR2_X1  g0656(.A(KEYINPUT100), .B(KEYINPUT37), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n853), .A2(new_n855), .A3(new_n471), .A4(new_n857), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n855), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n476), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  XOR2_X1   g0664(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n865));
  NAND2_X1  g0665(.A1(new_n457), .A2(new_n458), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n427), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n390), .B1(new_n426), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n471), .B1(new_n868), .B2(new_n680), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n868), .A2(new_n454), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT37), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n425), .A2(KEYINPUT16), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n456), .B1(new_n460), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n854), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n860), .A2(new_n871), .B1(new_n476), .B2(new_n875), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n864), .A2(new_n865), .B1(new_n876), .B2(KEYINPUT38), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n360), .A2(new_n682), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n383), .A2(new_n386), .A3(new_n878), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n360), .B(new_n682), .C1(new_n381), .C2(new_n382), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n881), .A2(new_n841), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n737), .A2(new_n882), .A3(KEYINPUT40), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n852), .B1(new_n877), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n881), .A2(new_n841), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n732), .A2(KEYINPUT31), .A3(new_n682), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT31), .B1(new_n732), .B2(new_n682), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n885), .B1(new_n888), .B2(new_n722), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n871), .A2(new_n860), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n476), .A2(new_n875), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n890), .A2(new_n891), .A3(KEYINPUT38), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT38), .B1(new_n890), .B2(new_n891), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n889), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT40), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n890), .A2(new_n891), .A3(KEYINPUT38), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n859), .A2(new_n860), .B1(new_n476), .B2(new_n862), .ZN(new_n898));
  INV_X1    g0698(.A(new_n865), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n900), .A2(KEYINPUT102), .A3(KEYINPUT40), .A4(new_n889), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n884), .A2(new_n896), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n480), .A2(new_n737), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n902), .A2(new_n903), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n904), .A2(G330), .A3(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT39), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n899), .B1(new_n861), .B2(new_n863), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n907), .B1(new_n892), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT38), .ZN(new_n910));
  INV_X1    g0710(.A(new_n891), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n853), .A2(new_n855), .A3(new_n471), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n873), .A2(new_n453), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n874), .A2(new_n913), .A3(new_n471), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n912), .A2(new_n857), .B1(new_n914), .B2(KEYINPUT37), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n910), .B1(new_n911), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n916), .A2(KEYINPUT39), .A3(new_n897), .ZN(new_n917));
  INV_X1    g0717(.A(new_n383), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n685), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n909), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n672), .A2(new_n854), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n916), .A2(new_n897), .ZN(new_n923));
  INV_X1    g0723(.A(new_n881), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n685), .B(new_n841), .C1(new_n659), .C2(new_n668), .ZN(new_n925));
  INV_X1    g0725(.A(new_n839), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n922), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n921), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n480), .B1(new_n718), .B2(new_n720), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n675), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n929), .B(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n851), .B1(new_n906), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n932), .B2(new_n906), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n528), .A2(KEYINPUT35), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n528), .A2(KEYINPUT35), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n935), .A2(G116), .A3(new_n228), .A4(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT36), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n415), .A2(G77), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n939), .A2(new_n232), .B1(G50), .B2(new_n357), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n940), .A2(G1), .A3(new_n353), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n934), .A2(new_n938), .A3(new_n941), .ZN(G367));
  OAI21_X1  g0742(.A(new_n535), .B1(new_n532), .B2(new_n685), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n715), .A2(new_n682), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n691), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n527), .B1(new_n943), .B2(new_n661), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n946), .A2(KEYINPUT42), .B1(new_n685), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(KEYINPUT42), .B2(new_n946), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n597), .A2(new_n598), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n682), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n653), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n593), .B2(new_n951), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT43), .B1(new_n953), .B2(KEYINPUT103), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(KEYINPUT103), .B2(new_n953), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n949), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n949), .B2(new_n956), .ZN(new_n958));
  INV_X1    g0758(.A(new_n945), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n958), .B1(new_n700), .B2(new_n959), .ZN(new_n960));
  OR3_X1    g0760(.A1(new_n958), .A2(new_n700), .A3(new_n959), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n703), .B(KEYINPUT41), .Z(new_n962));
  NOR3_X1   g0762(.A1(new_n691), .A2(new_n692), .A3(new_n959), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT45), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT44), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n693), .B2(new_n945), .ZN(new_n966));
  OAI211_X1 g0766(.A(KEYINPUT44), .B(new_n959), .C1(new_n691), .C2(new_n692), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n964), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT104), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n700), .ZN(new_n972));
  INV_X1    g0772(.A(new_n700), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n969), .A2(new_n970), .A3(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n694), .A2(new_n683), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n975), .A2(new_n691), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(new_n699), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n977), .A2(new_n739), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n972), .A2(new_n974), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n962), .B1(new_n979), .B2(new_n740), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n960), .B(new_n961), .C1(new_n980), .C2(new_n746), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n757), .B1(new_n223), .B2(new_n303), .C1(new_n764), .C2(new_n243), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n750), .A2(new_n982), .ZN(new_n983));
  AOI22_X1  g0783(.A1(G58), .A2(new_n792), .B1(new_n795), .B2(G77), .ZN(new_n984));
  INV_X1    g0784(.A(new_n781), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G159), .A2(new_n985), .B1(new_n787), .B2(G50), .ZN(new_n986));
  AOI22_X1  g0786(.A1(G150), .A2(new_n824), .B1(new_n829), .B2(G137), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n783), .A2(new_n357), .ZN(new_n988));
  INV_X1    g0788(.A(new_n784), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n429), .B(new_n988), .C1(G143), .C2(new_n989), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n984), .A2(new_n986), .A3(new_n987), .A4(new_n990), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n550), .A2(new_n781), .B1(new_n779), .B2(new_n620), .ZN(new_n992));
  AOI22_X1  g0792(.A1(G283), .A2(new_n787), .B1(new_n829), .B2(G317), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n803), .B2(new_n784), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n992), .B(new_n994), .C1(G107), .C2(new_n830), .ZN(new_n995));
  INV_X1    g0795(.A(new_n409), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n795), .A2(G97), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n791), .A2(new_n625), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT46), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n991), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT47), .Z(new_n1002));
  OAI221_X1 g0802(.A(new_n983), .B1(new_n811), .B2(new_n953), .C1(new_n1002), .C2(new_n769), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n981), .A2(new_n1003), .ZN(G387));
  OAI21_X1  g0804(.A(new_n763), .B1(new_n240), .B2(new_n255), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n760), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1005), .B1(new_n1006), .B2(new_n705), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n297), .A2(G50), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1009), .A2(KEYINPUT50), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(KEYINPUT50), .ZN(new_n1011));
  AOI21_X1  g0811(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1010), .A2(new_n705), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n1007), .A2(new_n1013), .B1(new_n530), .B2(new_n702), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n750), .B1(new_n1014), .B2(new_n758), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n792), .A2(G294), .B1(G283), .B2(new_n830), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G317), .A2(new_n824), .B1(new_n787), .B2(G303), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1017), .B1(new_n803), .B2(new_n781), .C1(new_n801), .C2(new_n784), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT48), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1016), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n1019), .B2(new_n1018), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1021), .A2(KEYINPUT49), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n996), .B1(new_n798), .B2(new_n772), .C1(new_n794), .C2(new_n625), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(KEYINPUT49), .B2(new_n1021), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n781), .A2(new_n296), .B1(new_n772), .B2(new_n315), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n784), .A2(new_n417), .B1(new_n786), .B2(new_n357), .ZN(new_n1027));
  NOR3_X1   g0827(.A1(new_n996), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n792), .A2(G77), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1028), .A2(new_n997), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n830), .A2(new_n577), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n202), .B2(new_n779), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT105), .Z(new_n1033));
  OAI21_X1  g0833(.A(new_n1025), .B1(new_n1030), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1015), .B1(new_n1034), .B2(new_n756), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n689), .A2(new_n690), .A3(new_n755), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n746), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n978), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n703), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n977), .A2(new_n739), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1037), .B1(new_n1038), .B2(new_n977), .C1(new_n1040), .C2(new_n1041), .ZN(G393));
  NOR2_X1   g0842(.A1(new_n969), .A2(new_n973), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n700), .B1(new_n964), .B2(new_n968), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1039), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT109), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1047), .A2(new_n703), .A3(new_n979), .A4(new_n1048), .ZN(new_n1049));
  NOR3_X1   g0849(.A1(new_n1043), .A2(new_n1038), .A3(new_n1044), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n959), .A2(new_n755), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n763), .A2(new_n252), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1052), .B(new_n757), .C1(new_n362), .C2(new_n223), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n750), .A2(new_n1053), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT106), .Z(new_n1055));
  AOI22_X1  g0855(.A1(new_n792), .A2(new_n210), .B1(G143), .B2(new_n829), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT107), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n783), .A2(new_n290), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1058), .B(new_n996), .C1(G50), .C2(new_n985), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n297), .A2(new_n786), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n784), .A2(new_n315), .B1(new_n779), .B2(new_n417), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT51), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n794), .A2(new_n447), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1060), .B(new_n1063), .C1(new_n1062), .C2(new_n1061), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1057), .A2(new_n1059), .A3(new_n1064), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G317), .A2(new_n989), .B1(new_n824), .B2(G311), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(KEYINPUT108), .B(KEYINPUT52), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1066), .B(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n429), .B1(new_n772), .B2(new_n801), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n781), .A2(new_n620), .B1(new_n786), .B2(new_n550), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1069), .B(new_n1070), .C1(G116), .C2(new_n830), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n792), .A2(G283), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1068), .A2(new_n796), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n769), .B1(new_n1065), .B2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1055), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1050), .B1(new_n1051), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1049), .A2(new_n1076), .ZN(G390));
  INV_X1    g0877(.A(G330), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n888), .B2(new_n722), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n480), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n930), .A2(new_n675), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n839), .B1(new_n843), .B2(new_n841), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n881), .B1(new_n1079), .B2(new_n841), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n738), .A2(new_n885), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1083), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n841), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n924), .B1(new_n738), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1079), .A2(new_n882), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n840), .A2(new_n308), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n717), .A2(new_n685), .A3(new_n1090), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1088), .A2(new_n1089), .A3(new_n926), .A4(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1081), .B1(new_n1086), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n909), .A2(new_n917), .ZN(new_n1095));
  OAI21_X1  g0895(.A(KEYINPUT110), .B1(new_n927), .B2(new_n920), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT110), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1097), .B(new_n919), .C1(new_n1082), .C2(new_n924), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1095), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1091), .A2(new_n926), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n919), .B(new_n900), .C1(new_n1100), .C2(new_n924), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1099), .A2(new_n1101), .A3(new_n1089), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1089), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1094), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n1085), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1107), .A2(new_n1102), .A3(new_n1093), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1105), .A2(new_n1108), .A3(new_n703), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n795), .A2(G68), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n784), .A2(new_n807), .B1(new_n779), .B2(new_n625), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n786), .A2(new_n362), .B1(new_n772), .B2(new_n550), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n267), .B(new_n1058), .C1(G107), .C2(new_n985), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n793), .A2(new_n1110), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n792), .A2(G150), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT53), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n267), .B1(new_n783), .B2(new_n417), .C1(new_n826), .C2(new_n781), .ZN(new_n1118));
  INV_X1    g0918(.A(G128), .ZN(new_n1119));
  INV_X1    g0919(.A(G132), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n784), .A2(new_n1119), .B1(new_n779), .B2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(KEYINPUT54), .B(G143), .ZN(new_n1122));
  INV_X1    g0922(.A(G125), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n786), .A2(new_n1122), .B1(new_n772), .B2(new_n1123), .ZN(new_n1124));
  NOR3_X1   g0924(.A1(new_n1118), .A2(new_n1121), .A3(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n202), .B2(new_n794), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1115), .B1(new_n1117), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT112), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n769), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n1128), .B2(new_n1127), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n837), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1130), .B(new_n750), .C1(new_n388), .C2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g0932(.A(new_n1132), .B(KEYINPUT113), .Z(new_n1133));
  INV_X1    g0933(.A(new_n1095), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1133), .B1(new_n1134), .B2(new_n754), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1107), .A2(new_n746), .A3(new_n1102), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1136), .A2(KEYINPUT111), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1136), .A2(KEYINPUT111), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1109), .B(new_n1135), .C1(new_n1137), .C2(new_n1138), .ZN(G378));
  NAND4_X1  g0939(.A1(new_n884), .A2(new_n896), .A3(G330), .A4(new_n901), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT116), .ZN(new_n1141));
  XOR2_X1   g0941(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1142));
  NAND2_X1  g0942(.A1(new_n320), .A2(new_n854), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n347), .A2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n347), .A2(new_n1143), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n1144), .A2(new_n1145), .A3(KEYINPUT115), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(KEYINPUT115), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1142), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1148), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1142), .ZN(new_n1151));
  NOR3_X1   g0951(.A1(new_n1150), .A2(new_n1151), .A3(new_n1146), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1141), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1151), .B1(new_n1150), .B2(new_n1146), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1147), .A2(new_n1142), .A3(new_n1148), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1154), .A2(new_n1155), .A3(KEYINPUT116), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  AND2_X1   g0957(.A1(new_n1140), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1153), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1140), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n929), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT117), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1140), .A2(new_n1157), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n929), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1163), .B(new_n1164), .C1(new_n1140), .C2(new_n1159), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1161), .A2(new_n1162), .A3(new_n1165), .ZN(new_n1166));
  OAI211_X1 g0966(.A(KEYINPUT117), .B(new_n929), .C1(new_n1158), .C2(new_n1160), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n930), .A2(new_n675), .A3(new_n1080), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1108), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1166), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT57), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1171), .B1(new_n1161), .B2(new_n1165), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n704), .B1(new_n1173), .B2(new_n1169), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1166), .A2(new_n746), .A3(new_n1167), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n781), .A2(new_n362), .B1(new_n786), .B2(new_n303), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT114), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1178), .B(new_n1029), .C1(new_n246), .C2(new_n794), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n996), .A2(new_n254), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n989), .A2(G116), .B1(new_n829), .B2(G283), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n530), .B2(new_n779), .ZN(new_n1182));
  NOR4_X1   g0982(.A1(new_n1179), .A2(new_n988), .A3(new_n1180), .A4(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(KEYINPUT58), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1180), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n781), .A2(new_n1120), .B1(new_n786), .B2(new_n826), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n784), .A2(new_n1123), .B1(new_n779), .B2(new_n1119), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1187), .B(new_n1188), .C1(G150), .C2(new_n830), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n791), .B2(new_n1122), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n795), .A2(G159), .ZN(new_n1193));
  AOI211_X1 g0993(.A(G33), .B(G41), .C1(new_n829), .C2(G124), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1186), .B1(KEYINPUT58), .B2(new_n1183), .C1(new_n1191), .C2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(new_n756), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n749), .B1(new_n202), .B2(new_n837), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1197), .B(new_n1198), .C1(new_n1199), .C2(new_n754), .ZN(new_n1200));
  AND2_X1   g1000(.A1(new_n1176), .A2(new_n1200), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1175), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(G375));
  OAI22_X1  g1003(.A1(new_n781), .A2(new_n625), .B1(new_n786), .B2(new_n530), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT118), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n429), .B1(new_n772), .B2(new_n620), .C1(new_n784), .C2(new_n550), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n795), .B2(G77), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1205), .B(new_n1207), .C1(new_n362), .C2(new_n791), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1031), .B1(new_n807), .B2(new_n779), .ZN(new_n1209));
  XOR2_X1   g1009(.A(new_n1209), .B(KEYINPUT119), .Z(new_n1210));
  NOR2_X1   g1010(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1212), .A2(KEYINPUT120), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n996), .B1(new_n795), .B2(G58), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n784), .A2(new_n1120), .B1(new_n786), .B2(new_n315), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G128), .B2(new_n829), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n826), .A2(new_n779), .B1(new_n781), .B2(new_n1122), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G50), .B2(new_n830), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n792), .A2(G159), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1214), .A2(new_n1216), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT120), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1220), .B1(new_n1211), .B2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n756), .B1(new_n1213), .B2(new_n1222), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1223), .B(new_n750), .C1(G68), .C2(new_n1131), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n924), .B2(new_n753), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1086), .A2(new_n1092), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1225), .B1(new_n1226), .B2(new_n746), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1093), .A2(new_n962), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1081), .A2(new_n1086), .A3(new_n1092), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1227), .B1(new_n1228), .B2(new_n1230), .ZN(G381));
  NAND2_X1  g1031(.A1(G378), .A2(KEYINPUT121), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1136), .B(KEYINPUT111), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT121), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1233), .A2(new_n1234), .A3(new_n1109), .A4(new_n1135), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1202), .A2(new_n1232), .A3(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(G390), .ZN(new_n1237));
  NOR4_X1   g1037(.A1(G393), .A2(G396), .A3(G384), .A4(G381), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1236), .A2(new_n1239), .A3(G387), .ZN(new_n1240));
  XOR2_X1   g1040(.A(new_n1240), .B(KEYINPUT122), .Z(G407));
  OAI211_X1 g1041(.A(G407), .B(G213), .C1(G343), .C2(new_n1236), .ZN(G409));
  AOI21_X1  g1042(.A(G390), .B1(new_n981), .B2(new_n1003), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(G393), .B(new_n813), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(G390), .A2(new_n981), .A3(new_n1003), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1245), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1246), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1248), .B1(new_n1249), .B2(new_n1243), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1175), .A2(G378), .A3(new_n1201), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1200), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1161), .A2(new_n1165), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1253), .B1(new_n1254), .B2(new_n746), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n1170), .B2(new_n962), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1232), .A2(new_n1235), .A3(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1252), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(G213), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1259), .A2(G343), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT126), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT125), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(new_n1226), .B2(new_n1168), .ZN(new_n1268));
  OAI21_X1  g1068(.A(KEYINPUT124), .B1(new_n1268), .B2(new_n1230), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT124), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1270), .B(new_n1229), .C1(new_n1093), .C2(new_n1267), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT60), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n703), .B1(new_n1229), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1265), .B1(new_n1272), .B2(new_n1275), .ZN(new_n1276));
  AOI211_X1 g1076(.A(KEYINPUT125), .B(new_n1274), .C1(new_n1269), .C2(new_n1271), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1227), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(new_n1278), .B(G384), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(KEYINPUT62), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT127), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1258), .A2(KEYINPUT126), .A3(new_n1261), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1264), .A2(new_n1281), .A3(new_n1282), .A4(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT61), .ZN(new_n1285));
  INV_X1    g1085(.A(G2897), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1261), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1279), .A2(new_n1287), .ZN(new_n1288));
  OR2_X1    g1088(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1289));
  AOI21_X1  g1089(.A(G384), .B1(new_n1289), .B2(new_n1227), .ZN(new_n1290));
  OAI211_X1 g1090(.A(G384), .B(new_n1227), .C1(new_n1276), .C2(new_n1277), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  OAI22_X1  g1092(.A1(new_n1290), .A2(new_n1292), .B1(new_n1286), .B2(new_n1261), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1288), .A2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT126), .B1(new_n1258), .B2(new_n1261), .ZN(new_n1295));
  AOI211_X1 g1095(.A(new_n1263), .B(new_n1260), .C1(new_n1252), .C2(new_n1257), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1294), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1284), .A2(new_n1285), .A3(new_n1297), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1295), .A2(new_n1296), .A3(new_n1280), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1258), .A2(new_n1261), .A3(new_n1279), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT62), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(KEYINPUT127), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1299), .A2(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1251), .B1(new_n1298), .B2(new_n1304), .ZN(new_n1305));
  AND2_X1   g1105(.A1(new_n1294), .A2(new_n1262), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT63), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1300), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1264), .A2(KEYINPUT63), .A3(new_n1283), .A4(new_n1279), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1251), .A2(KEYINPUT61), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1308), .A2(new_n1309), .A3(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1305), .A2(new_n1311), .ZN(G405));
  NAND2_X1  g1112(.A1(new_n1232), .A2(new_n1235), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1202), .A2(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1314), .B1(G378), .B2(new_n1202), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1279), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1319));
  OR3_X1    g1119(.A1(new_n1318), .A2(new_n1251), .A3(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1251), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(G402));
endmodule


