//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT65), .B1(new_n188), .B2(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n188), .A2(KEYINPUT65), .A3(G143), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT67), .B(G128), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT1), .B1(new_n194), .B2(G146), .ZN(new_n195));
  AOI22_X1  g009(.A1(new_n191), .A2(new_n192), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(G146), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n190), .A2(new_n197), .A3(new_n198), .A4(G128), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n187), .B1(new_n196), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT11), .ZN(new_n202));
  INV_X1    g016(.A(G134), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(G137), .ZN(new_n204));
  INV_X1    g018(.A(G137), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(KEYINPUT11), .A3(G134), .ZN(new_n206));
  INV_X1    g020(.A(G131), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n203), .A2(G137), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n204), .A2(new_n206), .A3(new_n207), .A4(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n203), .A2(G137), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n205), .A2(G134), .ZN(new_n211));
  OAI21_X1  g025(.A(G131), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n188), .A2(KEYINPUT65), .A3(G143), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n214), .B1(new_n190), .B2(new_n189), .ZN(new_n215));
  AND2_X1   g029(.A1(KEYINPUT67), .A2(G128), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(KEYINPUT67), .A2(G128), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  AOI22_X1  g033(.A1(new_n217), .A2(new_n219), .B1(KEYINPUT1), .B2(new_n190), .ZN(new_n220));
  OAI211_X1 g034(.A(KEYINPUT70), .B(new_n199), .C1(new_n215), .C2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n201), .A2(new_n213), .A3(new_n221), .ZN(new_n222));
  XOR2_X1   g036(.A(KEYINPUT2), .B(G113), .Z(new_n223));
  INV_X1    g037(.A(G119), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G116), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n226));
  INV_X1    g040(.A(G116), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(KEYINPUT68), .A2(G116), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(G119), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n223), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n223), .A2(new_n230), .A3(new_n225), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT69), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n223), .A2(new_n230), .A3(KEYINPUT69), .A4(new_n225), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n231), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n204), .A2(new_n206), .A3(new_n208), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G131), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(KEYINPUT66), .A3(new_n209), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT65), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n240), .B1(new_n194), .B2(G146), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n194), .A2(G146), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n192), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT0), .ZN(new_n244));
  INV_X1    g058(.A(G128), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n244), .A2(new_n245), .A3(KEYINPUT64), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT64), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n248), .B1(KEYINPUT0), .B2(G128), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n246), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n190), .A2(new_n197), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n243), .A2(new_n250), .B1(new_n246), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n237), .A2(new_n253), .A3(G131), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n239), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n222), .A2(new_n236), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(KEYINPUT28), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(KEYINPUT71), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n222), .A2(new_n236), .A3(new_n260), .A4(new_n255), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n222), .A2(new_n255), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n234), .A2(new_n235), .ZN(new_n263));
  INV_X1    g077(.A(new_n231), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n259), .A2(new_n261), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n258), .B1(new_n267), .B2(KEYINPUT28), .ZN(new_n268));
  NOR2_X1   g082(.A1(G237), .A2(G953), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G210), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n270), .B(KEYINPUT27), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT26), .B(G101), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n271), .B(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT29), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(G902), .B1(new_n268), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n199), .B1(new_n215), .B2(new_n220), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n213), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n255), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n265), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT72), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n280), .A2(new_n265), .A3(new_n283), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n282), .A2(new_n259), .A3(new_n261), .A4(new_n284), .ZN(new_n285));
  AOI211_X1 g099(.A(new_n274), .B(new_n258), .C1(new_n285), .C2(KEYINPUT28), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT30), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n287), .B1(new_n222), .B2(new_n255), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n255), .A2(new_n287), .A3(new_n279), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n265), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n259), .A2(new_n261), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n274), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n275), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n277), .B1(new_n286), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G472), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n290), .A2(new_n259), .A3(new_n261), .A4(new_n273), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT31), .ZN(new_n298));
  INV_X1    g112(.A(new_n292), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT31), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n299), .A2(new_n300), .A3(new_n273), .A4(new_n290), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n258), .B1(new_n285), .B2(KEYINPUT28), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n298), .B(new_n301), .C1(new_n302), .C2(new_n273), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT32), .ZN(new_n304));
  NOR2_X1   g118(.A1(G472), .A2(G902), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n304), .B1(new_n303), .B2(new_n305), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n296), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n224), .A2(G128), .ZN(new_n309));
  AND2_X1   g123(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n310));
  NOR2_X1   g124(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n311));
  OAI22_X1  g125(.A1(new_n310), .A2(new_n311), .B1(new_n224), .B2(G128), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n216), .A2(new_n218), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G119), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT23), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n309), .B(new_n312), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n314), .A2(new_n309), .ZN(new_n317));
  XOR2_X1   g131(.A(KEYINPUT24), .B(G110), .Z(new_n318));
  AOI22_X1  g132(.A1(new_n316), .A2(G110), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G140), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G125), .ZN(new_n321));
  INV_X1    g135(.A(G125), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G140), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n321), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n322), .A2(KEYINPUT74), .A3(G140), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(KEYINPUT16), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT16), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n321), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n188), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n327), .A2(new_n329), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(G146), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n319), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  OAI22_X1  g147(.A1(new_n316), .A2(G110), .B1(new_n317), .B2(new_n318), .ZN(new_n334));
  INV_X1    g148(.A(new_n330), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n321), .A2(new_n323), .A3(new_n188), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n334), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT22), .B(G137), .ZN(new_n339));
  INV_X1    g153(.A(G953), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(G221), .A3(G234), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n339), .B(new_n341), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n333), .A2(new_n338), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n342), .B1(new_n333), .B2(new_n338), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G902), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(KEYINPUT25), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n333), .A2(new_n338), .ZN(new_n348));
  INV_X1    g162(.A(new_n342), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n333), .A2(new_n338), .A3(new_n342), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n346), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT25), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n347), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G217), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(G234), .B2(new_n346), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n357), .A2(G902), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n345), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n358), .A2(KEYINPUT75), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT75), .ZN(new_n362));
  INV_X1    g176(.A(new_n357), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n363), .B1(new_n347), .B2(new_n354), .ZN(new_n364));
  INV_X1    g178(.A(new_n360), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n362), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n308), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT9), .B(G234), .ZN(new_n369));
  OAI21_X1  g183(.A(G221), .B1(new_n369), .B2(G902), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n370), .B(KEYINPUT76), .ZN(new_n371));
  XOR2_X1   g185(.A(new_n371), .B(KEYINPUT77), .Z(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT78), .B(G101), .ZN(new_n374));
  INV_X1    g188(.A(G104), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT3), .B1(new_n375), .B2(G107), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT3), .ZN(new_n377));
  INV_X1    g191(.A(G107), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(G104), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n375), .A2(G107), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n374), .A2(new_n376), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n380), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n375), .A2(G107), .ZN(new_n383));
  OAI21_X1  g197(.A(G101), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n381), .A2(KEYINPUT10), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n201), .A2(new_n221), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n376), .A2(new_n379), .A3(new_n380), .ZN(new_n387));
  AOI22_X1  g201(.A1(new_n381), .A2(KEYINPUT4), .B1(G101), .B2(new_n387), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n387), .A2(KEYINPUT4), .A3(G101), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n252), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n239), .A2(new_n254), .ZN(new_n391));
  AOI22_X1  g205(.A1(new_n195), .A2(G128), .B1(new_n190), .B2(new_n197), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n381), .B(new_n384), .C1(new_n200), .C2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT10), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n386), .A2(new_n390), .A3(new_n391), .A4(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(G110), .B(G140), .ZN(new_n397));
  INV_X1    g211(.A(G227), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(G953), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n397), .B(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT80), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT79), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n239), .A2(new_n405), .A3(new_n254), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n381), .A2(new_n384), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n393), .B1(new_n407), .B2(new_n278), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT12), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n406), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n409), .B1(new_n406), .B2(new_n408), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n396), .A2(KEYINPUT80), .A3(new_n401), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n404), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n386), .A2(new_n395), .A3(new_n390), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(new_n254), .A3(new_n239), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n396), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n400), .ZN(new_n419));
  AOI211_X1 g233(.A(G469), .B(G902), .C1(new_n415), .C2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n406), .A2(new_n408), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT12), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n422), .A2(new_n396), .A3(new_n410), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n400), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n417), .A2(new_n396), .A3(new_n401), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(G469), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(G469), .A2(G902), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n373), .B1(new_n420), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT81), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g245(.A(KEYINPUT81), .B(new_n373), .C1(new_n420), .C2(new_n428), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n434));
  XNOR2_X1  g248(.A(G113), .B(G122), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(new_n375), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n325), .A2(new_n326), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT84), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n325), .A2(KEYINPUT84), .A3(new_n326), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(G146), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n337), .ZN(new_n442));
  INV_X1    g256(.A(G237), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(new_n340), .A3(G214), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n194), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n269), .A2(G143), .A3(G214), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(KEYINPUT18), .A2(G131), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n447), .B(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n442), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT86), .ZN(new_n451));
  INV_X1    g265(.A(new_n446), .ZN(new_n452));
  AOI21_X1  g266(.A(G143), .B1(new_n269), .B2(G214), .ZN(new_n453));
  OAI21_X1  g267(.A(G131), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT85), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT85), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n447), .A2(new_n456), .A3(G131), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n451), .B1(new_n458), .B2(KEYINPUT17), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT17), .ZN(new_n460));
  AOI211_X1 g274(.A(KEYINPUT86), .B(new_n460), .C1(new_n455), .C2(new_n457), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n327), .A2(new_n188), .A3(new_n329), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n445), .A2(new_n207), .A3(new_n446), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n455), .A2(new_n457), .A3(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n463), .B(new_n335), .C1(new_n465), .C2(KEYINPUT17), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n436), .B(new_n450), .C1(new_n462), .C2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n439), .A2(KEYINPUT19), .A3(new_n440), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT19), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n321), .A2(new_n323), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n335), .B(new_n465), .C1(new_n471), .C2(G146), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n450), .ZN(new_n473));
  INV_X1    g287(.A(new_n436), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n467), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(G475), .A2(G902), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n434), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n477), .ZN(new_n480));
  AOI211_X1 g294(.A(KEYINPUT20), .B(new_n480), .C1(new_n467), .C2(new_n475), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n450), .B1(new_n462), .B2(new_n466), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n474), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n467), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n346), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n479), .A2(new_n482), .B1(new_n486), .B2(G475), .ZN(new_n487));
  NOR3_X1   g301(.A1(new_n369), .A2(new_n356), .A3(G953), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n228), .A2(G122), .A3(new_n229), .ZN(new_n490));
  INV_X1    g304(.A(G122), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G116), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(new_n378), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT14), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n228), .A2(new_n494), .A3(G122), .A4(new_n229), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n496), .A2(KEYINPUT92), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(G107), .B1(new_n496), .B2(KEYINPUT92), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n493), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(KEYINPUT90), .B1(new_n193), .B2(new_n194), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT90), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n313), .A2(new_n502), .A3(G143), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT88), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n505), .B1(G128), .B2(new_n194), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n245), .A2(KEYINPUT88), .A3(G143), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n504), .A2(new_n203), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n502), .B1(new_n313), .B2(G143), .ZN(new_n511));
  NOR4_X1   g325(.A1(new_n216), .A2(new_n218), .A3(KEYINPUT90), .A4(new_n194), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(G134), .B1(new_n513), .B2(new_n508), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n500), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n516), .B1(new_n506), .B2(new_n507), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n505), .A2(new_n194), .A3(G128), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT88), .B1(new_n245), .B2(G143), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT13), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n520), .A2(KEYINPUT89), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n520), .A2(KEYINPUT89), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n518), .B(new_n519), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n517), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(G134), .B1(new_n513), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n510), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n490), .A2(new_n378), .A3(new_n492), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n378), .B1(new_n490), .B2(new_n492), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n527), .A2(new_n528), .A3(KEYINPUT87), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT87), .ZN(new_n530));
  AND2_X1   g344(.A1(KEYINPUT68), .A2(G116), .ZN(new_n531));
  NOR2_X1   g345(.A1(KEYINPUT68), .A2(G116), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n531), .A2(new_n532), .A3(new_n491), .ZN(new_n533));
  INV_X1    g347(.A(new_n492), .ZN(new_n534));
  OAI21_X1  g348(.A(G107), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n530), .B1(new_n535), .B2(new_n493), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n529), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT91), .B1(new_n526), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(KEYINPUT87), .B1(new_n527), .B2(new_n528), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n535), .A2(new_n530), .A3(new_n493), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT91), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n541), .A2(new_n542), .A3(new_n510), .A4(new_n525), .ZN(new_n543));
  AOI211_X1 g357(.A(new_n489), .B(new_n515), .C1(new_n538), .C2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n538), .A2(new_n543), .ZN(new_n545));
  INV_X1    g359(.A(new_n515), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n488), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n346), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT93), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT93), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n550), .B(new_n346), .C1(new_n544), .C2(new_n547), .ZN(new_n551));
  INV_X1    g365(.A(G478), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT94), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n553), .A2(KEYINPUT15), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(KEYINPUT15), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n552), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n549), .A2(new_n551), .A3(new_n557), .ZN(new_n558));
  OR2_X1    g372(.A1(new_n548), .A2(new_n557), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n487), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(G214), .B1(G237), .B2(G902), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(G210), .B1(G237), .B2(G902), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(G110), .B(G122), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n230), .A2(KEYINPUT5), .A3(new_n225), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n567), .B(G113), .C1(KEYINPUT5), .C2(new_n225), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n263), .A2(new_n407), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n388), .A2(new_n389), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(new_n236), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n566), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n569), .B(new_n565), .C1(new_n236), .C2(new_n571), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(new_n574), .A3(KEYINPUT6), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT6), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n576), .B(new_n566), .C1(new_n570), .C2(new_n572), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n278), .A2(G125), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n252), .A2(new_n322), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(KEYINPUT82), .B(G224), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n340), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n580), .B(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n575), .A2(new_n577), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n582), .A2(KEYINPUT7), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT83), .B1(new_n580), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT83), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n589), .B(new_n586), .C1(new_n578), .C2(new_n579), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n580), .A2(new_n587), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n565), .B(KEYINPUT8), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n407), .B1(new_n263), .B2(new_n568), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n593), .B1(new_n570), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n574), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n346), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n564), .B1(new_n585), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n597), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n599), .A2(new_n563), .A3(new_n584), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n562), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(G234), .A2(G237), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n602), .A2(G952), .A3(new_n340), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n602), .A2(G902), .A3(G953), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT21), .B(G898), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n601), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n560), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n368), .A2(new_n433), .A3(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(new_n610), .B(new_n374), .Z(G3));
  INV_X1    g425(.A(KEYINPUT95), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n515), .B1(new_n538), .B2(new_n543), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n612), .B1(new_n613), .B2(new_n488), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n614), .B(KEYINPUT33), .C1(new_n544), .C2(new_n547), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n517), .A2(new_n523), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n203), .B1(new_n616), .B2(new_n504), .ZN(new_n617));
  AOI211_X1 g431(.A(G134), .B(new_n508), .C1(new_n501), .C2(new_n503), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n542), .B1(new_n619), .B2(new_n541), .ZN(new_n620));
  INV_X1    g434(.A(new_n543), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n546), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n489), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n613), .A2(new_n488), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT33), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n623), .B(new_n624), .C1(new_n612), .C2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n615), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n552), .A2(G902), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(KEYINPUT96), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n549), .A2(new_n551), .A3(new_n552), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT96), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n627), .A2(new_n632), .A3(new_n628), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n608), .ZN(new_n635));
  AOI21_X1  g449(.A(G902), .B1(new_n484), .B2(new_n467), .ZN(new_n636));
  INV_X1    g450(.A(G475), .ZN(new_n637));
  OAI22_X1  g451(.A1(new_n478), .A2(new_n481), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n634), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(G472), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n640), .B1(new_n303), .B2(new_n346), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n305), .B2(new_n303), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n433), .A2(new_n642), .A3(new_n367), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT34), .B(G104), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  AND2_X1   g460(.A1(new_n642), .A2(new_n367), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n558), .A2(new_n559), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n648), .A2(new_n638), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n647), .A2(new_n433), .A3(new_n635), .A4(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT35), .B(G107), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G9));
  NAND2_X1  g466(.A1(new_n348), .A2(KEYINPUT97), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT97), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n333), .A2(new_n338), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n349), .A2(KEYINPUT36), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n653), .A2(new_n657), .A3(new_n655), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n659), .A2(new_n359), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(KEYINPUT98), .B1(new_n358), .B2(new_n661), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n659), .A2(new_n359), .A3(new_n660), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT98), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n364), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n609), .A2(new_n433), .A3(new_n642), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT37), .B(G110), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT99), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n667), .B(new_n669), .ZN(G12));
  AND3_X1   g484(.A1(new_n433), .A2(new_n308), .A3(new_n666), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n558), .A2(new_n559), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT100), .ZN(new_n673));
  INV_X1    g487(.A(G900), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n603), .B1(new_n604), .B2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n672), .A2(new_n673), .A3(new_n487), .A4(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n672), .A2(new_n487), .A3(new_n676), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT100), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n671), .A2(new_n601), .A3(new_n677), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G128), .ZN(G30));
  INV_X1    g495(.A(new_n433), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n675), .B(KEYINPUT39), .ZN(new_n683));
  OR2_X1    g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OR2_X1    g498(.A1(new_n684), .A2(KEYINPUT40), .ZN(new_n685));
  OR2_X1    g499(.A1(new_n306), .A2(new_n307), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n299), .A2(new_n290), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n273), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n688), .B1(new_n273), .B2(new_n267), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT101), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n346), .B1(new_n689), .B2(new_n690), .ZN(new_n692));
  OAI21_X1  g506(.A(G472), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n686), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n364), .A2(new_n663), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n585), .A2(new_n597), .A3(new_n564), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n563), .B1(new_n599), .B2(new_n584), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT38), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n672), .A2(new_n561), .A3(new_n638), .ZN(new_n702));
  NOR4_X1   g516(.A1(new_n695), .A2(new_n697), .A3(new_n701), .A4(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n684), .A2(KEYINPUT40), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n685), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT102), .B(G143), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G45));
  AND4_X1   g521(.A1(new_n308), .A2(new_n433), .A3(new_n666), .A4(new_n601), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n633), .A2(new_n631), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n632), .B1(new_n627), .B2(new_n628), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n638), .B(new_n676), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(KEYINPUT103), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT103), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n634), .A2(new_n713), .A3(new_n638), .A4(new_n676), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n708), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G146), .ZN(G48));
  AND3_X1   g530(.A1(new_n404), .A2(new_n413), .A3(new_n414), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n401), .B1(new_n417), .B2(new_n396), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(G469), .B1(new_n719), .B2(G902), .ZN(new_n720));
  INV_X1    g534(.A(G469), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n721), .B(new_n346), .C1(new_n717), .C2(new_n718), .ZN(new_n722));
  INV_X1    g536(.A(new_n371), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n720), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n308), .A2(new_n367), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n639), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g541(.A(KEYINPUT41), .B(G113), .Z(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G15));
  NOR4_X1   g543(.A1(new_n726), .A2(new_n608), .A3(new_n648), .A4(new_n638), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(new_n227), .ZN(G18));
  AND4_X1   g545(.A1(new_n607), .A2(new_n487), .A3(new_n558), .A4(new_n559), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n561), .B1(new_n698), .B2(new_n699), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n724), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n732), .A2(new_n308), .A3(new_n734), .A4(new_n666), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G119), .ZN(G21));
  NAND2_X1  g550(.A1(new_n638), .A2(new_n561), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n737), .B1(new_n559), .B2(new_n558), .ZN(new_n738));
  INV_X1    g552(.A(new_n305), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n298), .A2(new_n301), .ZN(new_n740));
  OR2_X1    g554(.A1(new_n268), .A2(new_n273), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n358), .A2(new_n360), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n641), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n700), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n724), .A2(new_n606), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n738), .A2(new_n744), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G122), .ZN(G24));
  NAND2_X1  g562(.A1(new_n725), .A2(new_n601), .ZN(new_n749));
  INV_X1    g563(.A(new_n641), .ZN(new_n750));
  INV_X1    g564(.A(new_n742), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n751), .A3(new_n697), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n712), .A2(new_n714), .A3(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G125), .ZN(G27));
  NAND2_X1  g569(.A1(new_n712), .A2(new_n714), .ZN(new_n756));
  INV_X1    g570(.A(new_n743), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n308), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g572(.A(new_n427), .B(KEYINPUT104), .Z(new_n759));
  NAND2_X1  g573(.A1(new_n426), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n371), .B1(new_n761), .B2(new_n722), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT105), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n598), .A2(new_n600), .A3(new_n561), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n723), .B1(new_n420), .B2(new_n760), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n765), .B1(new_n766), .B2(KEYINPUT105), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n758), .A2(new_n764), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT42), .B1(new_n756), .B2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n308), .A2(new_n367), .A3(new_n767), .A4(new_n764), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT42), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n771), .A2(new_n712), .A3(new_n772), .A4(new_n714), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(new_n207), .ZN(G33));
  INV_X1    g589(.A(KEYINPUT106), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n771), .A2(new_n776), .A3(new_n677), .A4(new_n679), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n679), .A2(new_n677), .ZN(new_n778));
  OAI21_X1  g592(.A(KEYINPUT106), .B1(new_n778), .B2(new_n770), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G134), .ZN(G36));
  NAND2_X1  g595(.A1(new_n634), .A2(new_n487), .ZN(new_n782));
  XOR2_X1   g596(.A(new_n782), .B(KEYINPUT43), .Z(new_n783));
  NOR2_X1   g597(.A1(new_n642), .A2(new_n696), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT44), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n424), .A2(KEYINPUT45), .A3(new_n425), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT45), .B1(new_n424), .B2(new_n425), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n786), .A2(new_n787), .A3(new_n721), .ZN(new_n788));
  INV_X1    g602(.A(new_n759), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n790), .A2(KEYINPUT46), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n722), .B1(new_n790), .B2(KEYINPUT46), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n723), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR4_X1   g607(.A1(new_n785), .A2(new_n683), .A3(new_n765), .A4(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n783), .A2(KEYINPUT44), .A3(new_n784), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G137), .ZN(G39));
  INV_X1    g611(.A(new_n756), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n308), .A2(new_n367), .A3(new_n765), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(KEYINPUT107), .A3(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT47), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n793), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n793), .A2(new_n801), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT107), .B1(new_n798), .B2(new_n799), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(new_n320), .ZN(G42));
  INV_X1    g622(.A(new_n765), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n720), .A2(new_n722), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n811), .A2(KEYINPUT115), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(KEYINPUT115), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n812), .A2(new_n372), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n809), .B1(new_n804), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n783), .A2(new_n603), .A3(new_n744), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n701), .A2(new_n562), .A3(new_n725), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n820), .B(KEYINPUT117), .Z(new_n821));
  OR3_X1    g635(.A1(new_n816), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n819), .B1(new_n816), .B2(new_n821), .ZN(new_n823));
  AOI22_X1  g637(.A1(KEYINPUT116), .A2(new_n818), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n724), .A2(new_n765), .ZN(new_n825));
  AND4_X1   g639(.A1(new_n367), .A2(new_n695), .A3(new_n603), .A4(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n634), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n826), .A2(new_n487), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n783), .A2(new_n603), .A3(new_n825), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n828), .B1(new_n829), .B2(new_n752), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n830), .B1(new_n817), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT51), .B1(new_n824), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(G952), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n827), .A2(new_n487), .ZN(new_n835));
  AOI211_X1 g649(.A(new_n834), .B(G953), .C1(new_n826), .C2(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n836), .B1(new_n749), .B2(new_n816), .ZN(new_n837));
  INV_X1    g651(.A(new_n758), .ZN(new_n838));
  OR3_X1    g652(.A1(new_n829), .A2(KEYINPUT48), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT48), .B1(new_n829), .B2(new_n838), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n837), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n822), .A2(new_n823), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n829), .A2(new_n752), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n818), .A2(new_n843), .A3(KEYINPUT51), .A4(new_n828), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n841), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n833), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n735), .B(new_n747), .C1(new_n639), .C2(new_n726), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(new_n730), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n849), .A2(new_n769), .A3(new_n773), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n650), .A2(new_n667), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT108), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n610), .B(new_n852), .C1(new_n639), .C2(new_n643), .ZN(new_n853));
  INV_X1    g667(.A(new_n560), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n854), .A2(new_n635), .A3(new_n433), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n308), .A2(new_n367), .ZN(new_n856));
  OAI22_X1  g670(.A1(new_n639), .A2(new_n643), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(KEYINPUT108), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n851), .A2(new_n853), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n767), .A2(new_n764), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n860), .A2(new_n752), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n712), .A2(new_n861), .A3(new_n714), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT111), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT111), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n712), .A2(new_n861), .A3(new_n714), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n598), .A2(new_n600), .A3(new_n561), .A4(new_n676), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT109), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n648), .A2(new_n868), .A3(new_n869), .A4(new_n487), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT109), .B1(new_n560), .B2(new_n867), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n433), .A2(new_n308), .A3(new_n666), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT110), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT110), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n671), .A2(new_n875), .A3(new_n870), .A4(new_n871), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n777), .A2(new_n779), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n850), .A2(new_n859), .A3(new_n866), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n696), .A2(new_n676), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT112), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n702), .A2(new_n700), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n880), .A2(new_n881), .A3(new_n694), .A4(new_n762), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n715), .A2(new_n882), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n680), .A2(new_n754), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT52), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n715), .A2(new_n680), .A3(new_n754), .A4(new_n882), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT52), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n878), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n883), .A2(new_n884), .A3(KEYINPUT52), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n886), .A2(new_n887), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n891), .A2(KEYINPUT113), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT113), .B1(new_n891), .B2(new_n892), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n878), .A2(KEYINPUT53), .ZN(new_n897));
  OAI221_X1 g711(.A(KEYINPUT54), .B1(new_n847), .B2(new_n890), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n877), .A2(new_n866), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n849), .A2(new_n769), .A3(KEYINPUT53), .A4(new_n773), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n851), .A2(new_n853), .A3(new_n858), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT113), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n903), .B1(new_n885), .B2(new_n888), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n891), .A2(KEYINPUT113), .A3(new_n892), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n902), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT114), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT54), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n847), .B1(new_n878), .B2(new_n889), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT114), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n902), .A2(new_n904), .A3(new_n910), .A4(new_n905), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n907), .A2(new_n908), .A3(new_n909), .A4(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n846), .A2(new_n898), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n834), .A2(new_n340), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n743), .A2(new_n372), .A3(new_n562), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n701), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n917), .B1(KEYINPUT49), .B2(new_n810), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n782), .A2(new_n694), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n918), .B(new_n919), .C1(KEYINPUT49), .C2(new_n810), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n915), .A2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT118), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n915), .A2(KEYINPUT118), .A3(new_n920), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(G75));
  NAND3_X1  g739(.A1(new_n907), .A2(new_n909), .A3(new_n911), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n926), .A2(G210), .A3(G902), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n927), .A2(KEYINPUT119), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(KEYINPUT119), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n575), .A2(new_n577), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(new_n583), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT55), .Z(new_n932));
  NOR2_X1   g746(.A1(new_n932), .A2(KEYINPUT56), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n928), .A2(new_n929), .A3(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n340), .A2(G952), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT56), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n927), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n935), .B1(new_n937), .B2(new_n932), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n934), .A2(new_n938), .ZN(G51));
  NAND3_X1  g753(.A1(new_n926), .A2(G902), .A3(new_n788), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n910), .B1(new_n895), .B2(new_n902), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n911), .A2(new_n909), .ZN(new_n943));
  OAI21_X1  g757(.A(KEYINPUT54), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n912), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n759), .B(KEYINPUT57), .Z(new_n946));
  AOI21_X1  g760(.A(new_n719), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n941), .B1(new_n947), .B2(KEYINPUT120), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT120), .ZN(new_n949));
  INV_X1    g763(.A(new_n946), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n950), .B1(new_n944), .B2(new_n912), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n949), .B1(new_n951), .B2(new_n719), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n935), .B1(new_n948), .B2(new_n952), .ZN(G54));
  INV_X1    g767(.A(new_n476), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n926), .A2(G902), .ZN(new_n955));
  NAND2_X1  g769(.A1(KEYINPUT58), .A2(G475), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n935), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n955), .A2(new_n954), .A3(new_n956), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(G60));
  NAND2_X1  g775(.A1(G478), .A2(G902), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT59), .Z(new_n963));
  AOI21_X1  g777(.A(new_n963), .B1(new_n898), .B2(new_n912), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n958), .B1(new_n964), .B2(new_n627), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n963), .B1(new_n615), .B2(new_n626), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n945), .A2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT121), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n945), .A2(KEYINPUT121), .A3(new_n966), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n965), .B1(new_n969), .B2(new_n970), .ZN(G63));
  NAND2_X1  g785(.A1(G217), .A2(G902), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT60), .Z(new_n973));
  NAND4_X1  g787(.A1(new_n926), .A2(new_n660), .A3(new_n659), .A4(new_n973), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n926), .A2(new_n973), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n958), .B(new_n974), .C1(new_n975), .C2(new_n345), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT61), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n976), .B(new_n977), .ZN(G66));
  INV_X1    g792(.A(new_n605), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n340), .B1(new_n979), .B2(new_n581), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n859), .A2(new_n849), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n980), .B1(new_n981), .B2(new_n340), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n930), .B1(G898), .B2(new_n340), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT122), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n982), .B(new_n984), .ZN(G69));
  OAI211_X1 g799(.A(new_n368), .B(new_n809), .C1(new_n835), .C2(new_n649), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n986), .A2(new_n684), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n987), .B1(new_n794), .B2(new_n795), .ZN(new_n988));
  INV_X1    g802(.A(new_n807), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n884), .A2(new_n715), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n705), .ZN(new_n991));
  OR2_X1    g805(.A1(new_n991), .A2(KEYINPUT62), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(KEYINPUT62), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n988), .A2(new_n989), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n340), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n471), .B(KEYINPUT123), .Z(new_n996));
  NOR2_X1   g810(.A1(new_n288), .A2(new_n289), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n340), .A2(G900), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n793), .A2(new_n683), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n1001), .A2(new_n881), .A3(new_n758), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT126), .ZN(new_n1003));
  INV_X1    g817(.A(new_n780), .ZN(new_n1004));
  NOR4_X1   g818(.A1(new_n807), .A2(new_n1003), .A3(new_n774), .A4(new_n1004), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n796), .A2(KEYINPUT125), .A3(new_n990), .ZN(new_n1006));
  AOI21_X1  g820(.A(KEYINPUT125), .B1(new_n796), .B2(new_n990), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1000), .B1(new_n1008), .B2(new_n340), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n999), .B1(new_n1009), .B2(new_n998), .ZN(new_n1010));
  OAI21_X1  g824(.A(G953), .B1(new_n398), .B2(new_n674), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1011), .B(KEYINPUT124), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1010), .B(new_n1012), .ZN(G72));
  NAND2_X1  g827(.A1(G472), .A2(G902), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1014), .B(KEYINPUT63), .Z(new_n1015));
  OAI21_X1  g829(.A(new_n1015), .B1(new_n994), .B2(new_n981), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT127), .ZN(new_n1017));
  OR2_X1    g831(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1018), .A2(new_n273), .A3(new_n687), .A4(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1015), .B1(new_n1008), .B2(new_n981), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n687), .A2(new_n273), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n935), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1015), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1024), .B1(new_n293), .B2(new_n297), .ZN(new_n1025));
  OAI221_X1 g839(.A(new_n1025), .B1(new_n847), .B2(new_n890), .C1(new_n896), .C2(new_n897), .ZN(new_n1026));
  AND3_X1   g840(.A1(new_n1020), .A2(new_n1023), .A3(new_n1026), .ZN(G57));
endmodule


