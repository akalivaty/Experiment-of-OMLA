//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 1 1 1 0 1 1 0 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1124,
    new_n1125;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT64), .Z(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n458), .A2(KEYINPUT65), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(G567), .B2(new_n455), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(KEYINPUT65), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G137), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT3), .B(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n472), .A2(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n467), .A2(G136), .ZN(new_n479));
  XOR2_X1   g054(.A(new_n479), .B(KEYINPUT66), .Z(new_n480));
  NOR2_X1   g055(.A1(new_n466), .A2(new_n473), .ZN(new_n481));
  NOR2_X1   g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT67), .ZN(new_n483));
  INV_X1    g058(.A(G112), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n469), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  AOI22_X1  g060(.A1(G124), .A2(new_n481), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n480), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n489), .B1(new_n490), .B2(G2105), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(new_n481), .B2(G126), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT68), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n497), .A2(new_n474), .A3(new_n498), .A4(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n464), .B2(new_n465), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n473), .A2(G138), .ZN(new_n505));
  INV_X1    g080(.A(new_n465), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n498), .B1(new_n508), .B2(new_n497), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n492), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(KEYINPUT71), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(KEYINPUT5), .A3(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT72), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n517), .A2(KEYINPUT72), .A3(new_n518), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n523), .A2(G88), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n518), .A2(G543), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n525), .A2(KEYINPUT70), .A3(G50), .ZN(new_n526));
  AOI21_X1  g101(.A(KEYINPUT70), .B1(new_n525), .B2(G50), .ZN(new_n527));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n526), .A2(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n524), .A2(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n518), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G51), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n514), .A2(new_n516), .ZN(new_n537));
  NAND2_X1  g112(.A1(G63), .A2(G651), .ZN(new_n538));
  OAI221_X1 g113(.A(new_n534), .B1(new_n535), .B2(new_n536), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n539), .B1(new_n523), .B2(G89), .ZN(G168));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G64), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n543), .A2(G651), .B1(G52), .B2(new_n525), .ZN(new_n544));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n521), .A2(new_n522), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT73), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n547), .B(new_n548), .ZN(G171));
  NAND2_X1  g124(.A1(new_n523), .A2(G81), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n517), .A2(G56), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n528), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(KEYINPUT74), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n553), .A2(KEYINPUT74), .B1(G43), .B2(new_n525), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n550), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  AND3_X1   g138(.A1(new_n525), .A2(new_n563), .A3(G53), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n563), .B1(new_n525), .B2(G53), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n517), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n566));
  OAI22_X1  g141(.A1(new_n564), .A2(new_n565), .B1(new_n528), .B2(new_n566), .ZN(new_n567));
  AND3_X1   g142(.A1(new_n521), .A2(G91), .A3(new_n522), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(G299));
  XNOR2_X1  g145(.A(new_n547), .B(KEYINPUT73), .ZN(G301));
  INV_X1    g146(.A(G168), .ZN(G286));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n573));
  AND3_X1   g148(.A1(new_n521), .A2(G87), .A3(new_n522), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n575));
  INV_X1    g150(.A(G49), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n576), .B2(new_n535), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n573), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n517), .A2(G74), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n579), .A2(G651), .B1(G49), .B2(new_n525), .ZN(new_n580));
  INV_X1    g155(.A(G87), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n580), .B(KEYINPUT75), .C1(new_n581), .C2(new_n546), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n578), .A2(new_n582), .ZN(G288));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n537), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n586), .A2(G651), .B1(G48), .B2(new_n525), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n521), .A2(G86), .A3(new_n522), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n528), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(KEYINPUT76), .ZN(new_n592));
  XOR2_X1   g167(.A(KEYINPUT77), .B(G47), .Z(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n535), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g169(.A(KEYINPUT78), .B(G85), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n546), .A2(new_n595), .B1(new_n591), .B2(KEYINPUT76), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G290));
  NAND3_X1  g173(.A1(new_n523), .A2(KEYINPUT10), .A3(G92), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  INV_X1    g175(.A(G92), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n546), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT79), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n537), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n607), .A2(G651), .B1(G54), .B2(new_n525), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g186(.A(new_n610), .B1(G868), .B2(G171), .ZN(G321));
  NAND2_X1  g187(.A1(G286), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n569), .ZN(G297));
  OAI21_X1  g189(.A(new_n613), .B1(G868), .B2(new_n569), .ZN(G280));
  INV_X1    g190(.A(new_n609), .ZN(new_n616));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G860), .ZN(G148));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n556), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n609), .A2(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n619), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n474), .A2(new_n470), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  INV_X1    g201(.A(G2100), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n467), .A2(G135), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n481), .A2(G123), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n473), .A2(G111), .ZN(new_n632));
  OAI21_X1  g207(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n630), .B(new_n631), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(G2096), .Z(new_n635));
  NAND3_X1  g210(.A1(new_n628), .A2(new_n629), .A3(new_n635), .ZN(G156));
  INV_X1    g211(.A(KEYINPUT14), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n640), .B2(new_n639), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n642), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  AND3_X1   g225(.A1(new_n649), .A2(G14), .A3(new_n650), .ZN(G401));
  INV_X1    g226(.A(KEYINPUT18), .ZN(new_n652));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(KEYINPUT17), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n653), .A2(new_n654), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n652), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2096), .B(G2100), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2072), .B(G2078), .Z(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n655), .B2(KEYINPUT18), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT80), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n660), .B(new_n663), .ZN(G227));
  XOR2_X1   g239(.A(KEYINPUT81), .B(KEYINPUT19), .Z(new_n665));
  XNOR2_X1  g240(.A(G1971), .B(G1976), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1956), .B(G2474), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT20), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n668), .A2(new_n669), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n667), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n674), .A2(new_n670), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n672), .B(new_n675), .C1(new_n667), .C2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT83), .ZN(new_n678));
  XOR2_X1   g253(.A(G1991), .B(G1996), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT82), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n678), .B(new_n684), .ZN(G229));
  INV_X1    g260(.A(G29), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G26), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT28), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n467), .A2(G140), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n481), .A2(G128), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n473), .A2(G116), .ZN(new_n691));
  OAI21_X1  g266(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n689), .B(new_n690), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G29), .ZN(new_n694));
  AND2_X1   g269(.A1(new_n694), .A2(KEYINPUT87), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(KEYINPUT87), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n688), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G2067), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT95), .B(KEYINPUT23), .Z(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G20), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n700), .B(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(new_n569), .B2(new_n701), .ZN(new_n704));
  INV_X1    g279(.A(G1956), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G1341), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n557), .A2(new_n701), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n701), .B2(G19), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n699), .B(new_n706), .C1(new_n707), .C2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n686), .A2(G35), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT93), .Z(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n487), .B2(G29), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G2090), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n713), .B(new_n715), .Z(new_n716));
  NAND2_X1  g291(.A1(new_n709), .A2(new_n707), .ZN(new_n717));
  NOR2_X1   g292(.A1(G4), .A2(G16), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n616), .B2(G16), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n716), .B(new_n717), .C1(G1348), .C2(new_n719), .ZN(new_n720));
  AOI211_X1 g295(.A(new_n710), .B(new_n720), .C1(G1348), .C2(new_n719), .ZN(new_n721));
  NOR2_X1   g296(.A1(G168), .A2(new_n701), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n701), .B2(G21), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT90), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G1966), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n701), .A2(G5), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G171), .B2(new_n701), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(G1961), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n724), .ZN(new_n730));
  INV_X1    g305(.A(G1966), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n730), .A2(new_n731), .B1(new_n727), .B2(G1961), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n686), .A2(G33), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT25), .ZN(new_n734));
  NAND2_X1  g309(.A1(G103), .A2(G2104), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(G2105), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n473), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n467), .A2(G139), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n738), .B1(new_n473), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT88), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n733), .B1(new_n742), .B2(new_n686), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2072), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n686), .A2(G27), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G164), .B2(new_n686), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G2078), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n467), .A2(G141), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n481), .A2(G129), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n470), .A2(G105), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT26), .Z(new_n752));
  NAND4_X1  g327(.A1(new_n748), .A2(new_n749), .A3(new_n750), .A4(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n754), .A2(new_n686), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n686), .B2(G32), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT27), .B(G1996), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT31), .B(G11), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT30), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n686), .B1(new_n760), .B2(G28), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n761), .A2(KEYINPUT91), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(G28), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n761), .B2(KEYINPUT91), .ZN(new_n764));
  OAI221_X1 g339(.A(new_n759), .B1(new_n762), .B2(new_n764), .C1(new_n634), .C2(new_n686), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n756), .B2(new_n757), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT89), .B(KEYINPUT24), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G34), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n768), .A2(G29), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G160), .B2(G29), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n770), .A2(G2084), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n770), .A2(G2084), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n758), .A2(new_n766), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  NOR3_X1   g348(.A1(new_n744), .A2(new_n747), .A3(new_n773), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n729), .A2(new_n732), .A3(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT92), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n721), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n776), .B2(new_n775), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n701), .A2(G22), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G166), .B2(new_n701), .ZN(new_n780));
  INV_X1    g355(.A(G1971), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  MUX2_X1   g357(.A(G6), .B(G305), .S(G16), .Z(new_n783));
  XOR2_X1   g358(.A(KEYINPUT32), .B(G1981), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n580), .B1(new_n546), .B2(new_n581), .ZN(new_n786));
  MUX2_X1   g361(.A(G23), .B(new_n786), .S(G16), .Z(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT33), .B(G1976), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n782), .A2(new_n785), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(KEYINPUT34), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n467), .A2(G131), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT84), .ZN(new_n793));
  OAI21_X1  g368(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n794));
  INV_X1    g369(.A(G107), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(G2105), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n481), .B2(G119), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  MUX2_X1   g373(.A(G25), .B(new_n798), .S(G29), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT85), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT35), .B(G1991), .Z(new_n801));
  OR2_X1    g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT86), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n701), .B1(G290), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n597), .A2(KEYINPUT86), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n805), .A2(new_n806), .B1(new_n701), .B2(G24), .ZN(new_n807));
  INV_X1    g382(.A(G1986), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n802), .A2(new_n803), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT34), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n782), .A2(new_n811), .A3(new_n785), .A4(new_n789), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n791), .A2(new_n809), .A3(new_n810), .A4(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT36), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n778), .A2(new_n814), .ZN(G150));
  NOR2_X1   g390(.A1(G150), .A2(KEYINPUT96), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT96), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n778), .B2(new_n814), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n816), .A2(new_n818), .ZN(G311));
  XNOR2_X1  g394(.A(KEYINPUT97), .B(G93), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n546), .A2(new_n820), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  INV_X1    g397(.A(G55), .ZN(new_n823));
  OAI22_X1  g398(.A1(new_n822), .A2(new_n528), .B1(new_n823), .B2(new_n535), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(G860), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT37), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n616), .A2(G559), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT38), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n557), .A2(new_n825), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n826), .A2(new_n556), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n830), .B(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT98), .ZN(new_n837));
  AOI21_X1  g412(.A(G860), .B1(new_n834), .B2(new_n835), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n828), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT99), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(G145));
  XNOR2_X1  g416(.A(new_n798), .B(new_n625), .ZN(new_n842));
  AOI22_X1  g417(.A1(G130), .A2(new_n481), .B1(new_n467), .B2(G142), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT100), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n844), .A2(new_n473), .A3(G118), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n844), .B1(new_n473), .B2(G118), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n846), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n843), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n842), .B(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n510), .B(new_n693), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n754), .ZN(new_n852));
  MUX2_X1   g427(.A(new_n740), .B(new_n742), .S(new_n852), .Z(new_n853));
  INV_X1    g428(.A(KEYINPUT102), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n850), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n854), .B2(new_n853), .ZN(new_n856));
  XNOR2_X1  g431(.A(G160), .B(new_n634), .ZN(new_n857));
  XNOR2_X1  g432(.A(G162), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT103), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n849), .B(KEYINPUT101), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n856), .B(new_n859), .C1(new_n853), .C2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(G37), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n860), .B(new_n853), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(new_n858), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n861), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g441(.A1(new_n826), .A2(new_n619), .ZN(new_n867));
  XNOR2_X1  g442(.A(G305), .B(KEYINPUT105), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(G303), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n597), .B(new_n786), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT42), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n833), .B(new_n621), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n616), .A2(new_n569), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT41), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n569), .B1(new_n603), .B2(new_n608), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n609), .A2(G299), .ZN(new_n881));
  OAI21_X1  g456(.A(KEYINPUT41), .B1(new_n881), .B2(new_n878), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n880), .A2(new_n882), .A3(KEYINPUT104), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n881), .A2(new_n878), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n885), .A3(new_n877), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n875), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n884), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n887), .B1(new_n888), .B2(new_n875), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n874), .B(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n867), .B1(new_n890), .B2(new_n619), .ZN(G295));
  OAI21_X1  g466(.A(new_n867), .B1(new_n890), .B2(new_n619), .ZN(G331));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n557), .A2(new_n825), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n826), .A2(new_n556), .ZN(new_n895));
  OAI21_X1  g470(.A(G301), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(G171), .A2(new_n831), .A3(new_n832), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n896), .A2(G168), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(G168), .B1(new_n896), .B2(new_n897), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n883), .B(new_n886), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n899), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n896), .A2(G168), .A3(new_n897), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n884), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n873), .B1(new_n904), .B2(KEYINPUT106), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n900), .A2(new_n903), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(G37), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n900), .A2(new_n903), .A3(new_n873), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n893), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n873), .ZN(new_n913));
  AOI22_X1  g488(.A1(new_n901), .A2(new_n902), .B1(new_n880), .B2(new_n882), .ZN(new_n914));
  NOR3_X1   g489(.A1(new_n898), .A2(new_n899), .A3(new_n888), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n916), .A2(new_n909), .A3(new_n862), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT107), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n916), .A2(new_n909), .A3(KEYINPUT107), .A4(new_n862), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(KEYINPUT43), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n912), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n922), .B1(new_n912), .B2(new_n921), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n910), .B1(new_n908), .B2(new_n909), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n911), .A2(new_n862), .A3(new_n916), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI22_X1  g502(.A1(new_n923), .A2(new_n924), .B1(KEYINPUT44), .B2(new_n927), .ZN(G397));
  XNOR2_X1  g503(.A(KEYINPUT68), .B(KEYINPUT4), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT69), .B1(new_n502), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n930), .A2(new_n503), .A3(new_n501), .ZN(new_n931));
  AOI21_X1  g506(.A(G1384), .B1(new_n931), .B2(new_n492), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n932), .A2(KEYINPUT45), .ZN(new_n933));
  INV_X1    g508(.A(G40), .ZN(new_n934));
  NOR3_X1   g509(.A1(new_n472), .A2(new_n477), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n936), .A2(G1996), .A3(new_n753), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT109), .ZN(new_n938));
  INV_X1    g513(.A(new_n936), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n693), .B(new_n698), .ZN(new_n940));
  INV_X1    g515(.A(G1996), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n940), .B1(new_n941), .B2(new_n754), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n938), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n798), .B(new_n801), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n943), .B1(new_n936), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n597), .B(new_n808), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n945), .B1(new_n939), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G1384), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n510), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT45), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n935), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n731), .B1(new_n951), .B2(new_n933), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n949), .A2(KEYINPUT113), .A3(KEYINPUT50), .ZN(new_n953));
  AOI22_X1  g528(.A1(new_n467), .A2(G137), .B1(G101), .B2(new_n470), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n475), .A2(new_n476), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n954), .B(G40), .C1(new_n473), .C2(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n956), .B1(new_n932), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT113), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT50), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n959), .B1(new_n932), .B2(new_n960), .ZN(new_n961));
  XOR2_X1   g536(.A(KEYINPUT121), .B(G2084), .Z(new_n962));
  NAND4_X1  g537(.A1(new_n953), .A2(new_n958), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n952), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(G8), .B1(new_n964), .B2(G286), .ZN(new_n965));
  AOI21_X1  g540(.A(G168), .B1(new_n952), .B2(new_n963), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT51), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n968), .B(G8), .C1(new_n964), .C2(G286), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n970), .A2(KEYINPUT62), .ZN(new_n971));
  INV_X1    g546(.A(G2078), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n956), .B1(new_n932), .B2(KEYINPUT45), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT110), .B1(new_n949), .B2(new_n950), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n932), .A2(new_n975), .A3(KEYINPUT45), .ZN(new_n976));
  OAI211_X1 g551(.A(KEYINPUT111), .B(new_n973), .C1(new_n974), .C2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n949), .A2(KEYINPUT110), .A3(new_n950), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n975), .B1(new_n932), .B2(KEYINPUT45), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT111), .B1(new_n981), .B2(new_n973), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n972), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n951), .A2(new_n933), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n984), .A2(G2078), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n953), .A2(new_n958), .A3(new_n961), .ZN(new_n988));
  INV_X1    g563(.A(G1961), .ZN(new_n989));
  AOI22_X1  g564(.A1(new_n986), .A2(new_n987), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(G301), .B1(new_n985), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT62), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n993), .B1(new_n967), .B2(new_n969), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n971), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n973), .B1(new_n974), .B2(new_n976), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(G2078), .B1(new_n998), .B2(new_n977), .ZN(new_n999));
  OAI211_X1 g574(.A(G301), .B(new_n990), .C1(new_n999), .C2(KEYINPUT53), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT54), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n970), .B1(new_n1001), .B2(new_n991), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n569), .B(KEYINPUT57), .ZN(new_n1003));
  XNOR2_X1  g578(.A(KEYINPUT56), .B(G2072), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n981), .A2(new_n973), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n932), .A2(new_n960), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1006), .B(new_n935), .C1(new_n932), .C2(new_n957), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n705), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1003), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G1348), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n949), .A2(new_n956), .ZN(new_n1011));
  AOI22_X1  g586(.A1(new_n988), .A2(new_n1010), .B1(new_n698), .B2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1012), .A2(new_n609), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1003), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1009), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1009), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT61), .ZN(new_n1017));
  OR3_X1    g592(.A1(new_n1016), .A2(new_n1014), .A3(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(KEYINPUT58), .B(G1341), .ZN(new_n1019));
  OAI22_X1  g594(.A1(new_n996), .A2(G1996), .B1(new_n1011), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1020), .A2(KEYINPUT122), .A3(new_n557), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT59), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT59), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1020), .A2(KEYINPUT122), .A3(new_n1023), .A4(new_n557), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n1012), .A2(KEYINPUT60), .A3(new_n609), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n609), .B1(new_n1012), .B2(KEYINPUT60), .ZN(new_n1027));
  OAI22_X1  g602(.A1(new_n1026), .A2(new_n1027), .B1(KEYINPUT60), .B2(new_n1012), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1017), .B1(new_n1016), .B2(new_n1014), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1018), .A2(new_n1025), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1002), .B1(new_n1015), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT123), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n992), .A2(new_n1032), .A3(new_n1000), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n985), .A2(KEYINPUT123), .A3(G301), .A4(new_n990), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n995), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n580), .B(G1976), .C1(new_n581), .C2(new_n546), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1039), .B(G8), .C1(new_n949), .C2(new_n956), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G8), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1043), .B1(new_n935), .B2(new_n932), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1044), .A2(KEYINPUT116), .A3(new_n1039), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1042), .A2(new_n1045), .A3(KEYINPUT52), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1042), .A2(new_n1045), .A3(KEYINPUT117), .A4(KEYINPUT52), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT49), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n521), .A2(G86), .A3(new_n522), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n517), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1053));
  INV_X1    g628(.A(G48), .ZN(new_n1054));
  OAI22_X1  g629(.A1(new_n1053), .A2(new_n528), .B1(new_n1054), .B2(new_n535), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n1052), .A2(G1981), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G1981), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1057), .B1(new_n587), .B2(new_n588), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1051), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(G1981), .B1(new_n1052), .B2(new_n1055), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n587), .A2(new_n1057), .A3(new_n588), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(KEYINPUT49), .A3(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(new_n1044), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G1976), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n578), .A2(new_n1064), .A3(new_n582), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1065), .A2(new_n1066), .A3(new_n1044), .A4(new_n1039), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1063), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1038), .B1(new_n1050), .B2(new_n1069), .ZN(new_n1070));
  AOI211_X1 g645(.A(KEYINPUT120), .B(new_n1068), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1071));
  NAND2_X1  g646(.A1(G303), .A2(G8), .ZN(new_n1072));
  XOR2_X1   g647(.A(new_n1072), .B(KEYINPUT55), .Z(new_n1073));
  NAND3_X1  g648(.A1(new_n998), .A2(new_n781), .A3(new_n977), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n1075));
  AOI21_X1  g650(.A(G2090), .B1(new_n1007), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1076), .B1(new_n1075), .B2(new_n1007), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1043), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1078));
  OAI22_X1  g653(.A1(new_n1070), .A2(new_n1071), .B1(new_n1073), .B2(new_n1078), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n978), .A2(new_n982), .A3(G1971), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n988), .A2(G2090), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT114), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT114), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1081), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1074), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1082), .A2(G8), .A3(new_n1073), .A4(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(KEYINPUT115), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1085), .A2(G8), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT115), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1088), .A2(new_n1089), .A3(new_n1073), .A4(new_n1082), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1079), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  AOI211_X1 g667(.A(new_n1043), .B(G286), .C1(new_n952), .C2(new_n963), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT63), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  AND4_X1   g669(.A1(KEYINPUT63), .A2(new_n1050), .A3(new_n1069), .A4(new_n1093), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1082), .A2(G8), .A3(new_n1085), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1095), .B1(new_n1096), .B2(new_n1073), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1097), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1098));
  OAI22_X1  g673(.A1(new_n1037), .A2(new_n1092), .B1(new_n1094), .B2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1087), .A2(new_n1090), .A3(new_n1050), .A4(new_n1069), .ZN(new_n1100));
  AOI211_X1 g675(.A(G1976), .B(G288), .C1(new_n1059), .C2(new_n1062), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1044), .B1(new_n1101), .B2(new_n1056), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1100), .A2(KEYINPUT118), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT118), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n947), .B1(new_n1099), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT46), .B1(new_n939), .B2(new_n941), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1107), .B(KEYINPUT124), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n753), .B1(KEYINPUT46), .B2(new_n941), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n940), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1108), .B1(new_n936), .B2(new_n1110), .ZN(new_n1111));
  XOR2_X1   g686(.A(new_n1111), .B(KEYINPUT47), .Z(new_n1112));
  NAND4_X1  g687(.A1(new_n943), .A2(new_n801), .A3(new_n793), .A4(new_n797), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n693), .A2(G2067), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n936), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NOR3_X1   g690(.A1(G290), .A2(new_n936), .A3(G1986), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1116), .B(KEYINPUT125), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1117), .B(KEYINPUT48), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1118), .A2(new_n945), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1112), .A2(new_n1115), .A3(new_n1119), .ZN(new_n1120));
  XOR2_X1   g695(.A(new_n1120), .B(KEYINPUT126), .Z(new_n1121));
  NAND2_X1  g696(.A1(new_n1106), .A2(new_n1121), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g697(.A1(G229), .A2(new_n462), .A3(G401), .A4(G227), .ZN(new_n1124));
  NAND2_X1  g698(.A1(new_n865), .A2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g699(.A1(new_n927), .A2(new_n1125), .ZN(G308));
  INV_X1    g700(.A(G308), .ZN(G225));
endmodule


