

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X2 U323 ( .A(n361), .B(n360), .ZN(n576) );
  XNOR2_X1 U324 ( .A(n448), .B(KEYINPUT121), .ZN(n564) );
  XNOR2_X1 U325 ( .A(n446), .B(n445), .ZN(n528) );
  XNOR2_X1 U326 ( .A(n309), .B(n308), .ZN(n554) );
  XNOR2_X1 U327 ( .A(n414), .B(n291), .ZN(n308) );
  XNOR2_X1 U328 ( .A(n477), .B(n476), .ZN(n500) );
  AND2_X1 U329 ( .A1(G232GAT), .A2(G233GAT), .ZN(n291) );
  NOR2_X1 U330 ( .A1(n525), .A2(n519), .ZN(n387) );
  XNOR2_X1 U331 ( .A(KEYINPUT10), .B(KEYINPUT79), .ZN(n294) );
  XNOR2_X1 U332 ( .A(n375), .B(n294), .ZN(n299) );
  NAND2_X1 U333 ( .A1(n528), .A2(n465), .ZN(n453) );
  INV_X1 U334 ( .A(KEYINPUT37), .ZN(n473) );
  XNOR2_X1 U335 ( .A(n473), .B(KEYINPUT106), .ZN(n474) );
  NOR2_X1 U336 ( .A1(n447), .A2(n528), .ZN(n448) );
  XNOR2_X1 U337 ( .A(n475), .B(n474), .ZN(n515) );
  INV_X1 U338 ( .A(G43GAT), .ZN(n478) );
  XNOR2_X1 U339 ( .A(G183GAT), .B(KEYINPUT122), .ZN(n450) );
  XNOR2_X1 U340 ( .A(n478), .B(KEYINPUT40), .ZN(n479) );
  XNOR2_X1 U341 ( .A(n451), .B(n450), .ZN(G1350GAT) );
  XNOR2_X1 U342 ( .A(n480), .B(n479), .ZN(G1330GAT) );
  XOR2_X1 U343 ( .A(KEYINPUT80), .B(G218GAT), .Z(n293) );
  XNOR2_X1 U344 ( .A(G36GAT), .B(G190GAT), .ZN(n292) );
  XNOR2_X1 U345 ( .A(n293), .B(n292), .ZN(n375) );
  INV_X1 U346 ( .A(n299), .ZN(n297) );
  XOR2_X1 U347 ( .A(G29GAT), .B(G134GAT), .Z(n389) );
  XNOR2_X1 U348 ( .A(n389), .B(KEYINPUT9), .ZN(n295) );
  XOR2_X1 U349 ( .A(n295), .B(KEYINPUT11), .Z(n298) );
  INV_X1 U350 ( .A(n298), .ZN(n296) );
  NAND2_X1 U351 ( .A1(n297), .A2(n296), .ZN(n301) );
  NAND2_X1 U352 ( .A1(n299), .A2(n298), .ZN(n300) );
  NAND2_X1 U353 ( .A1(n301), .A2(n300), .ZN(n307) );
  XOR2_X1 U354 ( .A(G43GAT), .B(KEYINPUT8), .Z(n303) );
  XNOR2_X1 U355 ( .A(KEYINPUT70), .B(KEYINPUT7), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n303), .B(n302), .ZN(n331) );
  XOR2_X1 U357 ( .A(G92GAT), .B(G106GAT), .Z(n305) );
  XNOR2_X1 U358 ( .A(G99GAT), .B(G85GAT), .ZN(n304) );
  XNOR2_X1 U359 ( .A(n305), .B(n304), .ZN(n350) );
  XNOR2_X1 U360 ( .A(n331), .B(n350), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n309) );
  XOR2_X1 U362 ( .A(G50GAT), .B(G162GAT), .Z(n414) );
  XNOR2_X1 U363 ( .A(KEYINPUT81), .B(n554), .ZN(n565) );
  XNOR2_X1 U364 ( .A(KEYINPUT36), .B(n565), .ZN(n583) );
  XOR2_X1 U365 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n311) );
  NAND2_X1 U366 ( .A1(G231GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U367 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U368 ( .A(n312), .B(KEYINPUT83), .Z(n317) );
  XNOR2_X1 U369 ( .A(G71GAT), .B(G57GAT), .ZN(n313) );
  XNOR2_X1 U370 ( .A(n313), .B(KEYINPUT13), .ZN(n359) );
  XOR2_X1 U371 ( .A(G211GAT), .B(KEYINPUT82), .Z(n315) );
  XNOR2_X1 U372 ( .A(G8GAT), .B(G183GAT), .ZN(n314) );
  XNOR2_X1 U373 ( .A(n315), .B(n314), .ZN(n382) );
  XNOR2_X1 U374 ( .A(n359), .B(n382), .ZN(n316) );
  XNOR2_X1 U375 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U376 ( .A(KEYINPUT14), .B(G64GAT), .Z(n319) );
  XNOR2_X1 U377 ( .A(G155GAT), .B(G78GAT), .ZN(n318) );
  XNOR2_X1 U378 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U379 ( .A(n321), .B(n320), .Z(n323) );
  XOR2_X1 U380 ( .A(G22GAT), .B(G15GAT), .Z(n328) );
  XOR2_X1 U381 ( .A(G1GAT), .B(G127GAT), .Z(n388) );
  XNOR2_X1 U382 ( .A(n328), .B(n388), .ZN(n322) );
  XNOR2_X1 U383 ( .A(n323), .B(n322), .ZN(n580) );
  NOR2_X1 U384 ( .A1(n583), .A2(n580), .ZN(n324) );
  XNOR2_X1 U385 ( .A(KEYINPUT45), .B(n324), .ZN(n363) );
  XOR2_X1 U386 ( .A(G141GAT), .B(G113GAT), .Z(n326) );
  XNOR2_X1 U387 ( .A(G29GAT), .B(G1GAT), .ZN(n325) );
  XNOR2_X1 U388 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U389 ( .A(n327), .B(G36GAT), .Z(n330) );
  XNOR2_X1 U390 ( .A(n328), .B(G50GAT), .ZN(n329) );
  XNOR2_X1 U391 ( .A(n330), .B(n329), .ZN(n335) );
  XOR2_X1 U392 ( .A(n331), .B(KEYINPUT68), .Z(n333) );
  NAND2_X1 U393 ( .A1(G229GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U394 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U395 ( .A(n335), .B(n334), .Z(n343) );
  XOR2_X1 U396 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n337) );
  XNOR2_X1 U397 ( .A(KEYINPUT66), .B(KEYINPUT30), .ZN(n336) );
  XNOR2_X1 U398 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U399 ( .A(KEYINPUT69), .B(G8GAT), .Z(n339) );
  XNOR2_X1 U400 ( .A(G169GAT), .B(G197GAT), .ZN(n338) );
  XNOR2_X1 U401 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U402 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n343), .B(n342), .ZN(n573) );
  INV_X1 U404 ( .A(n573), .ZN(n544) );
  XOR2_X1 U405 ( .A(G176GAT), .B(G64GAT), .Z(n373) );
  XOR2_X1 U406 ( .A(KEYINPUT75), .B(KEYINPUT73), .Z(n345) );
  XNOR2_X1 U407 ( .A(G120GAT), .B(KEYINPUT72), .ZN(n344) );
  XNOR2_X1 U408 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U409 ( .A(n373), .B(n346), .Z(n348) );
  NAND2_X1 U410 ( .A1(G230GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U411 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U412 ( .A(n349), .B(KEYINPUT32), .ZN(n352) );
  XOR2_X1 U413 ( .A(n350), .B(KEYINPUT31), .Z(n351) );
  XNOR2_X1 U414 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U415 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n354) );
  XNOR2_X1 U416 ( .A(KEYINPUT71), .B(KEYINPUT33), .ZN(n353) );
  XNOR2_X1 U417 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U418 ( .A(n356), .B(n355), .ZN(n361) );
  XOR2_X1 U419 ( .A(G78GAT), .B(G204GAT), .Z(n358) );
  XNOR2_X1 U420 ( .A(G148GAT), .B(KEYINPUT74), .ZN(n357) );
  XNOR2_X1 U421 ( .A(n358), .B(n357), .ZN(n415) );
  XOR2_X1 U422 ( .A(n359), .B(n415), .Z(n360) );
  NOR2_X1 U423 ( .A1(n544), .A2(n576), .ZN(n362) );
  NAND2_X1 U424 ( .A1(n363), .A2(n362), .ZN(n370) );
  XNOR2_X1 U425 ( .A(n576), .B(KEYINPUT41), .ZN(n549) );
  NOR2_X1 U426 ( .A1(n573), .A2(n549), .ZN(n365) );
  XNOR2_X1 U427 ( .A(KEYINPUT115), .B(KEYINPUT46), .ZN(n364) );
  XNOR2_X1 U428 ( .A(n365), .B(n364), .ZN(n367) );
  XOR2_X1 U429 ( .A(n580), .B(KEYINPUT114), .Z(n535) );
  NOR2_X1 U430 ( .A1(n554), .A2(n535), .ZN(n366) );
  NAND2_X1 U431 ( .A1(n367), .A2(n366), .ZN(n368) );
  XOR2_X1 U432 ( .A(n368), .B(KEYINPUT47), .Z(n369) );
  NAND2_X1 U433 ( .A1(n370), .A2(n369), .ZN(n372) );
  INV_X1 U434 ( .A(KEYINPUT48), .ZN(n371) );
  XNOR2_X1 U435 ( .A(n372), .B(n371), .ZN(n525) );
  NAND2_X1 U436 ( .A1(G226GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U437 ( .A(n374), .B(n373), .ZN(n386) );
  XNOR2_X1 U438 ( .A(n375), .B(KEYINPUT95), .ZN(n376) );
  XNOR2_X1 U439 ( .A(n376), .B(KEYINPUT96), .ZN(n379) );
  XNOR2_X1 U440 ( .A(G204GAT), .B(G92GAT), .ZN(n377) );
  XOR2_X1 U441 ( .A(G197GAT), .B(KEYINPUT21), .Z(n412) );
  XNOR2_X1 U442 ( .A(n377), .B(n412), .ZN(n378) );
  XOR2_X1 U443 ( .A(n379), .B(n378), .Z(n384) );
  XOR2_X1 U444 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n381) );
  XNOR2_X1 U445 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n380) );
  XNOR2_X1 U446 ( .A(n381), .B(n380), .ZN(n443) );
  XNOR2_X1 U447 ( .A(n443), .B(n382), .ZN(n383) );
  XNOR2_X1 U448 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U449 ( .A(n386), .B(n385), .ZN(n519) );
  XNOR2_X1 U450 ( .A(n387), .B(KEYINPUT54), .ZN(n408) );
  XOR2_X1 U451 ( .A(G85GAT), .B(G162GAT), .Z(n391) );
  XNOR2_X1 U452 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U453 ( .A(n391), .B(n390), .ZN(n405) );
  XOR2_X1 U454 ( .A(G148GAT), .B(KEYINPUT93), .Z(n393) );
  XNOR2_X1 U455 ( .A(KEYINPUT92), .B(KEYINPUT4), .ZN(n392) );
  XNOR2_X1 U456 ( .A(n393), .B(n392), .ZN(n397) );
  XOR2_X1 U457 ( .A(G57GAT), .B(KEYINPUT6), .Z(n395) );
  XNOR2_X1 U458 ( .A(KEYINPUT5), .B(KEYINPUT1), .ZN(n394) );
  XNOR2_X1 U459 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U460 ( .A(n397), .B(n396), .Z(n403) );
  XOR2_X1 U461 ( .A(G120GAT), .B(KEYINPUT85), .Z(n399) );
  XNOR2_X1 U462 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n398) );
  XNOR2_X1 U463 ( .A(n399), .B(n398), .ZN(n444) );
  XOR2_X1 U464 ( .A(G155GAT), .B(KEYINPUT2), .Z(n401) );
  XNOR2_X1 U465 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n400) );
  XNOR2_X1 U466 ( .A(n401), .B(n400), .ZN(n420) );
  XNOR2_X1 U467 ( .A(n444), .B(n420), .ZN(n402) );
  XNOR2_X1 U468 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U469 ( .A(n405), .B(n404), .Z(n407) );
  NAND2_X1 U470 ( .A1(G225GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U471 ( .A(n407), .B(n406), .ZN(n462) );
  XNOR2_X1 U472 ( .A(KEYINPUT94), .B(n462), .ZN(n517) );
  NAND2_X1 U473 ( .A1(n408), .A2(n517), .ZN(n409) );
  XNOR2_X1 U474 ( .A(n409), .B(KEYINPUT64), .ZN(n571) );
  XOR2_X1 U475 ( .A(KEYINPUT22), .B(KEYINPUT90), .Z(n411) );
  XNOR2_X1 U476 ( .A(KEYINPUT91), .B(KEYINPUT23), .ZN(n410) );
  XNOR2_X1 U477 ( .A(n411), .B(n410), .ZN(n413) );
  XOR2_X1 U478 ( .A(n413), .B(n412), .Z(n417) );
  XNOR2_X1 U479 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U480 ( .A(n417), .B(n416), .ZN(n426) );
  XOR2_X1 U481 ( .A(G211GAT), .B(G218GAT), .Z(n419) );
  XNOR2_X1 U482 ( .A(G22GAT), .B(G106GAT), .ZN(n418) );
  XNOR2_X1 U483 ( .A(n419), .B(n418), .ZN(n424) );
  XOR2_X1 U484 ( .A(n420), .B(KEYINPUT24), .Z(n422) );
  NAND2_X1 U485 ( .A1(G228GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U486 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U487 ( .A(n424), .B(n423), .Z(n425) );
  XNOR2_X1 U488 ( .A(n426), .B(n425), .ZN(n465) );
  NOR2_X1 U489 ( .A1(n571), .A2(n465), .ZN(n427) );
  XNOR2_X1 U490 ( .A(n427), .B(KEYINPUT55), .ZN(n447) );
  XOR2_X1 U491 ( .A(G134GAT), .B(G99GAT), .Z(n429) );
  XNOR2_X1 U492 ( .A(G43GAT), .B(G190GAT), .ZN(n428) );
  XNOR2_X1 U493 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U494 ( .A(G176GAT), .B(G71GAT), .Z(n431) );
  XNOR2_X1 U495 ( .A(G15GAT), .B(G127GAT), .ZN(n430) );
  XNOR2_X1 U496 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U497 ( .A(n433), .B(n432), .Z(n438) );
  XOR2_X1 U498 ( .A(KEYINPUT20), .B(KEYINPUT87), .Z(n435) );
  NAND2_X1 U499 ( .A1(G227GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U500 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U501 ( .A(KEYINPUT86), .B(n436), .ZN(n437) );
  XNOR2_X1 U502 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U503 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n440) );
  XNOR2_X1 U504 ( .A(G183GAT), .B(KEYINPUT65), .ZN(n439) );
  XNOR2_X1 U505 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U506 ( .A(n442), .B(n441), .Z(n446) );
  XNOR2_X1 U507 ( .A(n444), .B(n443), .ZN(n445) );
  INV_X1 U508 ( .A(n564), .ZN(n449) );
  NAND2_X1 U509 ( .A1(n449), .A2(n535), .ZN(n451) );
  XOR2_X1 U510 ( .A(KEYINPUT38), .B(KEYINPUT107), .Z(n477) );
  NOR2_X1 U511 ( .A1(n576), .A2(n573), .ZN(n452) );
  XNOR2_X1 U512 ( .A(n452), .B(KEYINPUT78), .ZN(n486) );
  XNOR2_X1 U513 ( .A(KEYINPUT27), .B(n519), .ZN(n466) );
  XOR2_X1 U514 ( .A(KEYINPUT99), .B(KEYINPUT26), .Z(n454) );
  XNOR2_X1 U515 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U516 ( .A(KEYINPUT98), .B(n455), .ZN(n570) );
  OR2_X1 U517 ( .A1(n466), .A2(n570), .ZN(n461) );
  XOR2_X1 U518 ( .A(KEYINPUT25), .B(KEYINPUT101), .Z(n459) );
  NOR2_X1 U519 ( .A1(n528), .A2(n519), .ZN(n456) );
  NOR2_X1 U520 ( .A1(n465), .A2(n456), .ZN(n457) );
  XNOR2_X1 U521 ( .A(n457), .B(KEYINPUT100), .ZN(n458) );
  XNOR2_X1 U522 ( .A(n459), .B(n458), .ZN(n460) );
  NAND2_X1 U523 ( .A1(n461), .A2(n460), .ZN(n463) );
  NAND2_X1 U524 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U525 ( .A(n464), .B(KEYINPUT102), .ZN(n470) );
  XNOR2_X1 U526 ( .A(KEYINPUT28), .B(n465), .ZN(n493) );
  NOR2_X1 U527 ( .A1(n517), .A2(n466), .ZN(n467) );
  XNOR2_X1 U528 ( .A(n467), .B(KEYINPUT97), .ZN(n526) );
  NOR2_X1 U529 ( .A1(n493), .A2(n526), .ZN(n468) );
  NAND2_X1 U530 ( .A1(n468), .A2(n528), .ZN(n469) );
  NAND2_X1 U531 ( .A1(n470), .A2(n469), .ZN(n484) );
  NAND2_X1 U532 ( .A1(n580), .A2(n484), .ZN(n471) );
  XOR2_X1 U533 ( .A(KEYINPUT105), .B(n471), .Z(n472) );
  NOR2_X1 U534 ( .A1(n472), .A2(n583), .ZN(n475) );
  NAND2_X1 U535 ( .A1(n486), .A2(n515), .ZN(n476) );
  NOR2_X1 U536 ( .A1(n528), .A2(n500), .ZN(n480) );
  XOR2_X1 U537 ( .A(KEYINPUT16), .B(KEYINPUT84), .Z(n483) );
  INV_X1 U538 ( .A(n580), .ZN(n481) );
  NAND2_X1 U539 ( .A1(n481), .A2(n565), .ZN(n482) );
  XNOR2_X1 U540 ( .A(n483), .B(n482), .ZN(n485) );
  AND2_X1 U541 ( .A1(n485), .A2(n484), .ZN(n503) );
  NAND2_X1 U542 ( .A1(n503), .A2(n486), .ZN(n494) );
  NOR2_X1 U543 ( .A1(n517), .A2(n494), .ZN(n487) );
  XOR2_X1 U544 ( .A(KEYINPUT34), .B(n487), .Z(n488) );
  XNOR2_X1 U545 ( .A(G1GAT), .B(n488), .ZN(G1324GAT) );
  NOR2_X1 U546 ( .A1(n519), .A2(n494), .ZN(n490) );
  XNOR2_X1 U547 ( .A(G8GAT), .B(KEYINPUT103), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n490), .B(n489), .ZN(G1325GAT) );
  NOR2_X1 U549 ( .A1(n528), .A2(n494), .ZN(n492) );
  XNOR2_X1 U550 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n492), .B(n491), .ZN(G1326GAT) );
  INV_X1 U552 ( .A(n493), .ZN(n529) );
  NOR2_X1 U553 ( .A1(n529), .A2(n494), .ZN(n495) );
  XOR2_X1 U554 ( .A(KEYINPUT104), .B(n495), .Z(n496) );
  XNOR2_X1 U555 ( .A(G22GAT), .B(n496), .ZN(G1327GAT) );
  NOR2_X1 U556 ( .A1(n500), .A2(n517), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n497), .B(KEYINPUT39), .ZN(n498) );
  XNOR2_X1 U558 ( .A(G29GAT), .B(n498), .ZN(G1328GAT) );
  NOR2_X1 U559 ( .A1(n500), .A2(n519), .ZN(n499) );
  XOR2_X1 U560 ( .A(G36GAT), .B(n499), .Z(G1329GAT) );
  NOR2_X1 U561 ( .A1(n500), .A2(n529), .ZN(n501) );
  XOR2_X1 U562 ( .A(G50GAT), .B(n501), .Z(n502) );
  XNOR2_X1 U563 ( .A(KEYINPUT108), .B(n502), .ZN(G1331GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT109), .B(n549), .Z(n558) );
  NOR2_X1 U565 ( .A1(n544), .A2(n558), .ZN(n516) );
  NAND2_X1 U566 ( .A1(n516), .A2(n503), .ZN(n512) );
  NOR2_X1 U567 ( .A1(n517), .A2(n512), .ZN(n505) );
  XNOR2_X1 U568 ( .A(KEYINPUT42), .B(KEYINPUT110), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U570 ( .A(G57GAT), .B(n506), .Z(G1332GAT) );
  NOR2_X1 U571 ( .A1(n519), .A2(n512), .ZN(n508) );
  XNOR2_X1 U572 ( .A(G64GAT), .B(KEYINPUT111), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(G1333GAT) );
  NOR2_X1 U574 ( .A1(n528), .A2(n512), .ZN(n510) );
  XNOR2_X1 U575 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U577 ( .A(G71GAT), .B(n511), .ZN(G1334GAT) );
  NOR2_X1 U578 ( .A1(n529), .A2(n512), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  NAND2_X1 U581 ( .A1(n516), .A2(n515), .ZN(n522) );
  NOR2_X1 U582 ( .A1(n517), .A2(n522), .ZN(n518) );
  XOR2_X1 U583 ( .A(G85GAT), .B(n518), .Z(G1336GAT) );
  NOR2_X1 U584 ( .A1(n519), .A2(n522), .ZN(n520) );
  XOR2_X1 U585 ( .A(G92GAT), .B(n520), .Z(G1337GAT) );
  NOR2_X1 U586 ( .A1(n528), .A2(n522), .ZN(n521) );
  XOR2_X1 U587 ( .A(G99GAT), .B(n521), .Z(G1338GAT) );
  NOR2_X1 U588 ( .A1(n529), .A2(n522), .ZN(n523) );
  XOR2_X1 U589 ( .A(KEYINPUT44), .B(n523), .Z(n524) );
  XNOR2_X1 U590 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  NOR2_X1 U591 ( .A1(n525), .A2(n526), .ZN(n527) );
  XOR2_X1 U592 ( .A(KEYINPUT116), .B(n527), .Z(n543) );
  NOR2_X1 U593 ( .A1(n528), .A2(n543), .ZN(n530) );
  NAND2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n540) );
  NOR2_X1 U595 ( .A1(n573), .A2(n540), .ZN(n532) );
  XNOR2_X1 U596 ( .A(G113GAT), .B(KEYINPUT117), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(G1340GAT) );
  NOR2_X1 U598 ( .A1(n558), .A2(n540), .ZN(n534) );
  XNOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(G1341GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n538) );
  INV_X1 U602 ( .A(n540), .ZN(n536) );
  NAND2_X1 U603 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U605 ( .A(G127GAT), .B(n539), .Z(G1342GAT) );
  NOR2_X1 U606 ( .A1(n565), .A2(n540), .ZN(n542) );
  XNOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(G1343GAT) );
  XOR2_X1 U609 ( .A(G141GAT), .B(KEYINPUT119), .Z(n546) );
  NOR2_X1 U610 ( .A1(n543), .A2(n570), .ZN(n555) );
  NAND2_X1 U611 ( .A1(n555), .A2(n544), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n548) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n551) );
  INV_X1 U616 ( .A(n555), .ZN(n552) );
  NOR2_X1 U617 ( .A1(n549), .A2(n552), .ZN(n550) );
  XOR2_X1 U618 ( .A(n551), .B(n550), .Z(G1345GAT) );
  NOR2_X1 U619 ( .A1(n580), .A2(n552), .ZN(n553) );
  XOR2_X1 U620 ( .A(G155GAT), .B(n553), .Z(G1346GAT) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U623 ( .A1(n573), .A2(n564), .ZN(n557) );
  XOR2_X1 U624 ( .A(G169GAT), .B(n557), .Z(G1348GAT) );
  NOR2_X1 U625 ( .A1(n564), .A2(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(n561), .ZN(G1349GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n563) );
  XNOR2_X1 U630 ( .A(G190GAT), .B(KEYINPUT124), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n563), .B(n562), .ZN(n567) );
  NOR2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U633 ( .A(n567), .B(n566), .Z(G1351GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n569) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(n575) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(KEYINPUT125), .B(n572), .ZN(n582) );
  NOR2_X1 U639 ( .A1(n573), .A2(n582), .ZN(n574) );
  XOR2_X1 U640 ( .A(n575), .B(n574), .Z(G1352GAT) );
  XOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT61), .Z(n579) );
  INV_X1 U642 ( .A(n582), .ZN(n577) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n582), .ZN(n581) );
  XOR2_X1 U646 ( .A(G211GAT), .B(n581), .Z(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(KEYINPUT62), .B(n584), .Z(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

