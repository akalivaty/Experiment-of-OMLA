//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1285, new_n1286, new_n1287, new_n1289, new_n1290, new_n1291,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n207), .B(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n205), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n202), .A2(G50), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  AOI211_X1 g0022(.A(new_n209), .B(new_n217), .C1(new_n220), .C2(new_n222), .ZN(G361));
  XOR2_X1   g0023(.A(G238), .B(G244), .Z(new_n224));
  XNOR2_X1  g0024(.A(G226), .B(G232), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G264), .B(G270), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n228), .B(new_n231), .ZN(G358));
  XNOR2_X1  g0032(.A(G68), .B(G77), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G58), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT66), .B(G50), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G87), .B(G97), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G351));
  INV_X1    g0040(.A(G33), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(KEYINPUT3), .ZN(new_n242));
  INV_X1    g0042(.A(KEYINPUT3), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g0045(.A(KEYINPUT7), .B1(new_n245), .B2(new_n219), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT7), .ZN(new_n247));
  AOI211_X1 g0047(.A(new_n247), .B(G20), .C1(new_n242), .C2(new_n244), .ZN(new_n248));
  OAI21_X1  g0048(.A(G68), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G58), .ZN(new_n250));
  INV_X1    g0050(.A(G68), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g0052(.A(G20), .B1(new_n252), .B2(new_n201), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G159), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n249), .A2(KEYINPUT16), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT16), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT3), .B(G33), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n247), .B1(new_n260), .B2(G20), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n245), .A2(KEYINPUT7), .A3(new_n219), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n251), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n259), .B1(new_n263), .B2(new_n256), .ZN(new_n264));
  NAND3_X1  g0064(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n218), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n258), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G13), .A3(G20), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT68), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT68), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n271), .A2(new_n268), .A3(G13), .A4(G20), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n266), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT8), .B(G58), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n277), .B1(new_n268), .B2(G20), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n270), .A2(new_n272), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n276), .A2(new_n278), .B1(new_n279), .B2(new_n277), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n267), .A2(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT67), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n282), .A2(new_n283), .A3(new_n218), .ZN(new_n284));
  AND2_X1   g0084(.A1(G1), .A2(G13), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G41), .ZN(new_n286));
  AOI21_X1  g0086(.A(KEYINPUT67), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT78), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n268), .B1(G41), .B2(G45), .ZN(new_n290));
  INV_X1    g0090(.A(G274), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AND2_X1   g0092(.A1(new_n290), .A2(G232), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n288), .B(new_n289), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n283), .B1(new_n282), .B2(new_n218), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n285), .A2(KEYINPUT67), .A3(new_n286), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n295), .A2(new_n296), .A3(G232), .A4(new_n290), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n292), .A2(new_n295), .A3(new_n296), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n297), .A2(new_n298), .A3(KEYINPUT78), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n242), .A2(new_n244), .A3(G226), .A4(G1698), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT77), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n260), .A2(KEYINPUT77), .A3(G226), .A4(G1698), .ZN(new_n304));
  NAND2_X1  g0104(.A1(G33), .A2(G87), .ZN(new_n305));
  INV_X1    g0105(.A(G1698), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n260), .A2(G223), .A3(new_n306), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n303), .A2(new_n304), .A3(new_n305), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n285), .A2(new_n286), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n300), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G169), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n294), .A2(new_n299), .B1(new_n308), .B2(new_n310), .ZN(new_n315));
  INV_X1    g0115(.A(G179), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n281), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT18), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT18), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n281), .A2(new_n320), .A3(new_n314), .A4(new_n317), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n280), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n249), .A2(new_n257), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n274), .B1(new_n325), .B2(new_n259), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n324), .B1(new_n326), .B2(new_n258), .ZN(new_n327));
  INV_X1    g0127(.A(G190), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n300), .A2(new_n328), .A3(new_n311), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(G200), .B2(new_n315), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n327), .A2(KEYINPUT17), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT17), .B1(new_n327), .B2(new_n330), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT79), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n300), .A2(new_n328), .A3(new_n311), .ZN(new_n335));
  AOI21_X1  g0135(.A(G200), .B1(new_n300), .B2(new_n311), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n267), .B(new_n280), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT17), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n327), .A2(KEYINPUT17), .A3(new_n330), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT79), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n323), .B1(new_n334), .B2(new_n341), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n342), .A2(KEYINPUT80), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n342), .A2(KEYINPUT80), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n288), .A2(G226), .A3(new_n290), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n345), .A2(new_n298), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n260), .A2(G222), .A3(new_n306), .ZN(new_n347));
  INV_X1    g0147(.A(G77), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n260), .A2(G1698), .ZN(new_n349));
  INV_X1    g0149(.A(G223), .ZN(new_n350));
  OAI221_X1 g0150(.A(new_n347), .B1(new_n348), .B2(new_n260), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n310), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n346), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(G179), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n219), .A2(G33), .ZN(new_n355));
  INV_X1    g0155(.A(G150), .ZN(new_n356));
  INV_X1    g0156(.A(new_n254), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n277), .A2(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G50), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n219), .B1(new_n201), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n266), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n268), .A2(G20), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n273), .A2(new_n274), .A3(G50), .A4(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n279), .A2(new_n359), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n361), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(G169), .B1(new_n346), .B2(new_n352), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n354), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n346), .A2(new_n352), .A3(G190), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n361), .A2(KEYINPUT9), .A3(new_n364), .A4(new_n363), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT71), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT9), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n353), .A2(G200), .B1(new_n373), .B2(new_n365), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n371), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT72), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n353), .A2(G200), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n365), .A2(new_n373), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n378), .A2(new_n379), .A3(new_n370), .A4(new_n369), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT10), .B1(new_n380), .B2(new_n376), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n375), .A2(new_n376), .A3(KEYINPUT10), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n368), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT70), .B1(new_n273), .B2(new_n274), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT70), .ZN(new_n386));
  AOI211_X1 g0186(.A(new_n386), .B(new_n266), .C1(new_n270), .C2(new_n272), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n388), .A2(G68), .A3(new_n362), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT11), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT75), .B1(new_n357), .B2(new_n359), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT75), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n254), .A2(new_n392), .A3(G50), .ZN(new_n393));
  AND2_X1   g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n355), .A2(new_n348), .B1(new_n219), .B2(G68), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n390), .B(new_n266), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n395), .B1(new_n391), .B2(new_n393), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT11), .B1(new_n397), .B2(new_n274), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT76), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n279), .A2(new_n400), .A3(KEYINPUT12), .A4(new_n251), .ZN(new_n401));
  XNOR2_X1  g0201(.A(KEYINPUT76), .B(KEYINPUT12), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n273), .B2(G68), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n389), .A2(new_n399), .A3(new_n401), .A4(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n295), .A2(new_n296), .A3(G238), .A4(new_n290), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n298), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n260), .A2(G232), .A3(G1698), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n260), .A2(G226), .A3(new_n306), .ZN(new_n409));
  AND3_X1   g0209(.A1(KEYINPUT73), .A2(G33), .A3(G97), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT73), .B1(G33), .B2(G97), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n408), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n310), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n407), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT13), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n406), .B1(new_n310), .B2(new_n413), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT13), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n404), .B1(new_n420), .B2(G200), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n418), .B1(new_n407), .B2(new_n414), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT74), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT74), .B1(new_n417), .B2(new_n418), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n424), .A2(new_n425), .A3(G190), .A4(new_n419), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n421), .A2(new_n426), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n407), .A2(new_n414), .A3(new_n418), .ZN(new_n428));
  OAI21_X1  g0228(.A(G169), .B1(new_n428), .B2(new_n422), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT14), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT14), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n420), .A2(new_n431), .A3(G169), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n424), .A2(new_n425), .A3(G179), .A4(new_n419), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n430), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n427), .B1(new_n404), .B2(new_n434), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n288), .A2(new_n290), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n436), .A2(G244), .B1(new_n288), .B2(new_n292), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n260), .A2(G232), .A3(new_n306), .ZN(new_n438));
  INV_X1    g0238(.A(G107), .ZN(new_n439));
  INV_X1    g0239(.A(G238), .ZN(new_n440));
  OAI221_X1 g0240(.A(new_n438), .B1(new_n439), .B2(new_n260), .C1(new_n349), .C2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n310), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(G190), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n388), .A2(G77), .A3(new_n362), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n277), .B1(KEYINPUT69), .B2(new_n357), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(KEYINPUT69), .B2(new_n357), .ZN(new_n448));
  XNOR2_X1  g0248(.A(KEYINPUT15), .B(G87), .ZN(new_n449));
  OAI221_X1 g0249(.A(new_n448), .B1(new_n219), .B2(new_n348), .C1(new_n355), .C2(new_n449), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n450), .A2(new_n266), .B1(new_n348), .B2(new_n279), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n443), .A2(G200), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n445), .A2(new_n446), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n446), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n444), .A2(new_n316), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n443), .A2(new_n313), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n384), .A2(new_n435), .A3(new_n458), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n343), .A2(new_n344), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(G45), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(G1), .ZN(new_n462));
  INV_X1    g0262(.A(G41), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT5), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT5), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G41), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n462), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n467), .A2(new_n295), .A3(new_n296), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n291), .B1(KEYINPUT5), .B2(new_n463), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n295), .A2(new_n296), .A3(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n268), .B(G45), .C1(new_n463), .C2(KEYINPUT5), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT84), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT84), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n462), .A2(new_n473), .A3(new_n466), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n468), .A2(G257), .B1(new_n470), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G283), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n242), .A2(new_n244), .A3(G250), .A4(G1698), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n242), .A2(new_n244), .A3(G244), .A4(new_n306), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT4), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n477), .B(new_n478), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n479), .A2(new_n480), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n310), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(G169), .B1(new_n476), .B2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n467), .A2(new_n295), .A3(G257), .A4(new_n296), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n471), .A2(KEYINPUT84), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n473), .B1(new_n462), .B2(new_n466), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n295), .A2(new_n296), .A3(new_n469), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n485), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n479), .A2(new_n480), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n260), .A2(KEYINPUT4), .A3(G244), .A4(new_n306), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n491), .A2(new_n492), .A3(new_n477), .A4(new_n478), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n490), .B1(new_n310), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n484), .B1(new_n316), .B2(new_n494), .ZN(new_n495));
  XNOR2_X1  g0295(.A(G97), .B(G107), .ZN(new_n496));
  INV_X1    g0296(.A(G97), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT81), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(KEYINPUT6), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT6), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n500), .A2(KEYINPUT81), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n497), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(KEYINPUT81), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n498), .A2(KEYINPUT6), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT82), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n496), .B1(new_n502), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n496), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n507), .A2(new_n509), .A3(KEYINPUT83), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT83), .ZN(new_n511));
  INV_X1    g0311(.A(new_n496), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n513));
  AOI21_X1  g0313(.A(G97), .B1(new_n503), .B2(new_n504), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n511), .B1(new_n515), .B2(new_n508), .ZN(new_n516));
  OAI21_X1  g0316(.A(G20), .B1(new_n510), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(G107), .B1(new_n246), .B2(new_n248), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n254), .A2(G77), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n274), .B1(new_n517), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n279), .A2(G97), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n275), .B1(new_n268), .B2(G33), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n524), .B1(new_n525), .B2(new_n497), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n495), .B1(new_n522), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT83), .B1(new_n507), .B2(new_n509), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n515), .A2(new_n511), .A3(new_n508), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n219), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n266), .B1(new_n531), .B2(new_n520), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n494), .A2(G200), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n476), .A2(new_n483), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n534), .A2(G190), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n532), .B(new_n526), .C1(new_n533), .C2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n242), .A2(new_n244), .A3(new_n219), .A4(G68), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT85), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT85), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n260), .A2(new_n539), .A3(new_n219), .A4(G68), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT19), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n355), .B2(new_n497), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n538), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  NOR3_X1   g0343(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n544));
  OAI21_X1  g0344(.A(KEYINPUT19), .B1(new_n410), .B2(new_n411), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n544), .B1(new_n545), .B2(new_n219), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n266), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n268), .A2(G33), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n276), .A2(G87), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n279), .A2(new_n449), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n547), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n462), .A2(new_n291), .ZN(new_n552));
  INV_X1    g0352(.A(G250), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n461), .B2(G1), .ZN(new_n554));
  AND4_X1   g0354(.A1(new_n295), .A2(new_n552), .A3(new_n296), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n440), .A2(new_n306), .ZN(new_n556));
  INV_X1    g0356(.A(G244), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G1698), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n242), .A2(new_n556), .A3(new_n244), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(G33), .A2(G116), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n309), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n555), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n328), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(G200), .B2(new_n562), .ZN(new_n564));
  INV_X1    g0364(.A(new_n449), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n276), .A2(new_n565), .A3(new_n548), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n547), .A2(new_n566), .A3(new_n550), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n313), .B1(new_n555), .B2(new_n561), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n295), .A2(new_n552), .A3(new_n296), .A4(new_n554), .ZN(new_n569));
  NOR2_X1   g0369(.A1(G238), .A2(G1698), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n570), .B1(new_n557), .B2(G1698), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n571), .A2(new_n260), .B1(G33), .B2(G116), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n316), .B(new_n569), .C1(new_n572), .C2(new_n309), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n551), .A2(new_n564), .B1(new_n567), .B2(new_n574), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n528), .A2(new_n536), .A3(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n242), .A2(new_n244), .A3(new_n219), .A4(G87), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT22), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT22), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n260), .A2(new_n579), .A3(new_n219), .A4(G87), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(G116), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n355), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT23), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n219), .B2(G107), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n439), .A2(KEYINPUT23), .A3(G20), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n583), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT24), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT24), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n581), .A2(new_n590), .A3(new_n587), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n274), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n525), .A2(G107), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n279), .A2(KEYINPUT25), .A3(new_n439), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT25), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n273), .B2(G107), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n592), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT87), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n553), .A2(G1698), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n601), .A2(new_n242), .A3(new_n244), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT86), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n260), .A2(G257), .A3(G1698), .ZN(new_n604));
  NAND2_X1  g0404(.A1(G33), .A2(G294), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT86), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n601), .A2(new_n242), .A3(new_n244), .A4(new_n606), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n603), .A2(new_n604), .A3(new_n605), .A4(new_n607), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n608), .A2(new_n310), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n470), .A2(new_n475), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n467), .A2(new_n295), .A3(G264), .A4(new_n296), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n600), .B1(new_n613), .B2(new_n328), .ZN(new_n614));
  INV_X1    g0414(.A(G200), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n609), .B2(new_n612), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n468), .A2(G264), .B1(new_n470), .B2(new_n475), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n608), .A2(new_n310), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n617), .A2(new_n618), .A3(new_n600), .A4(new_n328), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n599), .B1(new_n614), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(G169), .B1(new_n617), .B2(new_n618), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(new_n316), .B2(new_n613), .ZN(new_n623));
  INV_X1    g0423(.A(new_n591), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n590), .B1(new_n581), .B2(new_n587), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n266), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n626), .A2(new_n593), .A3(new_n597), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n621), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n385), .ZN(new_n630));
  INV_X1    g0430(.A(new_n387), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n582), .B1(new_n268), .B2(G33), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n265), .A2(new_n218), .B1(G20), .B2(new_n582), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n477), .B(new_n219), .C1(G33), .C2(new_n497), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n634), .A2(KEYINPUT20), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT20), .B1(new_n634), .B2(new_n635), .ZN(new_n637));
  OAI22_X1  g0437(.A1(new_n636), .A2(new_n637), .B1(G116), .B2(new_n273), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n633), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(KEYINPUT21), .A2(G169), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n468), .A2(G270), .B1(new_n470), .B2(new_n475), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n242), .A2(new_n244), .A3(G257), .A4(new_n306), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n242), .A2(new_n244), .A3(G264), .A4(G1698), .ZN(new_n644));
  INV_X1    g0444(.A(G303), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n643), .B(new_n644), .C1(new_n645), .C2(new_n260), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n310), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n641), .B1(new_n642), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n288), .A2(G270), .A3(new_n467), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n647), .A2(new_n610), .A3(new_n649), .A4(G179), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n640), .B1(new_n648), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT21), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n647), .A2(new_n610), .A3(new_n649), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(G169), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n638), .B1(new_n388), .B2(new_n632), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n654), .A2(G200), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n658), .B(new_n656), .C1(new_n328), .C2(new_n654), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n652), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  AND4_X1   g0460(.A1(new_n460), .A2(new_n576), .A3(new_n629), .A4(new_n660), .ZN(G372));
  INV_X1    g0461(.A(new_n457), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n421), .A2(new_n426), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n434), .A2(new_n404), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n333), .B1(new_n331), .B2(new_n332), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n339), .A2(KEYINPUT79), .A3(new_n340), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n664), .A2(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n668), .A2(new_n322), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n382), .A2(new_n383), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n368), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n460), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n532), .A2(new_n526), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n673), .A2(new_n575), .A3(KEYINPUT26), .A4(new_n495), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(new_n575), .A3(new_n495), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT90), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT26), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n676), .B1(new_n675), .B2(new_n677), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n674), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n567), .A2(new_n574), .ZN(new_n681));
  XOR2_X1   g0481(.A(new_n681), .B(KEYINPUT89), .Z(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  AND4_X1   g0483(.A1(new_n528), .A2(new_n621), .A3(new_n536), .A4(new_n575), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n652), .A2(new_n657), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n617), .A2(new_n316), .A3(new_n618), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n613), .B2(G169), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT88), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n599), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT88), .B1(new_n623), .B2(new_n627), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n685), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n683), .B1(new_n684), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n680), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n671), .B1(new_n672), .B2(new_n694), .ZN(G369));
  NAND3_X1  g0495(.A1(new_n268), .A2(new_n219), .A3(G13), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G213), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G343), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n660), .B1(new_n656), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n640), .A2(new_n701), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n703), .B1(new_n685), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G330), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n629), .B1(new_n599), .B2(new_n702), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n628), .B2(new_n702), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n689), .A2(new_n690), .A3(new_n701), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n685), .A2(new_n701), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n711), .B1(new_n629), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n710), .A2(new_n713), .ZN(G399));
  INV_X1    g0514(.A(new_n206), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G41), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n544), .A2(new_n582), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n717), .A2(G1), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n221), .B2(new_n717), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT28), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT29), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n685), .A2(new_n628), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n683), .B1(new_n684), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n675), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT92), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n726), .A2(new_n727), .A3(KEYINPUT26), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n675), .A2(new_n677), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(KEYINPUT92), .A3(new_n674), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n725), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n723), .B1(new_n731), .B2(new_n702), .ZN(new_n732));
  AND4_X1   g0532(.A1(new_n657), .A2(new_n652), .A3(new_n659), .A4(new_n702), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n576), .A2(new_n629), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n617), .A2(new_n618), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n559), .A2(new_n560), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n310), .ZN(new_n737));
  AOI21_X1  g0537(.A(G179), .B1(new_n737), .B2(new_n569), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n534), .A2(new_n735), .A3(new_n654), .A4(new_n738), .ZN(new_n739));
  AND3_X1   g0539(.A1(new_n647), .A2(new_n610), .A3(new_n649), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n737), .A2(new_n569), .A3(new_n611), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n740), .A2(G179), .A3(new_n742), .A4(new_n618), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n494), .A2(KEYINPUT30), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n739), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n618), .A2(new_n562), .A3(new_n611), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n650), .ZN(new_n747));
  AOI21_X1  g0547(.A(KEYINPUT30), .B1(new_n747), .B2(new_n494), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n701), .B1(new_n745), .B2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT31), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(KEYINPUT91), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT91), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n749), .A2(new_n753), .A3(new_n750), .ZN(new_n754));
  OAI211_X1 g0554(.A(KEYINPUT31), .B(new_n701), .C1(new_n745), .C2(new_n748), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n734), .A2(new_n752), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G330), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI211_X1 g0558(.A(KEYINPUT29), .B(new_n701), .C1(new_n680), .C2(new_n692), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n732), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n722), .B1(new_n760), .B2(G1), .ZN(G364));
  NAND2_X1  g0561(.A1(new_n219), .A2(G13), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n268), .B1(new_n763), .B2(G45), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n716), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n707), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(G330), .B2(new_n705), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n260), .A2(new_n206), .ZN(new_n769));
  INV_X1    g0569(.A(G355), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n769), .A2(new_n770), .B1(G116), .B2(new_n206), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n236), .A2(G45), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n715), .A2(new_n260), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n774), .B1(new_n461), .B2(new_n222), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n771), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G13), .A2(G33), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n218), .B1(G20), .B2(new_n313), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n766), .B1(new_n776), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n219), .A2(new_n316), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n786), .A2(new_n328), .A3(G200), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G322), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n786), .A2(G190), .A3(G200), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G311), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n788), .A2(new_n789), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR4_X1   g0593(.A1(new_n219), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n260), .B(new_n793), .C1(G329), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n785), .A2(G200), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(G190), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  OR2_X1    g0598(.A1(KEYINPUT33), .A2(G317), .ZN(new_n799));
  NAND2_X1  g0599(.A1(KEYINPUT33), .A2(G317), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n796), .A2(new_n328), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G326), .ZN(new_n804));
  INV_X1    g0604(.A(G294), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n328), .A2(G179), .A3(G200), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n219), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n803), .A2(new_n804), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n801), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n316), .A2(G200), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT95), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NOR3_X1   g0612(.A1(new_n812), .A2(new_n219), .A3(G190), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G283), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n812), .A2(new_n219), .A3(new_n328), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G303), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n795), .A2(new_n809), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  AOI22_X1  g0617(.A1(G58), .A2(new_n787), .B1(new_n790), .B2(G77), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT93), .Z(new_n819));
  INV_X1    g0619(.A(new_n813), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(new_n439), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n815), .A2(G87), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n819), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n794), .ZN(new_n825));
  XOR2_X1   g0625(.A(KEYINPUT94), .B(G159), .Z(new_n826));
  NOR2_X1   g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT32), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n359), .A2(new_n803), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n245), .B(new_n829), .C1(new_n828), .C2(new_n827), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n798), .A2(new_n251), .B1(new_n497), .B2(new_n807), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n831), .A2(KEYINPUT96), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(KEYINPUT96), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n830), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n817), .B1(new_n824), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n784), .B1(new_n835), .B2(new_n781), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n705), .B2(new_n780), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n768), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(G396));
  AND2_X1   g0639(.A1(new_n458), .A2(new_n702), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n693), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n694), .A2(new_n701), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n457), .A2(new_n701), .ZN(new_n843));
  INV_X1    g0643(.A(new_n454), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n453), .B1(new_n844), .B2(new_n702), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n843), .B1(new_n845), .B2(new_n457), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n841), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n847), .A2(new_n757), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT98), .Z(new_n849));
  AOI21_X1  g0649(.A(new_n766), .B1(new_n847), .B2(new_n757), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n766), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n781), .A2(new_n777), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n852), .B1(new_n348), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n826), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n790), .A2(new_n855), .B1(new_n787), .B2(G143), .ZN(new_n856));
  INV_X1    g0656(.A(G137), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n856), .B1(new_n857), .B2(new_n803), .C1(new_n356), .C2(new_n798), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT34), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n858), .A2(new_n859), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n813), .A2(G68), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n815), .A2(G50), .ZN(new_n863));
  INV_X1    g0663(.A(new_n807), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(G58), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n245), .B1(new_n794), .B2(G132), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n862), .A2(new_n863), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n861), .A2(new_n867), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n245), .B1(new_n825), .B2(new_n792), .C1(new_n788), .C2(new_n805), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n813), .A2(G87), .ZN(new_n870));
  INV_X1    g0670(.A(new_n815), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n870), .B1(new_n871), .B2(new_n439), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n869), .B(new_n872), .C1(G97), .C2(new_n864), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n790), .A2(G116), .B1(new_n802), .B2(G303), .ZN(new_n874));
  INV_X1    g0674(.A(G283), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n874), .B1(new_n875), .B2(new_n798), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n876), .B(KEYINPUT97), .Z(new_n877));
  AOI22_X1  g0677(.A1(new_n860), .A2(new_n868), .B1(new_n873), .B2(new_n877), .ZN(new_n878));
  OAI221_X1 g0678(.A(new_n854), .B1(new_n782), .B2(new_n878), .C1(new_n846), .C2(new_n778), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n851), .A2(new_n879), .ZN(G384));
  INV_X1    g0680(.A(G330), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT99), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n327), .B2(new_n699), .ZN(new_n883));
  INV_X1    g0683(.A(new_n699), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n281), .A2(KEYINPUT99), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n342), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n318), .A2(new_n337), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT37), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n889), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT100), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(new_n281), .B2(new_n884), .ZN(new_n893));
  AOI211_X1 g0693(.A(KEYINPUT100), .B(new_n699), .C1(new_n267), .C2(new_n280), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT37), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n891), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n890), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT38), .B1(new_n888), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n666), .A2(new_n667), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n886), .B1(new_n900), .B2(new_n323), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n896), .B1(new_n891), .B2(new_n886), .ZN(new_n902));
  NOR4_X1   g0702(.A1(new_n889), .A2(new_n893), .A3(new_n894), .A4(KEYINPUT37), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT38), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT101), .B1(new_n899), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT38), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n902), .A2(new_n903), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n907), .B1(new_n901), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n888), .A2(KEYINPUT38), .A3(new_n898), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT101), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n906), .A2(new_n912), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n404), .B(new_n701), .C1(new_n427), .C2(new_n434), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n404), .A2(new_n701), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n665), .A2(new_n663), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n846), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n660), .A2(new_n621), .A3(new_n628), .A4(new_n702), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n528), .A2(new_n536), .A3(new_n575), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n751), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n755), .A2(KEYINPUT103), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT30), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n743), .B2(new_n534), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n534), .A2(new_n923), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n747), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n924), .A2(new_n926), .A3(new_n739), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT103), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n927), .A2(new_n928), .A3(KEYINPUT31), .A4(new_n701), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n922), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n921), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n918), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT40), .B1(new_n913), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT102), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n901), .B2(new_n904), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n888), .A2(new_n898), .A3(KEYINPUT102), .A4(KEYINPUT38), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n896), .B1(new_n891), .B2(new_n895), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n339), .A2(new_n340), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n322), .A2(new_n938), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n903), .A2(new_n937), .B1(new_n939), .B2(new_n895), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n907), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n935), .A2(new_n936), .A3(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT40), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n918), .A2(new_n931), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n933), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n672), .A2(new_n931), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n881), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n945), .B2(new_n946), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n843), .B1(new_n693), .B2(new_n840), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n913), .A2(new_n917), .A3(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(KEYINPUT39), .B1(new_n899), .B2(new_n905), .ZN(new_n952));
  AOI21_X1  g0752(.A(KEYINPUT39), .B1(new_n940), .B2(new_n907), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(new_n935), .A3(new_n936), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n665), .A2(new_n701), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n322), .A2(new_n699), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n951), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n460), .B1(new_n759), .B2(new_n732), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n671), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n959), .B(new_n961), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n948), .A2(new_n962), .B1(G1), .B2(new_n762), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n962), .B2(new_n948), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n220), .A2(G116), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n529), .A2(new_n530), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n965), .B1(new_n966), .B2(KEYINPUT35), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(KEYINPUT35), .B2(new_n966), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(KEYINPUT36), .Z(new_n969));
  OR3_X1    g0769(.A1(new_n221), .A2(new_n348), .A3(new_n252), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n359), .A2(G68), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n268), .B(G13), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n964), .A2(new_n973), .ZN(G367));
  NAND2_X1  g0774(.A1(new_n673), .A2(new_n701), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n975), .A2(new_n528), .A3(new_n536), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n673), .A2(new_n495), .A3(new_n701), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n629), .A2(new_n712), .ZN(new_n980));
  OAI21_X1  g0780(.A(KEYINPUT42), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n528), .B1(new_n976), .B2(new_n628), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n702), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NOR3_X1   g0784(.A1(new_n979), .A2(KEYINPUT42), .A3(new_n980), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT43), .ZN(new_n986));
  NOR3_X1   g0786(.A1(new_n682), .A2(new_n551), .A3(new_n702), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n551), .A2(new_n702), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n987), .B1(new_n575), .B2(new_n988), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n984), .A2(new_n985), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n986), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n990), .B(new_n991), .Z(new_n992));
  NOR2_X1   g0792(.A1(new_n710), .A2(new_n979), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n992), .B(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n716), .B(KEYINPUT41), .Z(new_n995));
  NAND2_X1  g0795(.A1(new_n713), .A2(new_n978), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT45), .Z(new_n997));
  NOR2_X1   g0797(.A1(new_n713), .A2(new_n978), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT44), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(new_n710), .Z(new_n1001));
  OAI21_X1  g0801(.A(new_n980), .B1(new_n709), .B2(new_n712), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(new_n707), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n760), .A2(new_n1003), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n995), .B1(new_n1005), .B2(new_n760), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n994), .B1(new_n1006), .B2(new_n765), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n783), .B1(new_n715), .B2(new_n565), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n231), .A2(new_n773), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n852), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n807), .A2(new_n251), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(new_n797), .B2(new_n855), .ZN(new_n1012));
  INV_X1    g0812(.A(G143), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1012), .B1(new_n1013), .B2(new_n803), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n813), .A2(G77), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n245), .B1(new_n787), .B2(G150), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1015), .B(new_n1016), .C1(new_n359), .C2(new_n791), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n871), .A2(new_n250), .B1(new_n857), .B2(new_n825), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1014), .B(new_n1017), .C1(KEYINPUT104), .C2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(KEYINPUT104), .B2(new_n1018), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT105), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n820), .A2(new_n497), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n787), .A2(G303), .B1(G317), .B2(new_n794), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1023), .B(new_n245), .C1(new_n875), .C2(new_n791), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G107), .A2(new_n864), .B1(new_n797), .B2(G294), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(new_n792), .C2(new_n803), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n815), .A2(G116), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT46), .Z(new_n1029));
  OAI21_X1  g0829(.A(new_n1021), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT47), .Z(new_n1031));
  OAI21_X1  g0831(.A(new_n1010), .B1(new_n1031), .B2(new_n782), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1033), .A2(KEYINPUT106), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n989), .A2(new_n779), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1033), .A2(KEYINPUT106), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1007), .A2(new_n1037), .ZN(G387));
  OR2_X1    g0838(.A1(new_n709), .A2(new_n780), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n719), .A2(new_n769), .B1(G107), .B2(new_n206), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n228), .A2(G45), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT107), .Z(new_n1042));
  NOR2_X1   g0842(.A1(new_n277), .A2(G50), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT50), .ZN(new_n1044));
  AOI211_X1 g0844(.A(G45), .B(new_n718), .C1(G68), .C2(G77), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n774), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1040), .B1(new_n1042), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n766), .B1(new_n1047), .B2(new_n783), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G303), .A2(new_n790), .B1(new_n787), .B2(G317), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n792), .B2(new_n798), .C1(new_n789), .C2(new_n803), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT48), .Z(new_n1051));
  AOI22_X1  g0851(.A1(new_n815), .A2(G294), .B1(new_n864), .B2(G283), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT108), .Z(new_n1053));
  NOR2_X1   g0853(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1054), .A2(KEYINPUT49), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n245), .B1(new_n825), .B2(new_n804), .C1(new_n820), .C2(new_n582), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(KEYINPUT49), .B2(new_n1054), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n788), .A2(new_n359), .B1(new_n825), .B2(new_n356), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n245), .B(new_n1059), .C1(G68), .C2(new_n790), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1022), .ZN(new_n1061));
  INV_X1    g0861(.A(G159), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n1062), .A2(new_n803), .B1(new_n798), .B2(new_n277), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n807), .A2(new_n449), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n815), .A2(G77), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1060), .A2(new_n1061), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1058), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1048), .B1(new_n1068), .B2(new_n781), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1039), .A2(new_n1069), .B1(new_n1003), .B2(new_n765), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1004), .A2(new_n716), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n760), .A2(new_n1003), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(G393));
  NOR2_X1   g0873(.A1(new_n978), .A2(new_n780), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT109), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n783), .B1(G97), .B2(new_n715), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n239), .A2(new_n773), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n852), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n822), .B1(new_n875), .B2(new_n871), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n245), .B1(new_n789), .B2(new_n825), .C1(new_n791), .C2(new_n805), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n798), .A2(new_n645), .B1(new_n582), .B2(new_n807), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n787), .A2(G311), .B1(new_n802), .B2(G317), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1083), .B(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n870), .B1(new_n871), .B2(new_n251), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n260), .B1(new_n1013), .B2(new_n825), .C1(new_n791), .C2(new_n277), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n807), .A2(new_n348), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n798), .A2(new_n359), .ZN(new_n1089));
  NOR4_X1   g0889(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n787), .A2(G159), .B1(new_n802), .B2(G150), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT51), .Z(new_n1092));
  AOI22_X1  g0892(.A1(new_n1082), .A2(new_n1085), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1075), .B(new_n1078), .C1(new_n782), .C2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1005), .A2(new_n716), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n1094), .B1(new_n764), .B2(new_n1001), .C1(new_n1095), .C2(new_n1097), .ZN(G390));
  INV_X1    g0898(.A(new_n956), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n917), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1099), .B1(new_n949), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1101), .A2(new_n952), .A3(new_n954), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n845), .A2(new_n457), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n730), .A2(new_n728), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n724), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n528), .A2(new_n621), .A3(new_n536), .A4(new_n575), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n682), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n702), .B(new_n1103), .C1(new_n1104), .C2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n843), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n917), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1111), .A2(new_n942), .A3(new_n1099), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1102), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(G330), .B1(new_n921), .B2(new_n930), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n918), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n756), .A2(G330), .A3(new_n846), .A4(new_n917), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1102), .A2(new_n1112), .A3(new_n1117), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n765), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n791), .A2(new_n497), .B1(new_n825), .B2(new_n805), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n260), .B(new_n1121), .C1(G116), .C2(new_n787), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1122), .A2(new_n823), .A3(new_n862), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1088), .B1(G283), .B2(new_n802), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n439), .B2(new_n798), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n815), .A2(G150), .ZN(new_n1126));
  XOR2_X1   g0926(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n1127));
  XNOR2_X1  g0927(.A(new_n1126), .B(new_n1127), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n798), .A2(new_n857), .B1(new_n1062), .B2(new_n807), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(G128), .B2(new_n802), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n813), .A2(G50), .ZN(new_n1131));
  XOR2_X1   g0931(.A(KEYINPUT54), .B(G143), .Z(new_n1132));
  AOI21_X1  g0932(.A(new_n245), .B1(new_n790), .B2(new_n1132), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n787), .A2(G132), .B1(G125), .B2(new_n794), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1130), .A2(new_n1131), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n1123), .A2(new_n1125), .B1(new_n1128), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT113), .ZN(new_n1137));
  OR2_X1    g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n782), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n852), .B1(new_n277), .B2(new_n853), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1140), .B(new_n1141), .C1(new_n955), .C2(new_n778), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1120), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1114), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n460), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n960), .A2(new_n671), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT111), .ZN(new_n1147));
  OAI211_X1 g0947(.A(G330), .B(new_n846), .C1(new_n921), .C2(new_n930), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n1100), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n1117), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1147), .B1(new_n1150), .B2(new_n1110), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1152), .A2(KEYINPUT111), .A3(new_n1117), .A4(new_n1149), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n917), .B1(new_n758), .B2(new_n846), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n950), .B1(new_n1155), .B2(new_n1115), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1146), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1119), .A2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1158), .A2(new_n717), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1157), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1143), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(G378));
  INV_X1    g0962(.A(new_n959), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n368), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n371), .A2(KEYINPUT72), .A3(new_n374), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n376), .A2(new_n375), .B1(new_n1165), .B2(KEYINPUT10), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n383), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1164), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n366), .A2(new_n699), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1169), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n384), .A2(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NOR3_X1   g0974(.A1(new_n1170), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n384), .A2(new_n1171), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1173), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1175), .A2(new_n1178), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n899), .A2(new_n905), .A3(KEYINPUT101), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n911), .B1(new_n909), .B2(new_n910), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n932), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n943), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n881), .B1(new_n942), .B2(new_n944), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1179), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT119), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1174), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1176), .A2(new_n1177), .A3(new_n1173), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1188), .A2(KEYINPUT119), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1187), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n932), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n906), .B2(new_n912), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1191), .B(new_n1184), .C1(new_n1193), .C2(KEYINPUT40), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1163), .B1(new_n1185), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1179), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1184), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1197), .B1(new_n933), .B2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1199), .A2(new_n959), .A3(new_n1194), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1146), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1196), .A2(new_n1200), .B1(new_n1201), .B2(new_n1160), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n716), .B1(new_n1202), .B2(KEYINPUT57), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1196), .A2(new_n1200), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1160), .A2(new_n1201), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n1204), .A2(KEYINPUT57), .A3(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1203), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT121), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n764), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n853), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n766), .B1(G50), .B2(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n260), .A2(G41), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1212), .B1(new_n875), .B2(new_n825), .C1(new_n791), .C2(new_n449), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n788), .A2(new_n439), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1011), .B(new_n1213), .C1(KEYINPUT114), .C2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n813), .A2(G58), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1215), .A2(new_n1066), .A3(new_n1216), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G97), .A2(new_n797), .B1(new_n802), .B2(G116), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1217), .B(new_n1218), .C1(KEYINPUT114), .C2(new_n1214), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n1219), .B(KEYINPUT115), .Z(new_n1220));
  XNOR2_X1  g1020(.A(KEYINPUT116), .B(KEYINPUT58), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n815), .A2(new_n1132), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n797), .A2(G132), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(G128), .A2(new_n787), .B1(new_n790), .B2(G137), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(G150), .A2(new_n864), .B1(new_n802), .B2(G125), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  XOR2_X1   g1028(.A(new_n1228), .B(KEYINPUT59), .Z(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  OR2_X1    g1030(.A1(new_n1230), .A2(KEYINPUT117), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(KEYINPUT117), .ZN(new_n1232));
  XOR2_X1   g1032(.A(KEYINPUT118), .B(G124), .Z(new_n1233));
  OAI211_X1 g1033(.A(new_n241), .B(new_n463), .C1(new_n825), .C2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(new_n813), .B2(new_n855), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1231), .A2(new_n1232), .A3(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1212), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1237), .B(new_n359), .C1(G33), .C2(G41), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1222), .A2(new_n1223), .A3(new_n1236), .A4(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1211), .B1(new_n1239), .B2(new_n781), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1191), .A2(new_n777), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  XOR2_X1   g1042(.A(new_n1242), .B(KEYINPUT120), .Z(new_n1243));
  OAI21_X1  g1043(.A(new_n1208), .B1(new_n1209), .B2(new_n1243), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n1199), .A2(new_n959), .A3(new_n1194), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n959), .B1(new_n1199), .B2(new_n1194), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n765), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1242), .B(KEYINPUT120), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(KEYINPUT121), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1244), .A2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(KEYINPUT122), .B1(new_n1207), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT57), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1202), .A2(KEYINPUT57), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(new_n716), .A3(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT122), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1256), .A2(new_n1257), .A3(new_n1244), .A4(new_n1249), .ZN(new_n1258));
  AND2_X1   g1058(.A1(new_n1251), .A2(new_n1258), .ZN(G375));
  NAND2_X1  g1059(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1146), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n995), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1157), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n766), .B1(G68), .B2(new_n1210), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1064), .B1(G294), .B2(new_n802), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(new_n582), .B2(new_n798), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n815), .A2(G97), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n260), .B1(new_n790), .B2(G107), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n787), .A2(G283), .B1(G303), .B2(new_n794), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1015), .A2(new_n1269), .A3(new_n1270), .A4(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n815), .A2(G159), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n245), .B1(new_n787), .B2(G137), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n790), .A2(G150), .B1(G128), .B2(new_n794), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1216), .A2(new_n1273), .A3(new_n1274), .A4(new_n1275), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(G132), .A2(new_n802), .B1(new_n797), .B2(new_n1132), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(new_n359), .B2(new_n807), .ZN(new_n1278));
  OAI22_X1  g1078(.A1(new_n1268), .A2(new_n1272), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1266), .B1(new_n1279), .B2(new_n781), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n917), .B2(new_n778), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n1261), .B2(new_n764), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1265), .A2(new_n1283), .ZN(G381));
  NOR4_X1   g1084(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1285));
  INV_X1    g1085(.A(G387), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  OR4_X1    g1087(.A1(G378), .A2(G375), .A3(new_n1287), .A4(G381), .ZN(G407));
  NAND2_X1  g1088(.A1(new_n700), .A2(G213), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1161), .A2(new_n1290), .ZN(new_n1291));
  OAI211_X1 g1091(.A(G407), .B(G213), .C1(G375), .C2(new_n1291), .ZN(G409));
  INV_X1    g1092(.A(new_n1242), .ZN(new_n1293));
  OAI21_X1  g1093(.A(KEYINPUT124), .B1(new_n1209), .B2(new_n1293), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1205), .B(new_n1263), .C1(new_n1245), .C2(new_n1246), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(KEYINPUT123), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT124), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1247), .A2(new_n1297), .A3(new_n1242), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT123), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1204), .A2(new_n1299), .A3(new_n1263), .A4(new_n1205), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1294), .A2(new_n1296), .A3(new_n1298), .A4(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1161), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(KEYINPUT125), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT125), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1301), .A2(new_n1304), .A3(new_n1161), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1256), .A2(G378), .A3(new_n1244), .A4(new_n1249), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1303), .A2(new_n1305), .A3(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1264), .A2(KEYINPUT60), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1262), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1261), .A2(KEYINPUT60), .A3(new_n1146), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1309), .A2(new_n716), .A3(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1283), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1312), .A2(new_n851), .A3(new_n879), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1311), .A2(G384), .A3(new_n1283), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1307), .A2(new_n1289), .A3(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(KEYINPUT62), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT61), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1290), .A2(G2897), .ZN(new_n1320));
  XNOR2_X1  g1120(.A(new_n1315), .B(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1305), .ZN(new_n1322));
  NOR3_X1   g1122(.A1(new_n1207), .A2(new_n1250), .A3(new_n1161), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1304), .B1(new_n1301), .B2(new_n1161), .ZN(new_n1324));
  NOR3_X1   g1124(.A1(new_n1322), .A2(new_n1323), .A3(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1321), .B1(new_n1325), .B2(new_n1290), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT62), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1307), .A2(new_n1327), .A3(new_n1289), .A4(new_n1316), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1318), .A2(new_n1319), .A3(new_n1326), .A4(new_n1328), .ZN(new_n1329));
  XNOR2_X1  g1129(.A(G393), .B(new_n838), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1330), .B1(G387), .B2(KEYINPUT126), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1331), .B1(G387), .B2(new_n1330), .ZN(new_n1332));
  INV_X1    g1132(.A(G390), .ZN(new_n1333));
  XNOR2_X1  g1133(.A(new_n1332), .B(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1329), .A2(new_n1334), .ZN(new_n1335));
  XNOR2_X1  g1135(.A(new_n1332), .B(G390), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1307), .A2(new_n1289), .ZN(new_n1337));
  AOI21_X1  g1137(.A(KEYINPUT61), .B1(new_n1337), .B2(new_n1321), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT63), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1317), .A2(new_n1339), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1307), .A2(KEYINPUT63), .A3(new_n1289), .A4(new_n1316), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1336), .A2(new_n1338), .A3(new_n1340), .A4(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1335), .A2(new_n1342), .ZN(G405));
  NAND3_X1  g1143(.A1(new_n1251), .A2(new_n1258), .A3(new_n1161), .ZN(new_n1344));
  OR2_X1    g1144(.A1(new_n1344), .A2(KEYINPUT127), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1344), .A2(KEYINPUT127), .A3(new_n1306), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1315), .B1(new_n1345), .B2(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1347), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1345), .A2(new_n1315), .A3(new_n1346), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1348), .A2(new_n1334), .A3(new_n1349), .ZN(new_n1350));
  AND3_X1   g1150(.A1(new_n1345), .A2(new_n1315), .A3(new_n1346), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1336), .B1(new_n1351), .B2(new_n1347), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1350), .A2(new_n1352), .ZN(G402));
endmodule


