//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 1 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1239, new_n1240, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1307, new_n1308;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  INV_X1    g0009(.A(G77), .ZN(new_n210));
  INV_X1    g0010(.A(G244), .ZN(new_n211));
  INV_X1    g0011(.A(G264), .ZN(new_n212));
  OAI22_X1  g0012(.A1(new_n210), .A2(new_n211), .B1(new_n206), .B2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT64), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n213), .B(new_n215), .C1(G50), .C2(G226), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G116), .A2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G58), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n216), .B(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n209), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n209), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT0), .Z(new_n228));
  OAI21_X1  g0028(.A(G50), .B1(G58), .B2(G68), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NOR3_X1   g0032(.A1(new_n225), .A2(new_n228), .A3(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n219), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G58), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  NAND2_X1  g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(G1), .A3(G13), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT3), .B(G33), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n252), .A2(G238), .A3(G1698), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n253), .B1(new_n206), .B2(new_n252), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NOR3_X1   g0059(.A1(new_n259), .A2(new_n219), .A3(G1698), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n251), .B1(new_n254), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G1), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n262), .B1(G41), .B2(G45), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  OR2_X1    g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT65), .ZN(new_n266));
  AND3_X1   g0066(.A1(new_n250), .A2(new_n266), .A3(new_n263), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n266), .B1(new_n250), .B2(new_n263), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G244), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n261), .A2(new_n265), .A3(new_n270), .ZN(new_n271));
  OR2_X1    g0071(.A1(new_n271), .A2(G179), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT8), .B(G58), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G20), .A2(G33), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n274), .A2(new_n275), .B1(G20), .B2(G77), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n230), .A2(G33), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT15), .B(G87), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n231), .ZN(new_n281));
  INV_X1    g0081(.A(G13), .ZN(new_n282));
  NOR3_X1   g0082(.A1(new_n282), .A2(new_n230), .A3(G1), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n279), .A2(new_n281), .B1(new_n210), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n281), .B1(new_n262), .B2(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n284), .B1(new_n210), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G169), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n271), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n272), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G97), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G226), .A2(G1698), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n294), .B1(new_n219), .B2(G1698), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n293), .B1(new_n295), .B2(new_n252), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n265), .B1(new_n296), .B2(new_n250), .ZN(new_n297));
  NOR3_X1   g0097(.A1(new_n267), .A2(new_n268), .A3(new_n222), .ZN(new_n298));
  OAI21_X1  g0098(.A(KEYINPUT13), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n268), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n250), .A2(new_n266), .A3(new_n263), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n300), .A2(G238), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n219), .A2(G1698), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(G226), .B2(G1698), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n292), .B1(new_n304), .B2(new_n259), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n251), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT13), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n302), .A2(new_n306), .A3(new_n307), .A4(new_n265), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n299), .A2(KEYINPUT66), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT66), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n310), .B(KEYINPUT13), .C1(new_n297), .C2(new_n298), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(G169), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT69), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n309), .A2(KEYINPUT69), .A3(G169), .A4(new_n311), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n314), .A2(KEYINPUT14), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT70), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n299), .B(KEYINPUT67), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT68), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n308), .B(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n319), .A2(G179), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT14), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n309), .A2(new_n323), .A3(G169), .A4(new_n311), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n314), .A2(KEYINPUT70), .A3(KEYINPUT14), .A4(new_n315), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n318), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n275), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n328), .A2(new_n202), .B1(new_n230), .B2(G68), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n277), .A2(new_n210), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n281), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT11), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n283), .ZN(new_n334));
  NOR3_X1   g0134(.A1(new_n334), .A2(KEYINPUT12), .A3(G68), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT12), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n336), .B1(new_n283), .B2(new_n221), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n335), .A2(new_n337), .B1(new_n286), .B2(new_n221), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n291), .B1(new_n327), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n319), .A2(G190), .A3(new_n321), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n309), .A2(G200), .A3(new_n311), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(new_n343), .A3(new_n339), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT7), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n230), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT72), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT71), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n350), .A2(KEYINPUT3), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n257), .A2(KEYINPUT71), .ZN(new_n352));
  OAI21_X1  g0152(.A(G33), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n349), .B1(new_n353), .B2(new_n256), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n257), .A2(KEYINPUT71), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n350), .A2(KEYINPUT3), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n255), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n257), .A2(G33), .ZN(new_n358));
  NOR3_X1   g0158(.A1(new_n357), .A2(KEYINPUT72), .A3(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n348), .B1(new_n354), .B2(new_n359), .ZN(new_n360));
  XNOR2_X1  g0160(.A(KEYINPUT71), .B(KEYINPUT3), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n256), .B1(new_n361), .B2(new_n255), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n346), .B1(new_n362), .B2(new_n230), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n360), .A2(G68), .A3(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n218), .A2(new_n221), .ZN(new_n366));
  OAI21_X1  g0166(.A(G20), .B1(new_n366), .B2(new_n201), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n275), .A2(G159), .ZN(new_n368));
  AND3_X1   g0168(.A1(new_n367), .A2(KEYINPUT73), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(KEYINPUT73), .B1(new_n367), .B2(new_n368), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n365), .A2(KEYINPUT16), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n259), .A2(new_n348), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n355), .A2(new_n356), .A3(new_n255), .ZN(new_n374));
  AOI21_X1  g0174(.A(G20), .B1(new_n374), .B2(new_n258), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n373), .B1(new_n375), .B2(new_n346), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n371), .B1(new_n221), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT16), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n372), .A2(new_n379), .A3(new_n281), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n274), .A2(new_n283), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n381), .B1(new_n286), .B2(new_n274), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n250), .A2(new_n263), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n265), .B1(new_n384), .B2(new_n219), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT74), .ZN(new_n386));
  XNOR2_X1  g0186(.A(new_n385), .B(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(G223), .A2(G1698), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G1698), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n390), .A2(G226), .ZN(new_n391));
  AND4_X1   g0191(.A1(new_n256), .A2(new_n353), .A3(new_n389), .A4(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(G87), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n255), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n251), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G190), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n387), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G200), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n357), .A2(new_n358), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n399), .A2(new_n389), .A3(new_n391), .ZN(new_n400));
  INV_X1    g0200(.A(new_n394), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n250), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n398), .B1(new_n402), .B2(new_n385), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n397), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n380), .A2(new_n383), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT75), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT17), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n406), .A2(new_n407), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n408), .B1(new_n405), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n380), .A2(new_n383), .ZN(new_n413));
  INV_X1    g0213(.A(G179), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n387), .A2(new_n395), .A3(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n288), .B1(new_n402), .B2(new_n385), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(KEYINPUT18), .B1(new_n413), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT18), .ZN(new_n420));
  AOI211_X1 g0220(.A(new_n420), .B(new_n417), .C1(new_n380), .C2(new_n383), .ZN(new_n421));
  OAI22_X1  g0221(.A1(new_n410), .A2(new_n412), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n285), .A2(G50), .ZN(new_n424));
  INV_X1    g0224(.A(G150), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n273), .A2(new_n277), .B1(new_n425), .B2(new_n328), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n426), .B1(G20), .B2(new_n203), .ZN(new_n427));
  INV_X1    g0227(.A(new_n281), .ZN(new_n428));
  OAI221_X1 g0228(.A(new_n424), .B1(G50), .B2(new_n334), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT9), .ZN(new_n430));
  NOR2_X1   g0230(.A1(G222), .A2(G1698), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n390), .A2(G223), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n252), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n433), .B(new_n251), .C1(G77), .C2(new_n252), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n265), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n435), .B1(G226), .B2(new_n269), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(G190), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n430), .B(new_n437), .C1(new_n398), .C2(new_n436), .ZN(new_n438));
  XNOR2_X1  g0238(.A(new_n438), .B(KEYINPUT10), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n436), .A2(new_n414), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n440), .B(new_n429), .C1(G169), .C2(new_n436), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n287), .B1(G200), .B2(new_n271), .ZN(new_n442));
  OR2_X1    g0242(.A1(new_n271), .A2(new_n396), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n423), .A2(new_n439), .A3(new_n441), .A4(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT78), .ZN(new_n447));
  NOR4_X1   g0247(.A1(new_n357), .A2(new_n211), .A3(G1698), .A4(new_n358), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n447), .B1(new_n448), .B2(KEYINPUT4), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n252), .A2(KEYINPUT4), .A3(G244), .A4(new_n390), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G283), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n252), .A2(G250), .A3(G1698), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n353), .A2(G244), .A3(new_n390), .A4(new_n256), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT4), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n454), .A2(KEYINPUT78), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n449), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n251), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n262), .A2(G45), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(new_n264), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT5), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G41), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT79), .B1(new_n461), .B2(G41), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT79), .ZN(new_n464));
  INV_X1    g0264(.A(G41), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT5), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n460), .A2(new_n462), .A3(new_n463), .A4(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n462), .A2(new_n262), .A3(G45), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n461), .A2(G41), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(new_n251), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G257), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n458), .A2(new_n467), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT80), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n472), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n476), .B1(new_n457), .B2(new_n251), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n477), .A2(KEYINPUT80), .A3(new_n467), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n475), .A2(G200), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n275), .A2(G77), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT76), .B(KEYINPUT6), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n205), .A2(G107), .ZN(new_n482));
  OR2_X1    g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G97), .A2(G107), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n481), .A2(new_n207), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n483), .A2(G20), .A3(new_n485), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n480), .B(new_n486), .C1(new_n376), .C2(new_n206), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n281), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n334), .B(new_n428), .C1(G1), .C2(new_n255), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G97), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n283), .A2(new_n205), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n488), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT77), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n487), .A2(new_n281), .B1(new_n205), .B2(new_n283), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n496), .A2(KEYINPUT77), .A3(new_n491), .ZN(new_n497));
  INV_X1    g0297(.A(new_n467), .ZN(new_n498));
  AOI211_X1 g0298(.A(new_n498), .B(new_n476), .C1(new_n457), .C2(new_n251), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n495), .A2(new_n497), .B1(new_n499), .B2(G190), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n477), .A2(G179), .A3(new_n467), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n501), .B1(new_n499), .B2(new_n288), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n479), .A2(new_n500), .B1(new_n502), .B2(new_n493), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n393), .A2(G20), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n256), .B(new_n504), .C1(new_n361), .C2(new_n255), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT84), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT84), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n353), .A2(new_n507), .A3(new_n256), .A4(new_n504), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n506), .A2(KEYINPUT22), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT22), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n252), .A2(new_n510), .A3(new_n504), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n230), .A2(G33), .A3(G116), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n230), .A2(G107), .ZN(new_n514));
  XNOR2_X1  g0314(.A(new_n514), .B(KEYINPUT23), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n512), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT24), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n512), .A2(KEYINPUT24), .A3(new_n513), .A4(new_n515), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(new_n281), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n490), .A2(G107), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n334), .A2(G107), .ZN(new_n523));
  XOR2_X1   g0323(.A(KEYINPUT85), .B(KEYINPUT25), .Z(new_n524));
  INV_X1    g0324(.A(KEYINPUT86), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n525), .ZN(new_n527));
  MUX2_X1   g0327(.A(new_n523), .B(new_n526), .S(new_n527), .Z(new_n528));
  INV_X1    g0328(.A(G294), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n255), .A2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  OR2_X1    g0331(.A1(G250), .A2(G1698), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n353), .A2(new_n256), .A3(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n390), .A2(G257), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n498), .B1(new_n535), .B2(new_n251), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n471), .A2(G264), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n538), .A2(new_n396), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n538), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n541), .A2(new_n398), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n522), .A2(new_n528), .A3(new_n540), .A4(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(G270), .B(new_n250), .C1(new_n468), .C2(new_n469), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT82), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n545), .A2(new_n546), .A3(new_n467), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n546), .B1(new_n545), .B2(new_n467), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n212), .A2(G1698), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n399), .B(new_n550), .C1(G257), .C2(G1698), .ZN(new_n551));
  XNOR2_X1  g0351(.A(KEYINPUT83), .B(G303), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n259), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n250), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n549), .A2(new_n554), .A3(new_n414), .ZN(new_n555));
  INV_X1    g0355(.A(G116), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n283), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n451), .B(new_n230), .C1(G33), .C2(new_n205), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n558), .B(new_n281), .C1(new_n230), .C2(G116), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT20), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n559), .A2(new_n560), .ZN(new_n562));
  OAI221_X1 g0362(.A(new_n557), .B1(new_n556), .B2(new_n489), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n555), .A2(new_n563), .ZN(new_n564));
  OR2_X1    g0364(.A1(new_n547), .A2(new_n548), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n551), .A2(new_n553), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n251), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(G169), .A3(new_n563), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT21), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n568), .A2(G200), .ZN(new_n572));
  INV_X1    g0372(.A(new_n563), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n565), .A2(new_n567), .A3(G190), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n568), .A2(KEYINPUT21), .A3(G169), .A4(new_n563), .ZN(new_n576));
  AND4_X1   g0376(.A1(new_n564), .A2(new_n571), .A3(new_n575), .A4(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(G238), .A2(G1698), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n578), .B1(new_n211), .B2(G1698), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n579), .B(new_n256), .C1(new_n255), .C2(new_n361), .ZN(new_n580));
  NAND2_X1  g0380(.A1(G33), .A2(G116), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n250), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n250), .A2(new_n459), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n460), .B1(new_n584), .B2(G250), .ZN(new_n585));
  AOI21_X1  g0385(.A(G169), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n585), .ZN(new_n587));
  NOR3_X1   g0387(.A1(new_n582), .A2(new_n587), .A3(G179), .ZN(new_n588));
  OAI21_X1  g0388(.A(KEYINPUT81), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n583), .A2(new_n414), .A3(new_n585), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT81), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n582), .A2(new_n587), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n590), .B(new_n591), .C1(new_n592), .C2(G169), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT19), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n230), .B1(new_n292), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(G87), .B2(new_n207), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n594), .B1(new_n277), .B2(new_n205), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n230), .A2(G68), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n596), .B(new_n597), .C1(new_n362), .C2(new_n598), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n599), .A2(new_n281), .B1(new_n283), .B2(new_n278), .ZN(new_n600));
  OR2_X1    g0400(.A1(new_n489), .A2(new_n278), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n589), .A2(new_n593), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n490), .A2(G87), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n592), .A2(G190), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n605), .B(new_n606), .C1(new_n398), .C2(new_n592), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n520), .A2(new_n521), .A3(new_n528), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n538), .A2(G179), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(new_n288), .B2(new_n538), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n608), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n503), .A2(new_n544), .A3(new_n577), .A4(new_n612), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n345), .A2(new_n446), .A3(new_n613), .ZN(G372));
  INV_X1    g0414(.A(KEYINPUT89), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n327), .A2(new_n340), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n290), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n405), .A2(new_n411), .ZN(new_n618));
  INV_X1    g0418(.A(new_n408), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n409), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n344), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n617), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n413), .A2(new_n418), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n420), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n413), .A2(KEYINPUT18), .A3(new_n418), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n615), .B1(new_n624), .B2(new_n628), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n615), .B(new_n628), .C1(new_n341), .C2(new_n622), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n439), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n441), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT90), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(KEYINPUT90), .B(new_n441), .C1(new_n629), .C2(new_n631), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n446), .A2(new_n345), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT87), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n582), .A2(new_n638), .ZN(new_n639));
  AOI211_X1 g0439(.A(KEYINPUT87), .B(new_n250), .C1(new_n580), .C2(new_n581), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n585), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n588), .B1(new_n641), .B2(new_n288), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT88), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI211_X1 g0444(.A(KEYINPUT88), .B(new_n588), .C1(new_n641), .C2(new_n288), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n602), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n497), .ZN(new_n647));
  AOI21_X1  g0447(.A(KEYINPUT77), .B1(new_n496), .B2(new_n491), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n641), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n606), .B(new_n605), .C1(new_n650), .C2(new_n398), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n646), .A2(new_n502), .A3(new_n649), .A4(new_n651), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n652), .A2(KEYINPUT26), .ZN(new_n653));
  INV_X1    g0453(.A(new_n651), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n609), .A2(new_n611), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n571), .A2(new_n564), .A3(new_n576), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n657), .A2(new_n503), .A3(new_n544), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n502), .A2(new_n493), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT26), .B1(new_n659), .B2(new_n608), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n653), .A2(new_n658), .A3(new_n646), .A4(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n637), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n636), .A2(new_n662), .ZN(G369));
  NOR2_X1   g0463(.A1(new_n282), .A2(G20), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n262), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G213), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(G343), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n563), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n577), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n656), .B2(new_n671), .ZN(new_n673));
  XNOR2_X1  g0473(.A(KEYINPUT91), .B(G330), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n655), .ZN(new_n677));
  INV_X1    g0477(.A(new_n670), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR3_X1   g0479(.A1(new_n609), .A2(new_n539), .A3(new_n542), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n680), .B1(new_n609), .B2(new_n670), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n679), .B1(new_n681), .B2(new_n677), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n656), .A2(new_n670), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n676), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n656), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n681), .A2(new_n686), .A3(new_n655), .A4(new_n678), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n687), .A2(new_n679), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n685), .A2(new_n688), .ZN(G399));
  INV_X1    g0489(.A(new_n226), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G41), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G1), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n393), .A2(new_n205), .A3(new_n206), .A4(new_n556), .ZN(new_n694));
  OAI22_X1  g0494(.A1(new_n693), .A2(new_n694), .B1(new_n229), .B2(new_n692), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT28), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n661), .A2(new_n678), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT29), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n659), .A2(new_n608), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT26), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n652), .A2(KEYINPUT26), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n658), .A2(new_n646), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n704), .A2(KEYINPUT29), .A3(new_n678), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n536), .A2(new_n537), .A3(new_n592), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n477), .A2(new_n555), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n555), .A2(new_n477), .A3(new_n706), .A4(KEYINPUT30), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n473), .A2(new_n414), .A3(new_n568), .A4(new_n641), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n709), .B(new_n710), .C1(new_n711), .C2(new_n541), .ZN(new_n712));
  XNOR2_X1  g0512(.A(KEYINPUT92), .B(KEYINPUT31), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(new_n670), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(new_n670), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n714), .B(new_n717), .C1(new_n613), .C2(new_n670), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n699), .A2(new_n705), .B1(new_n674), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n696), .B1(new_n719), .B2(G1), .ZN(G364));
  NOR2_X1   g0520(.A1(new_n230), .A2(new_n414), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n721), .A2(KEYINPUT95), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n396), .A2(G200), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n721), .A2(KEYINPUT95), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n721), .A2(G200), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n396), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n726), .A2(G58), .B1(G50), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(G190), .A2(G200), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n722), .A2(new_n730), .A3(new_n724), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n732), .A2(KEYINPUT96), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(KEYINPUT96), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n729), .B1(new_n736), .B2(new_n210), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT97), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n230), .A2(G179), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n739), .A2(G190), .A3(G200), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G87), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n739), .A2(new_n730), .ZN(new_n743));
  INV_X1    g0543(.A(G159), .ZN(new_n744));
  OAI21_X1  g0544(.A(KEYINPUT32), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n739), .A2(new_n396), .A3(G200), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n206), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n743), .A2(KEYINPUT32), .A3(new_n744), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n746), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n727), .A2(G190), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n259), .B1(new_n751), .B2(G68), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n230), .B1(new_n723), .B2(new_n414), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G97), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n738), .A2(new_n750), .A3(new_n752), .A4(new_n755), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT98), .Z(new_n757));
  INV_X1    g0557(.A(new_n728), .ZN(new_n758));
  INV_X1    g0558(.A(G326), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI22_X1  g0560(.A1(G322), .A2(new_n726), .B1(new_n732), .B2(G311), .ZN(new_n761));
  INV_X1    g0561(.A(new_n743), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G329), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n761), .A2(new_n259), .A3(new_n763), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n760), .B(new_n764), .C1(G294), .C2(new_n754), .ZN(new_n765));
  INV_X1    g0565(.A(G317), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(KEYINPUT33), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n766), .A2(KEYINPUT33), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n751), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n747), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G283), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n741), .A2(G303), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n765), .A2(new_n769), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n757), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n231), .B1(G20), .B2(new_n288), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G13), .A2(G33), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n776), .B(KEYINPUT94), .Z(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n775), .ZN(new_n780));
  OAI21_X1  g0580(.A(KEYINPUT72), .B1(new_n357), .B2(new_n358), .ZN(new_n781));
  OAI211_X1 g0581(.A(new_n349), .B(new_n256), .C1(new_n361), .C2(new_n255), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n690), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(G45), .B2(new_n244), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(G45), .B2(new_n229), .ZN(new_n788));
  NAND3_X1  g0588(.A1(G355), .A2(new_n252), .A3(new_n226), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(G116), .B2(new_n226), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT93), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n774), .A2(new_n775), .B1(new_n780), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n693), .B1(G45), .B2(new_n664), .ZN(new_n794));
  INV_X1    g0594(.A(new_n779), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n793), .B(new_n794), .C1(new_n673), .C2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n676), .A2(new_n794), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(new_n674), .B2(new_n673), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(G396));
  AND2_X1   g0600(.A1(new_n287), .A2(new_n670), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n290), .B1(new_n444), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n291), .A2(new_n678), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n697), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n804), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n661), .A2(new_n678), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n718), .A2(new_n674), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n808), .B(new_n809), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n810), .A2(new_n794), .ZN(new_n811));
  INV_X1    g0611(.A(G132), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n784), .B1(new_n812), .B2(new_n743), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n735), .A2(G159), .B1(G143), .B2(new_n726), .ZN(new_n814));
  INV_X1    g0614(.A(G137), .ZN(new_n815));
  INV_X1    g0615(.A(new_n751), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n814), .B1(new_n815), .B2(new_n758), .C1(new_n425), .C2(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT34), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n818), .B1(new_n218), .B2(new_n753), .C1(new_n221), .C2(new_n747), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n813), .B(new_n819), .C1(G50), .C2(new_n741), .ZN(new_n820));
  INV_X1    g0620(.A(G311), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n725), .A2(new_n529), .B1(new_n821), .B2(new_n743), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n735), .A2(G116), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n770), .A2(G87), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n751), .A2(G283), .B1(new_n728), .B2(G303), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n252), .B1(new_n754), .B2(G97), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n823), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n822), .B(new_n827), .C1(G107), .C2(new_n741), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n775), .B1(new_n820), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n775), .A2(new_n776), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n804), .A2(new_n777), .B1(new_n210), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n829), .A2(new_n794), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n811), .A2(new_n832), .ZN(G384));
  NAND3_X1  g0633(.A1(new_n712), .A2(KEYINPUT31), .A3(new_n670), .ZN(new_n834));
  INV_X1    g0634(.A(new_n713), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n715), .A2(new_n835), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n834), .B(new_n836), .C1(new_n613), .C2(new_n670), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n637), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT103), .ZN(new_n839));
  AND3_X1   g0639(.A1(new_n327), .A2(new_n340), .A3(new_n678), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n340), .A2(new_n670), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n327), .A2(new_n340), .B1(new_n344), .B2(new_n841), .ZN(new_n842));
  NOR3_X1   g0642(.A1(new_n840), .A2(new_n842), .A3(new_n804), .ZN(new_n843));
  OR2_X1    g0643(.A1(new_n369), .A2(new_n370), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n347), .B1(new_n781), .B2(new_n782), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n845), .A2(new_n363), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n844), .B1(new_n846), .B2(G68), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n428), .B1(new_n847), .B2(KEYINPUT16), .ZN(new_n848));
  NOR3_X1   g0648(.A1(new_n845), .A2(new_n221), .A3(new_n363), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n378), .B1(new_n849), .B2(new_n844), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n382), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n851), .A2(new_n668), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n422), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n405), .B1(new_n851), .B2(new_n417), .ZN(new_n854));
  OAI21_X1  g0654(.A(KEYINPUT37), .B1(new_n854), .B2(new_n852), .ZN(new_n855));
  INV_X1    g0655(.A(new_n668), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n413), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT37), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n625), .A2(new_n857), .A3(new_n858), .A4(new_n405), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n853), .A2(new_n860), .A3(KEYINPUT38), .ZN(new_n861));
  XNOR2_X1  g0661(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n857), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n422), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n625), .A2(new_n857), .A3(new_n405), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(KEYINPUT37), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n859), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n863), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n843), .B(new_n837), .C1(new_n861), .C2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n840), .A2(new_n842), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n837), .A2(new_n871), .A3(new_n806), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n380), .A2(new_n383), .A3(new_n404), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n850), .A2(new_n281), .A3(new_n372), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n417), .B1(new_n875), .B2(new_n383), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(new_n383), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n856), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n858), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n859), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n879), .B1(new_n621), .B2(new_n628), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n873), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n853), .A2(new_n860), .A3(KEYINPUT38), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT40), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n870), .A2(KEYINPUT40), .B1(new_n872), .B2(new_n886), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n839), .B(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n674), .ZN(new_n889));
  INV_X1    g0689(.A(new_n646), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n475), .A2(G200), .A3(new_n478), .ZN(new_n891));
  OAI22_X1  g0691(.A1(new_n647), .A2(new_n648), .B1(new_n396), .B2(new_n473), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n659), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n893), .A2(new_n680), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n890), .B1(new_n894), .B2(new_n657), .ZN(new_n895));
  MUX2_X1   g0695(.A(new_n700), .B(new_n652), .S(new_n701), .Z(new_n896));
  AOI21_X1  g0696(.A(new_n670), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n637), .B(new_n705), .C1(new_n897), .C2(KEYINPUT29), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT101), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT101), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n699), .A2(new_n900), .A3(new_n637), .A4(new_n705), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n636), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n889), .B(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n840), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n861), .A2(new_n869), .A3(KEYINPUT39), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT39), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n884), .B2(new_n885), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT100), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n869), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(new_n907), .A3(new_n885), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT38), .B1(new_n853), .B2(new_n860), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT39), .B1(new_n861), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT100), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n911), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n905), .B1(new_n909), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n628), .A2(new_n856), .ZN(new_n918));
  INV_X1    g0718(.A(new_n871), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(new_n807), .B2(new_n803), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n861), .A2(new_n912), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n918), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n917), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT102), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n904), .B(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n262), .B2(new_n664), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n483), .A2(new_n485), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT35), .ZN(new_n929));
  AOI211_X1 g0729(.A(new_n230), .B(new_n231), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n930), .B(G116), .C1(new_n929), .C2(new_n928), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT36), .ZN(new_n932));
  OAI21_X1  g0732(.A(G77), .B1(new_n218), .B2(new_n221), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n933), .A2(new_n229), .B1(G50), .B2(new_n221), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(G1), .A3(new_n282), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n927), .A2(new_n932), .A3(new_n935), .ZN(G367));
  AOI22_X1  g0736(.A1(new_n735), .A2(G50), .B1(G137), .B2(new_n762), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n770), .A2(G77), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n728), .A2(G143), .B1(new_n754), .B2(G68), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n425), .B2(new_n725), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(KEYINPUT107), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n252), .B1(new_n940), .B2(KEYINPUT107), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n816), .A2(new_n744), .B1(new_n218), .B2(new_n740), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n937), .A2(new_n938), .A3(new_n941), .A4(new_n944), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n816), .A2(new_n529), .B1(new_n205), .B2(new_n747), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n735), .B2(G283), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT46), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n741), .A2(G116), .ZN(new_n949));
  OAI221_X1 g0749(.A(new_n947), .B1(new_n948), .B2(new_n949), .C1(new_n821), .C2(new_n758), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n948), .B2(new_n949), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n726), .A2(new_n552), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n784), .B1(G107), .B2(new_n754), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(KEYINPUT106), .B(G317), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n762), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n945), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT47), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n775), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n780), .B1(new_n226), .B2(new_n278), .C1(new_n786), .C2(new_n240), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n959), .A2(new_n794), .A3(new_n960), .ZN(new_n961));
  OR3_X1    g0761(.A1(new_n646), .A2(new_n605), .A3(new_n678), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n646), .B(new_n651), .C1(new_n605), .C2(new_n678), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n964), .A2(new_n795), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n685), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n649), .A2(new_n670), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n503), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n649), .A2(new_n502), .A3(new_n670), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n967), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT104), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n973), .B(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n687), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n971), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT42), .Z(new_n978));
  AOI21_X1  g0778(.A(new_n655), .B1(new_n969), .B2(new_n970), .ZN(new_n979));
  INV_X1    g0779(.A(new_n659), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n678), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n978), .A2(new_n981), .B1(KEYINPUT43), .B2(new_n964), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n975), .B(new_n982), .Z(new_n983));
  AOI21_X1  g0783(.A(new_n262), .B1(new_n664), .B2(G45), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT45), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n688), .A2(new_n971), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT105), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n986), .A2(KEYINPUT105), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n985), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n989), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n991), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n688), .A2(new_n971), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT44), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n990), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  NOR3_X1   g0795(.A1(new_n683), .A2(new_n676), .A3(new_n684), .ZN(new_n996));
  NOR3_X1   g0796(.A1(new_n967), .A2(new_n996), .A3(new_n976), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n719), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n995), .A2(new_n999), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n1000), .A2(new_n719), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n691), .B(KEYINPUT41), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n984), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n966), .B1(new_n983), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(G387));
  INV_X1    g0806(.A(new_n984), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n997), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n691), .B1(new_n997), .B2(new_n719), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n753), .A2(new_n278), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n726), .A2(G50), .B1(G97), .B2(new_n770), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n221), .B2(new_n731), .C1(new_n210), .C2(new_n740), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1010), .B(new_n1012), .C1(new_n274), .C2(new_n751), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n783), .B1(G150), .B2(new_n762), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(new_n744), .C2(new_n758), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n735), .A2(new_n552), .B1(new_n726), .B2(new_n955), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT109), .Z(new_n1017));
  AOI22_X1  g0817(.A1(new_n751), .A2(G311), .B1(new_n728), .B2(G322), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT110), .Z(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT48), .ZN(new_n1021));
  INV_X1    g0821(.A(G283), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1021), .B1(new_n1022), .B2(new_n753), .C1(new_n529), .C2(new_n740), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT49), .Z(new_n1024));
  OAI221_X1 g0824(.A(new_n783), .B1(new_n556), .B2(new_n747), .C1(new_n759), .C2(new_n743), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1015), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT111), .Z(new_n1027));
  AND2_X1   g0827(.A1(new_n1027), .A2(new_n775), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n274), .A2(new_n202), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1029), .A2(KEYINPUT50), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n694), .B1(new_n1029), .B2(KEYINPUT50), .ZN(new_n1031));
  INV_X1    g0831(.A(G45), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(G68), .A2(G77), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n785), .B(new_n1034), .C1(new_n237), .C2(new_n1032), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n252), .A2(new_n694), .A3(new_n226), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(G107), .B2(new_n226), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT108), .Z(new_n1038));
  NAND2_X1  g0838(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n780), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n794), .B(new_n1040), .C1(new_n683), .C2(new_n795), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1008), .B1(new_n999), .B2(new_n1009), .C1(new_n1028), .C2(new_n1041), .ZN(G393));
  AOI22_X1  g0842(.A1(new_n735), .A2(new_n274), .B1(G50), .B2(new_n751), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT112), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1044), .B(new_n824), .C1(new_n221), .C2(new_n740), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n754), .A2(G77), .B1(new_n762), .B2(G143), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n784), .A2(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n726), .A2(G159), .B1(G150), .B2(new_n728), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT51), .ZN(new_n1049));
  NOR3_X1   g0849(.A1(new_n1045), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n821), .A2(new_n725), .B1(new_n758), .B2(new_n766), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT52), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n732), .A2(G294), .B1(G116), .B2(new_n754), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n259), .B1(new_n740), .B2(new_n1022), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n748), .B(new_n1054), .C1(G322), .C2(new_n762), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1052), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n552), .B2(new_n751), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n775), .B1(new_n1050), .B2(new_n1057), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n780), .B1(new_n205), .B2(new_n226), .C1(new_n786), .C2(new_n247), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n969), .A2(new_n779), .A3(new_n970), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1058), .A2(new_n794), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1000), .A2(KEYINPUT113), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n995), .A2(new_n967), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n990), .A2(new_n992), .A3(new_n685), .A4(new_n994), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n999), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n692), .B1(new_n1066), .B2(KEYINPUT113), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1062), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT114), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1064), .A2(new_n1007), .A3(new_n1065), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1070), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(G390));
  NAND3_X1  g0875(.A1(new_n837), .A2(G330), .A3(new_n806), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n919), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n704), .A2(new_n678), .A3(new_n802), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n718), .A2(new_n871), .A3(new_n674), .A4(new_n806), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1077), .A2(new_n803), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n718), .A2(new_n674), .A3(new_n806), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n872), .A2(G330), .B1(new_n1081), .B2(new_n919), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n807), .A2(new_n803), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1080), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n838), .A2(G330), .ZN(new_n1086));
  AND4_X1   g0886(.A1(new_n636), .A2(new_n1085), .A3(new_n902), .A4(new_n1086), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n909), .B(new_n915), .C1(new_n840), .C2(new_n920), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1079), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n865), .A2(new_n868), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n422), .A2(new_n852), .B1(new_n855), .B2(new_n859), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1090), .A2(new_n862), .B1(new_n1091), .B2(KEYINPUT38), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1092), .A2(new_n840), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1078), .A2(new_n803), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1093), .B1(new_n1094), .B2(new_n919), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1088), .A2(new_n1089), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1088), .A2(new_n1095), .B1(G330), .B2(new_n872), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1087), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n909), .A2(new_n915), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n920), .A2(new_n840), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1095), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n872), .A2(G330), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1085), .A2(new_n902), .A3(new_n636), .A4(new_n1086), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1104), .A2(new_n1105), .A3(new_n1096), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1099), .A2(new_n691), .A3(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n909), .A2(new_n777), .A3(new_n915), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n259), .B(new_n742), .C1(new_n725), .C2(new_n556), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n751), .A2(G107), .B1(new_n728), .B2(G283), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n736), .B2(new_n205), .ZN(new_n1111));
  XOR2_X1   g0911(.A(new_n1111), .B(KEYINPUT117), .Z(new_n1112));
  OAI221_X1 g0912(.A(new_n1112), .B1(new_n221), .B2(new_n747), .C1(new_n529), .C2(new_n743), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n1109), .B(new_n1113), .C1(G77), .C2(new_n754), .ZN(new_n1114));
  XOR2_X1   g0914(.A(KEYINPUT54), .B(G143), .Z(new_n1115));
  NAND2_X1  g0915(.A1(new_n735), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n741), .A2(G150), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT116), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(KEYINPUT53), .ZN(new_n1119));
  OR2_X1    g0919(.A1(new_n1118), .A2(KEYINPUT53), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n725), .A2(new_n812), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n252), .B1(new_n816), .B2(new_n815), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n1121), .B(new_n1122), .C1(G128), .C2(new_n728), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1116), .A2(new_n1119), .A3(new_n1120), .A4(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n747), .A2(new_n202), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n753), .A2(new_n744), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n762), .A2(G125), .ZN(new_n1127));
  NOR4_X1   g0927(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n775), .B1(new_n1114), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n830), .A2(new_n273), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1108), .A2(new_n794), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1104), .A2(new_n1096), .ZN(new_n1132));
  AOI21_X1  g0932(.A(KEYINPUT115), .B1(new_n1132), .B2(new_n1007), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT115), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1134), .B(new_n984), .C1(new_n1104), .C2(new_n1096), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1107), .B(new_n1131), .C1(new_n1133), .C2(new_n1135), .ZN(G378));
  OAI22_X1  g0936(.A1(new_n731), .A2(new_n278), .B1(new_n221), .B2(new_n753), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n784), .A2(G41), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n747), .A2(new_n218), .B1(new_n743), .B2(new_n1022), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(G77), .B2(new_n741), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  XOR2_X1   g0941(.A(new_n1141), .B(KEYINPUT118), .Z(new_n1142));
  AOI211_X1 g0942(.A(new_n1137), .B(new_n1142), .C1(G116), .C2(new_n728), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1143), .B1(new_n205), .B2(new_n816), .C1(new_n206), .C2(new_n725), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT58), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n255), .A2(new_n465), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n726), .A2(G128), .B1(new_n741), .B2(new_n1115), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n751), .A2(G132), .B1(new_n754), .B2(G150), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1147), .B(new_n1148), .C1(new_n815), .C2(new_n731), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G125), .B2(new_n728), .ZN(new_n1150));
  XOR2_X1   g0950(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n1151));
  XNOR2_X1  g0951(.A(new_n1150), .B(new_n1151), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1146), .B(new_n1152), .C1(G124), .C2(new_n762), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n770), .A2(G159), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1138), .A2(G50), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n1153), .A2(new_n1154), .B1(new_n1146), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1145), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n775), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n429), .A2(new_n856), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n439), .A2(new_n441), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1161), .B1(new_n439), .B2(new_n441), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1160), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1164), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1166), .A2(new_n1162), .A3(new_n1159), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n777), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n830), .A2(new_n202), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1158), .A2(new_n1170), .A3(new_n794), .A4(new_n1171), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n1172), .B(KEYINPUT120), .Z(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n843), .A2(new_n837), .ZN(new_n1175));
  OAI21_X1  g0975(.A(KEYINPUT40), .B1(new_n1175), .B2(new_n1092), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n872), .A2(new_n886), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1169), .B1(new_n1178), .B2(G330), .ZN(new_n1179));
  INV_X1    g0979(.A(G330), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1180), .B(new_n1168), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n917), .B(new_n923), .C1(new_n1179), .C2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1168), .B1(new_n887), .B2(new_n1180), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1178), .A2(G330), .A3(new_n1169), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1083), .A2(new_n871), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n1185), .A2(new_n921), .B1(new_n628), .B2(new_n856), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1183), .B(new_n1184), .C1(new_n1186), .C2(new_n916), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1182), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1174), .B1(new_n1007), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n902), .A2(new_n636), .A3(new_n1086), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1099), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(KEYINPUT57), .B1(new_n1193), .B2(new_n1188), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1105), .B1(new_n1104), .B2(new_n1096), .ZN(new_n1195));
  OAI21_X1  g0995(.A(KEYINPUT57), .B1(new_n1195), .B2(new_n1191), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1182), .A2(KEYINPUT121), .A3(new_n1187), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT121), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n924), .A2(new_n1198), .A3(new_n1184), .A4(new_n1183), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n691), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1194), .B1(new_n1201), .B2(KEYINPUT122), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT122), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1203), .B(new_n691), .C1(new_n1196), .C2(new_n1200), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1190), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(G375));
  INV_X1    g1006(.A(new_n1085), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1191), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1208), .A2(new_n1002), .A3(new_n1105), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n919), .A2(new_n776), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n735), .A2(G107), .B1(G116), .B2(new_n751), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n205), .B2(new_n740), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n762), .A2(G303), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n938), .A2(new_n259), .ZN(new_n1214));
  XOR2_X1   g1014(.A(new_n1214), .B(KEYINPUT123), .Z(new_n1215));
  AOI21_X1  g1015(.A(new_n1010), .B1(G294), .B2(new_n728), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n1022), .B2(new_n725), .ZN(new_n1217));
  NOR4_X1   g1017(.A1(new_n1212), .A2(new_n1213), .A3(new_n1215), .A4(new_n1217), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n732), .A2(G150), .B1(G128), .B2(new_n762), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1219), .B1(new_n218), .B2(new_n747), .C1(new_n744), .C2(new_n740), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n784), .B1(new_n815), .B2(new_n725), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n751), .A2(new_n1115), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n758), .A2(new_n812), .B1(new_n202), .B2(new_n753), .ZN(new_n1223));
  NOR4_X1   g1023(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n775), .B1(new_n1218), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n830), .A2(new_n221), .ZN(new_n1226));
  AND4_X1   g1026(.A1(new_n794), .A2(new_n1210), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n1085), .B2(new_n1007), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1209), .A2(new_n1228), .ZN(G381));
  NAND2_X1  g1029(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1230), .A2(new_n1071), .A3(new_n1061), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(KEYINPUT114), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1232), .A2(new_n1005), .A3(new_n1233), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(new_n1234), .A2(G396), .A3(G393), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(G375), .A2(G378), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(G381), .A2(G384), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .ZN(G407));
  INV_X1    g1038(.A(G213), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(new_n1236), .B2(new_n669), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(G407), .A2(new_n1240), .ZN(G409));
  INV_X1    g1041(.A(KEYINPUT60), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n691), .B(new_n1105), .C1(new_n1208), .C2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT60), .B1(new_n1191), .B2(new_n1207), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1228), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1245), .A2(new_n811), .A3(new_n832), .ZN(new_n1246));
  OAI211_X1 g1046(.A(G384), .B(new_n1228), .C1(new_n1243), .C2(new_n1244), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1239), .A2(G343), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1107), .A2(new_n1131), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n1253), .B(new_n1190), .C1(new_n1202), .C2(new_n1204), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1002), .B(new_n1188), .C1(new_n1195), .C2(new_n1191), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1197), .A2(new_n1007), .A3(new_n1199), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1255), .A2(new_n1172), .A3(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(KEYINPUT124), .B1(new_n1257), .B2(G378), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT124), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1255), .A2(new_n1172), .A3(new_n1256), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1253), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1248), .B(new_n1250), .C1(new_n1254), .C2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(KEYINPUT62), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1249), .A2(KEYINPUT125), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1248), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1249), .A2(G2897), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1248), .A2(G2897), .A3(new_n1249), .A4(new_n1265), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1262), .B1(G378), .B2(new_n1205), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1270), .B1(new_n1271), .B2(new_n1249), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT61), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1194), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT57), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(new_n1099), .B2(new_n1192), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n692), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1275), .B1(new_n1279), .B2(new_n1203), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1204), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G378), .B(new_n1189), .C1(new_n1280), .C2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1274), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT62), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1283), .A2(new_n1284), .A3(new_n1248), .A4(new_n1250), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1264), .A2(new_n1272), .A3(new_n1273), .A4(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(KEYINPUT127), .ZN(new_n1287));
  OAI21_X1  g1087(.A(G387), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT126), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1288), .A2(new_n1234), .A3(new_n1289), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(G393), .B(G396), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1291), .A2(new_n1288), .A3(new_n1289), .A4(new_n1234), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1283), .A2(new_n1250), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT61), .B1(new_n1296), .B2(new_n1270), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT127), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1297), .A2(new_n1298), .A3(new_n1285), .A4(new_n1264), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1287), .A2(new_n1295), .A3(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1272), .A2(KEYINPUT63), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT61), .B1(new_n1301), .B2(new_n1263), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1283), .A2(KEYINPUT63), .A3(new_n1248), .A4(new_n1250), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1302), .A2(new_n1303), .A3(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1300), .A2(new_n1305), .ZN(G405));
  XNOR2_X1  g1106(.A(new_n1205), .B(G378), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(new_n1307), .B(new_n1248), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(new_n1308), .B(new_n1295), .ZN(G402));
endmodule


