//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 1 0 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n572, new_n574, new_n575,
    new_n576, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n609, new_n611, new_n612,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1141, new_n1142,
    new_n1144;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT66), .B(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT67), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT68), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT69), .Z(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G236), .A3(G235), .A4(G238), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT70), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(new_n454), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G137), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G101), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT71), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI211_X1 g046(.A(KEYINPUT71), .B(G125), .C1(new_n464), .C2(new_n465), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n468), .B1(new_n474), .B2(G2105), .ZN(G160));
  NOR2_X1   g050(.A1(new_n464), .A2(new_n465), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT72), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  INV_X1    g054(.A(G2105), .ZN(new_n480));
  OAI21_X1  g055(.A(KEYINPUT73), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  OR2_X1    g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT73), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n484), .A2(new_n485), .A3(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT74), .B1(G100), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NOR3_X1   g065(.A1(KEYINPUT74), .A2(G100), .A3(G2105), .ZN(new_n491));
  OAI221_X1 g066(.A(G2104), .B1(G112), .B2(new_n480), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n479), .A2(new_n488), .A3(new_n492), .ZN(new_n493));
  XOR2_X1   g068(.A(new_n493), .B(KEYINPUT75), .Z(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  NAND2_X1  g070(.A1(G126), .A2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G2104), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(G102), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(new_n480), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n484), .A2(new_n497), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  OAI211_X1 g078(.A(G138), .B(new_n480), .C1(new_n464), .C2(new_n465), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n484), .A2(KEYINPUT4), .A3(G138), .A4(new_n480), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n503), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT76), .B1(new_n510), .B2(KEYINPUT6), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT76), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(new_n513), .A3(G651), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n511), .A2(new_n514), .B1(KEYINPUT6), .B2(new_n510), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  OAI21_X1  g091(.A(KEYINPUT77), .B1(new_n516), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT77), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n518), .A2(new_n519), .A3(KEYINPUT5), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n517), .A2(new_n520), .B1(new_n516), .B2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n515), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G50), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n522), .A2(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n510), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n526), .A2(new_n528), .ZN(G166));
  AND2_X1   g104(.A1(new_n515), .A2(new_n521), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT7), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n530), .A2(G89), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  XNOR2_X1  g108(.A(KEYINPUT78), .B(G51), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n524), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n521), .A2(G63), .ZN(new_n536));
  NAND3_X1  g111(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n510), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n535), .A2(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  INV_X1    g116(.A(G52), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n522), .A2(new_n541), .B1(new_n524), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n510), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n543), .A2(new_n545), .ZN(G171));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  INV_X1    g122(.A(G43), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n522), .A2(new_n547), .B1(new_n524), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n510), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(new_n521), .A2(G65), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n560), .A2(G651), .B1(new_n530), .B2(G91), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  AND2_X1   g137(.A1(KEYINPUT79), .A2(G53), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n515), .A2(G543), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(KEYINPUT9), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n515), .A2(new_n566), .A3(G543), .A4(new_n563), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n562), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(G299));
  XNOR2_X1  g146(.A(G171), .B(KEYINPUT80), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G301));
  INV_X1    g148(.A(KEYINPUT81), .ZN(new_n574));
  NAND2_X1  g149(.A1(G166), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT81), .B1(new_n526), .B2(new_n528), .ZN(new_n576));
  AND2_X1   g151(.A1(new_n575), .A2(new_n576), .ZN(G303));
  OAI21_X1  g152(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n578));
  INV_X1    g153(.A(G49), .ZN(new_n579));
  INV_X1    g154(.A(G87), .ZN(new_n580));
  OAI221_X1 g155(.A(new_n578), .B1(new_n524), .B2(new_n579), .C1(new_n580), .C2(new_n522), .ZN(new_n581));
  XOR2_X1   g156(.A(new_n581), .B(KEYINPUT82), .Z(G288));
  INV_X1    g157(.A(G86), .ZN(new_n583));
  INV_X1    g158(.A(G48), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n522), .A2(new_n583), .B1(new_n524), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n521), .A2(G61), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT83), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n510), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G305));
  INV_X1    g166(.A(new_n524), .ZN(new_n592));
  AOI22_X1  g167(.A1(G47), .A2(new_n592), .B1(new_n530), .B2(G85), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n510), .B2(new_n594), .ZN(G290));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NOR2_X1   g171(.A1(G301), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n592), .A2(G54), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n521), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n599));
  AND3_X1   g174(.A1(new_n530), .A2(KEYINPUT10), .A3(G92), .ZN(new_n600));
  AOI21_X1  g175(.A(KEYINPUT10), .B1(new_n530), .B2(G92), .ZN(new_n601));
  OAI221_X1 g176(.A(new_n598), .B1(new_n510), .B2(new_n599), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  XOR2_X1   g177(.A(new_n602), .B(KEYINPUT84), .Z(new_n603));
  AOI21_X1  g178(.A(new_n597), .B1(new_n603), .B2(new_n596), .ZN(G284));
  AOI21_X1  g179(.A(new_n597), .B1(new_n603), .B2(new_n596), .ZN(G321));
  NAND2_X1  g180(.A1(G286), .A2(G868), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G868), .B2(new_n570), .ZN(G297));
  OAI21_X1  g182(.A(new_n606), .B1(G868), .B2(new_n570), .ZN(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n603), .B1(new_n609), .B2(G860), .ZN(G148));
  NAND2_X1  g185(.A1(new_n603), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT85), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n487), .A2(G123), .ZN(new_n616));
  OR2_X1    g191(.A1(G99), .A2(G2105), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n617), .B(G2104), .C1(G111), .C2(new_n480), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(G135), .B2(new_n478), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT86), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n621), .A2(G2096), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(G2096), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n477), .A2(G2104), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2100), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n622), .A2(new_n623), .A3(new_n627), .ZN(G156));
  XOR2_X1   g203(.A(G2451), .B(G2454), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT16), .ZN(new_n630));
  XNOR2_X1  g205(.A(G1341), .B(G1348), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(new_n639), .A3(KEYINPUT14), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n634), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n634), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(new_n643), .A3(G14), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT87), .ZN(G401));
  INV_X1    g220(.A(KEYINPUT18), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2084), .B(G2090), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT88), .ZN(new_n648));
  XOR2_X1   g223(.A(G2067), .B(G2678), .Z(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(KEYINPUT17), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n648), .A2(new_n649), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n646), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2072), .B(G2078), .Z(new_n654));
  NOR2_X1   g229(.A1(new_n652), .A2(new_n646), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n656), .B1(new_n653), .B2(new_n654), .ZN(new_n657));
  XOR2_X1   g232(.A(G2096), .B(G2100), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT89), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(new_n659), .ZN(G227));
  XOR2_X1   g235(.A(G1971), .B(G1976), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1956), .B(G2474), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1961), .B(G1966), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n662), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n662), .A2(new_n665), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT20), .Z(new_n669));
  AOI211_X1 g244(.A(new_n667), .B(new_n669), .C1(new_n662), .C2(new_n666), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G1986), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1991), .B(G1996), .ZN(new_n674));
  INV_X1    g249(.A(G1981), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(new_n676), .ZN(G229));
  NAND3_X1  g252(.A1(new_n480), .A2(G103), .A3(G2104), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT25), .Z(new_n679));
  AOI22_X1  g254(.A1(new_n484), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n679), .B1(new_n680), .B2(new_n480), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n478), .B2(G139), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT99), .ZN(new_n683));
  MUX2_X1   g258(.A(G33), .B(new_n683), .S(G29), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT100), .ZN(new_n685));
  INV_X1    g260(.A(G2072), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n686), .ZN(new_n688));
  NAND3_X1  g263(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT26), .ZN(new_n690));
  AND3_X1   g265(.A1(new_n480), .A2(G105), .A3(G2104), .ZN(new_n691));
  AOI211_X1 g266(.A(new_n690), .B(new_n691), .C1(new_n487), .C2(G129), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n478), .A2(G141), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n695), .B2(G32), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT27), .B(G1996), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT24), .ZN(new_n699));
  INV_X1    g274(.A(G34), .ZN(new_n700));
  AOI21_X1  g275(.A(G29), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(new_n699), .B2(new_n700), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G160), .B2(new_n695), .ZN(new_n703));
  AOI22_X1  g278(.A1(new_n697), .A2(new_n698), .B1(G2084), .B2(new_n703), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n687), .A2(new_n688), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT101), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT90), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n707), .A2(G16), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n710), .A2(G19), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(new_n552), .B2(new_n710), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT96), .B(G1341), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n620), .A2(G29), .ZN(new_n715));
  NOR2_X1   g290(.A1(G164), .A2(new_n695), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G27), .B2(new_n695), .ZN(new_n717));
  INV_X1    g292(.A(G2078), .ZN(new_n718));
  AOI22_X1  g293(.A1(new_n715), .A2(KEYINPUT103), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  MUX2_X1   g294(.A(G21), .B(G286), .S(G16), .Z(new_n720));
  OAI221_X1 g295(.A(new_n719), .B1(new_n718), .B2(new_n717), .C1(new_n720), .C2(G1966), .ZN(new_n721));
  AOI211_X1 g296(.A(new_n714), .B(new_n721), .C1(G1966), .C2(new_n720), .ZN(new_n722));
  INV_X1    g297(.A(G4), .ZN(new_n723));
  MUX2_X1   g298(.A(new_n723), .B(new_n603), .S(G16), .Z(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT95), .B(G1348), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT102), .B(KEYINPUT31), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G11), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT30), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n695), .B1(new_n729), .B2(G28), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n729), .B2(G28), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  OAI221_X1 g307(.A(new_n732), .B1(KEYINPUT103), .B2(new_n715), .C1(new_n697), .C2(new_n698), .ZN(new_n733));
  INV_X1    g308(.A(G171), .ZN(new_n734));
  MUX2_X1   g309(.A(G5), .B(new_n734), .S(G16), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1961), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n695), .A2(G26), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT28), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n478), .A2(G140), .ZN(new_n739));
  OR2_X1    g314(.A1(G104), .A2(G2105), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n740), .B(G2104), .C1(G116), .C2(new_n480), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(KEYINPUT97), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(KEYINPUT97), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n487), .A2(G128), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n738), .B1(new_n746), .B2(new_n695), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT98), .B(G2067), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n749), .ZN(new_n751));
  OAI22_X1  g326(.A1(new_n747), .A2(new_n751), .B1(G2084), .B2(new_n703), .ZN(new_n752));
  NOR4_X1   g327(.A1(new_n733), .A2(new_n736), .A3(new_n750), .A4(new_n752), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n722), .A2(new_n726), .A3(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G2090), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n695), .A2(G35), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G162), .B2(new_n695), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT29), .Z(new_n758));
  AOI21_X1  g333(.A(new_n754), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n758), .A2(new_n755), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT104), .B(KEYINPUT23), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT105), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n708), .A2(G20), .A3(new_n709), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G299), .B2(G16), .ZN(new_n765));
  INV_X1    g340(.A(G1956), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(KEYINPUT106), .B1(new_n760), .B2(new_n767), .ZN(new_n768));
  OR3_X1    g343(.A1(new_n760), .A2(KEYINPUT106), .A3(new_n767), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n706), .A2(new_n759), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT36), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n710), .A2(G22), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G166), .B2(new_n710), .ZN(new_n773));
  INV_X1    g348(.A(G1971), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  MUX2_X1   g350(.A(G23), .B(new_n581), .S(G16), .Z(new_n776));
  XOR2_X1   g351(.A(KEYINPUT33), .B(G1976), .Z(new_n777));
  XOR2_X1   g352(.A(new_n776), .B(new_n777), .Z(new_n778));
  MUX2_X1   g353(.A(G6), .B(G305), .S(G16), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT93), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT32), .B(G1981), .Z(new_n781));
  AND2_X1   g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n775), .B(new_n778), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT34), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT94), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n710), .A2(G24), .ZN(new_n788));
  XNOR2_X1  g363(.A(G290), .B(KEYINPUT91), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(new_n710), .ZN(new_n790));
  INV_X1    g365(.A(G1986), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT92), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n792), .A2(new_n793), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n695), .A2(G25), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n478), .A2(G131), .ZN(new_n797));
  OR2_X1    g372(.A1(G95), .A2(G2105), .ZN(new_n798));
  INV_X1    g373(.A(G107), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n498), .B1(new_n799), .B2(G2105), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n487), .A2(G119), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n796), .B1(new_n803), .B2(new_n695), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT35), .B(G1991), .Z(new_n805));
  XOR2_X1   g380(.A(new_n804), .B(new_n805), .Z(new_n806));
  NOR3_X1   g381(.A1(new_n794), .A2(new_n795), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n786), .A2(new_n787), .A3(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n787), .B1(new_n786), .B2(new_n807), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n771), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n810), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n812), .A2(KEYINPUT36), .A3(new_n808), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n770), .B1(new_n811), .B2(new_n813), .ZN(G311));
  NAND2_X1  g389(.A1(new_n811), .A2(new_n813), .ZN(new_n815));
  INV_X1    g390(.A(new_n770), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(G150));
  NAND2_X1  g392(.A1(new_n603), .A2(G559), .ZN(new_n818));
  INV_X1    g393(.A(G93), .ZN(new_n819));
  INV_X1    g394(.A(G55), .ZN(new_n820));
  OAI22_X1  g395(.A1(new_n522), .A2(new_n819), .B1(new_n524), .B2(new_n820), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n822), .A2(new_n510), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT108), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n552), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n825), .B2(new_n824), .ZN(new_n827));
  INV_X1    g402(.A(new_n824), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n828), .A2(KEYINPUT108), .A3(new_n552), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n818), .B(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT107), .B(KEYINPUT38), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT39), .ZN(new_n834));
  AOI21_X1  g409(.A(G860), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n834), .B2(new_n833), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n824), .A2(G860), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT37), .Z(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(G145));
  XNOR2_X1  g414(.A(new_n802), .B(KEYINPUT110), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n625), .ZN(new_n841));
  OAI21_X1  g416(.A(G2104), .B1(new_n480), .B2(G118), .ZN(new_n842));
  INV_X1    g417(.A(G106), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n842), .B1(new_n843), .B2(new_n480), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n487), .A2(G130), .ZN(new_n845));
  AOI211_X1 g420(.A(new_n844), .B(new_n845), .C1(G142), .C2(new_n478), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n841), .B(new_n846), .Z(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n499), .A2(G2105), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n502), .A2(new_n849), .A3(G2104), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n496), .B1(new_n482), .B2(new_n483), .ZN(new_n851));
  OAI21_X1  g426(.A(KEYINPUT109), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n497), .B1(new_n464), .B2(new_n465), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n502), .A2(new_n849), .A3(G2104), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT109), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n852), .A2(new_n856), .A3(new_n506), .A4(new_n507), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n745), .B(new_n857), .Z(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n694), .ZN(new_n859));
  MUX2_X1   g434(.A(new_n683), .B(new_n682), .S(new_n859), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n848), .B(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n620), .B(G160), .Z(new_n862));
  XNOR2_X1  g437(.A(G162), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n860), .B(new_n847), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(new_n863), .ZN(new_n867));
  INV_X1    g442(.A(G37), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n865), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g445(.A1(new_n824), .A2(new_n596), .ZN(new_n871));
  XNOR2_X1  g446(.A(G290), .B(new_n590), .ZN(new_n872));
  XNOR2_X1  g447(.A(G166), .B(new_n581), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(KEYINPUT111), .B2(KEYINPUT42), .ZN(new_n875));
  XOR2_X1   g450(.A(KEYINPUT111), .B(KEYINPUT42), .Z(new_n876));
  OAI21_X1  g451(.A(new_n875), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT112), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n611), .B(new_n830), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n602), .B(new_n570), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  AOI22_X1  g456(.A1(new_n877), .A2(new_n878), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n880), .B(KEYINPUT41), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n882), .B1(new_n879), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n877), .A2(new_n878), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n871), .B1(new_n887), .B2(new_n596), .ZN(G295));
  OAI21_X1  g463(.A(new_n871), .B1(new_n887), .B2(new_n596), .ZN(G331));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n890));
  NAND2_X1  g465(.A1(G286), .A2(G171), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(G286), .B2(new_n572), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n892), .B(new_n830), .Z(new_n893));
  NOR2_X1   g468(.A1(new_n893), .A2(new_n881), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT113), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n892), .B(new_n830), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n895), .B1(new_n896), .B2(new_n883), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n893), .A2(new_n884), .A3(KEYINPUT113), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT43), .B1(new_n899), .B2(new_n874), .ZN(new_n900));
  INV_X1    g475(.A(new_n874), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(new_n899), .B2(KEYINPUT114), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT114), .ZN(new_n903));
  AOI211_X1 g478(.A(new_n903), .B(new_n894), .C1(new_n897), .C2(new_n898), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n868), .B(new_n900), .C1(new_n902), .C2(new_n904), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n899), .A2(new_n874), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n894), .B1(new_n884), .B2(new_n893), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n868), .B1(new_n907), .B2(new_n874), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT43), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n890), .B1(new_n905), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n899), .A2(new_n874), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n913), .A2(new_n908), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n868), .B(new_n911), .C1(new_n902), .C2(new_n904), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n914), .B1(KEYINPUT43), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n910), .B1(new_n916), .B2(new_n890), .ZN(G397));
  NAND2_X1  g492(.A1(G160), .A2(G40), .ZN(new_n918));
  XOR2_X1   g493(.A(KEYINPUT115), .B(G1384), .Z(new_n919));
  NAND2_X1  g494(.A1(new_n857), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(KEYINPUT116), .B(KEYINPUT45), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n694), .B(G1996), .ZN(new_n923));
  INV_X1    g498(.A(G2067), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n745), .B(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  XOR2_X1   g501(.A(new_n802), .B(new_n805), .Z(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(G290), .B(new_n791), .ZN(new_n929));
  AOI211_X1 g504(.A(new_n918), .B(new_n922), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT50), .ZN(new_n931));
  INV_X1    g506(.A(G1384), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n857), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n508), .A2(new_n932), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT50), .ZN(new_n935));
  INV_X1    g510(.A(G40), .ZN(new_n936));
  AOI211_X1 g511(.A(new_n936), .B(new_n468), .C1(new_n474), .C2(G2105), .ZN(new_n937));
  INV_X1    g512(.A(G2084), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n933), .A2(new_n935), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n939), .B(KEYINPUT119), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT45), .B1(new_n857), .B2(new_n932), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT118), .B1(new_n941), .B2(new_n918), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT118), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n855), .B1(new_n853), .B2(new_n854), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n506), .A2(new_n507), .ZN(new_n947));
  AOI21_X1  g522(.A(G1384), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n943), .B(new_n937), .C1(new_n948), .C2(KEYINPUT45), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n934), .A2(new_n921), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n942), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G1966), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n940), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G8), .ZN(new_n956));
  NOR2_X1   g531(.A1(G168), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n941), .A2(new_n918), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n950), .B1(new_n959), .B2(new_n943), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n960), .A2(KEYINPUT53), .A3(new_n718), .A4(new_n942), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n933), .A2(new_n935), .A3(new_n937), .ZN(new_n962));
  INV_X1    g537(.A(G1961), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n857), .A2(KEYINPUT45), .A3(new_n919), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n965), .A2(new_n937), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n934), .A2(new_n921), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(new_n718), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT53), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n961), .A2(new_n964), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n971), .A2(KEYINPUT62), .A3(new_n572), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n956), .B1(new_n940), .B2(new_n954), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n973), .A2(KEYINPUT51), .A3(new_n957), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n957), .B1(new_n973), .B2(KEYINPUT123), .ZN(new_n977));
  AOI21_X1  g552(.A(G1966), .B1(new_n960), .B2(new_n942), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT119), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n939), .B(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(G8), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT123), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n976), .B1(new_n977), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n975), .B1(new_n984), .B2(KEYINPUT124), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT124), .ZN(new_n986));
  AOI211_X1 g561(.A(new_n986), .B(new_n976), .C1(new_n977), .C2(new_n983), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n958), .B(new_n972), .C1(new_n985), .C2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(G305), .A2(G1981), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n590), .A2(new_n675), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT49), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n989), .A2(KEYINPUT49), .A3(new_n990), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n857), .A2(new_n932), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n918), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n996), .A2(new_n956), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n993), .A2(new_n994), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT117), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n966), .A2(new_n967), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n774), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1002), .B1(G2090), .B2(new_n962), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(G8), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n575), .A2(G8), .A3(new_n576), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1005), .B(KEYINPUT55), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n508), .A2(new_n931), .A3(new_n932), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n937), .B(new_n1008), .C1(new_n948), .C2(new_n931), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1009), .A2(G2090), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1010), .B1(new_n774), .B2(new_n1001), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1006), .B1(new_n956), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1976), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n997), .B1(new_n1013), .B2(new_n581), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT52), .ZN(new_n1015));
  NAND2_X1  g590(.A1(G288), .A2(new_n1013), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1015), .B1(new_n1018), .B2(new_n1014), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1000), .A2(new_n1007), .A3(new_n1012), .A4(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  OAI211_X1 g597(.A(KEYINPUT123), .B(G8), .C1(new_n978), .C2(new_n980), .ZN(new_n1023));
  INV_X1    g598(.A(new_n957), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n973), .A2(KEYINPUT123), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT51), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n974), .B1(new_n1027), .B2(new_n986), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n984), .A2(KEYINPUT124), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1028), .A2(new_n1029), .B1(new_n957), .B2(new_n955), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n561), .A2(new_n568), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1031), .B1(new_n561), .B2(new_n568), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1009), .A2(new_n766), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT56), .B(G2072), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n966), .A2(new_n967), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1034), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1039));
  INV_X1    g614(.A(G1348), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n962), .A2(new_n1040), .B1(new_n996), .B2(new_n924), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(new_n602), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1038), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT61), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1039), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1045), .B1(new_n1046), .B2(new_n1038), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1037), .A2(new_n1035), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1034), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1050), .A2(KEYINPUT61), .A3(new_n1039), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n962), .A2(new_n1040), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n996), .A2(new_n924), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1052), .A2(new_n1053), .A3(new_n602), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT60), .B1(new_n1042), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n602), .A2(KEYINPUT60), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1041), .A2(new_n1056), .ZN(new_n1057));
  AND4_X1   g632(.A1(new_n1047), .A2(new_n1051), .A3(new_n1055), .A4(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G1996), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n965), .A2(new_n967), .A3(new_n937), .A4(new_n1059), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n1060), .A2(KEYINPUT120), .ZN(new_n1061));
  XOR2_X1   g636(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n1062));
  XNOR2_X1  g637(.A(new_n1062), .B(G1341), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(new_n918), .B2(new_n995), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1060), .A2(KEYINPUT120), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1061), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT122), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1066), .A2(new_n552), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1069), .B1(new_n1066), .B2(new_n552), .ZN(new_n1072));
  OAI22_X1  g647(.A1(new_n1071), .A2(new_n1072), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1044), .B1(new_n1058), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n572), .B1(new_n969), .B2(new_n968), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1075), .A2(new_n961), .A3(new_n964), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n966), .A2(KEYINPUT53), .A3(new_n718), .A4(new_n922), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1077), .A2(new_n964), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1078), .A2(new_n970), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1076), .B1(new_n1079), .B2(new_n734), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n971), .A2(new_n572), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT54), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1080), .A2(KEYINPUT54), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI22_X1  g658(.A1(new_n1074), .A2(new_n1083), .B1(KEYINPUT62), .B2(new_n1081), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n988), .B(new_n1022), .C1(new_n1030), .C2(new_n1084), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1000), .A2(new_n1020), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1007), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n997), .ZN(new_n1089));
  NOR2_X1   g664(.A1(G288), .A2(G1976), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n1000), .A2(new_n1090), .B1(new_n675), .B2(new_n590), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1088), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT63), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n981), .A2(G286), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1093), .B1(new_n1021), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1093), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1086), .A2(new_n1007), .A3(new_n1094), .A4(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1092), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n930), .B1(new_n1085), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n925), .A2(new_n694), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n922), .A2(new_n918), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NOR3_X1   g678(.A1(new_n922), .A2(G1996), .A3(new_n918), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT46), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n1104), .A2(KEYINPUT46), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1103), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1107), .B(KEYINPUT47), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n803), .A2(new_n805), .ZN(new_n1109));
  OAI22_X1  g684(.A1(new_n926), .A2(new_n1109), .B1(G2067), .B2(new_n745), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1102), .B1(new_n926), .B2(new_n927), .ZN(new_n1111));
  NOR2_X1   g686(.A1(G290), .A2(G1986), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n1102), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT125), .B(KEYINPUT48), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1114), .B(KEYINPUT126), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1113), .B(new_n1115), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1102), .A2(new_n1110), .B1(new_n1111), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1108), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(KEYINPUT127), .B1(new_n1100), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT127), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1118), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1091), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1123), .A2(new_n997), .B1(new_n1087), .B2(new_n1086), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n958), .B1(new_n985), .B2(new_n987), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1081), .A2(KEYINPUT62), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1072), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1128), .A2(new_n1070), .B1(KEYINPUT122), .B2(KEYINPUT59), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1047), .A2(new_n1051), .A3(new_n1055), .A4(new_n1057), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1043), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1080), .A2(KEYINPUT54), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1127), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1021), .B1(new_n1126), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1125), .B1(new_n1136), .B2(new_n988), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1120), .B(new_n1121), .C1(new_n1137), .C2(new_n930), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1119), .A2(new_n1138), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g714(.A1(G229), .A2(new_n462), .A3(G401), .A4(G227), .ZN(new_n1141));
  NAND2_X1  g715(.A1(new_n1141), .A2(new_n869), .ZN(new_n1142));
  NOR2_X1   g716(.A1(new_n1142), .A2(new_n916), .ZN(G308));
  AND2_X1   g717(.A1(new_n915), .A2(KEYINPUT43), .ZN(new_n1144));
  OAI211_X1 g718(.A(new_n869), .B(new_n1141), .C1(new_n1144), .C2(new_n914), .ZN(G225));
endmodule


