//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 0 0 1 1 0 1 1 0 1 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n187));
  INV_X1    g001(.A(G221), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT9), .B(G234), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n188), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(G110), .B(G140), .ZN(new_n194));
  INV_X1    g008(.A(G953), .ZN(new_n195));
  AND2_X1   g009(.A1(new_n195), .A2(G227), .ZN(new_n196));
  XNOR2_X1  g010(.A(new_n194), .B(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT3), .B1(new_n199), .B2(G107), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G104), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n199), .A2(G107), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n200), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT79), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT79), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n200), .A2(new_n203), .A3(new_n207), .A4(new_n204), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(G101), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G101), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n200), .A2(new_n203), .A3(new_n210), .A4(new_n204), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT80), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n206), .A2(KEYINPUT80), .A3(G101), .A4(new_n208), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(KEYINPUT4), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G143), .ZN(new_n217));
  INV_X1    g031(.A(G143), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G146), .ZN(new_n219));
  AND2_X1   g033(.A1(KEYINPUT0), .A2(G128), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n217), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  OR2_X1    g035(.A1(KEYINPUT0), .A2(G128), .ZN(new_n222));
  NAND2_X1  g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(G143), .B(G146), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n221), .B(KEYINPUT64), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n217), .A2(new_n219), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT64), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n227), .A2(new_n228), .A3(new_n223), .A4(new_n222), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n206), .A2(new_n231), .A3(G101), .A4(new_n208), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n215), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT11), .ZN(new_n234));
  INV_X1    g048(.A(G134), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n234), .B1(new_n235), .B2(G137), .ZN(new_n236));
  INV_X1    g050(.A(G137), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(KEYINPUT11), .A3(G134), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n235), .A2(G137), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n236), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G131), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT65), .B(G131), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n242), .A2(new_n236), .A3(new_n238), .A4(new_n239), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n199), .A2(G107), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n202), .A2(G104), .ZN(new_n247));
  OAI21_X1  g061(.A(G101), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n211), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT1), .B1(new_n218), .B2(G146), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT81), .ZN(new_n251));
  OAI21_X1  g065(.A(G128), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT81), .B1(new_n217), .B2(KEYINPUT1), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n227), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n255));
  AND4_X1   g069(.A1(new_n255), .A2(new_n217), .A3(new_n219), .A4(G128), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n249), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n259));
  INV_X1    g073(.A(G128), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n260), .B1(new_n217), .B2(KEYINPUT1), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT66), .B1(new_n261), .B2(new_n225), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n250), .A2(G128), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT66), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n264), .A3(new_n227), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n256), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n211), .A2(new_n248), .A3(KEYINPUT10), .ZN(new_n267));
  OAI22_X1  g081(.A1(new_n258), .A2(new_n259), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n233), .A2(new_n245), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n232), .A2(new_n230), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n231), .B1(new_n209), .B2(new_n212), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n271), .B1(new_n272), .B2(new_n214), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n244), .B1(new_n273), .B2(new_n268), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n198), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  AOI221_X4 g089(.A(new_n256), .B1(new_n211), .B2(new_n248), .C1(new_n262), .C2(new_n265), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n244), .B1(new_n276), .B2(new_n258), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT12), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n249), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n255), .B1(G143), .B2(new_n216), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n260), .B1(new_n281), .B2(KEYINPUT81), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n250), .A2(new_n251), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n225), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n280), .B1(new_n284), .B2(new_n256), .ZN(new_n285));
  NOR3_X1   g099(.A1(new_n261), .A2(new_n225), .A3(KEYINPUT66), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n264), .B1(new_n263), .B2(new_n227), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n257), .B(new_n249), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(KEYINPUT12), .A3(new_n244), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n279), .A2(KEYINPUT83), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT83), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT12), .B1(new_n289), .B2(new_n244), .ZN(new_n293));
  AOI211_X1 g107(.A(new_n278), .B(new_n245), .C1(new_n285), .C2(new_n288), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n273), .A2(new_n268), .A3(new_n244), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT84), .B1(new_n297), .B2(new_n197), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT84), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n270), .A2(new_n299), .A3(new_n198), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n296), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n275), .B1(new_n301), .B2(KEYINPUT85), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT85), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n296), .A2(new_n298), .A3(new_n300), .A4(new_n303), .ZN(new_n304));
  AOI211_X1 g118(.A(G469), .B(G902), .C1(new_n302), .C2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G469), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n293), .A2(new_n294), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n197), .B1(new_n307), .B2(new_n297), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n270), .A2(new_n274), .A3(new_n198), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n306), .B1(new_n310), .B2(new_n191), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n193), .B1(new_n305), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(G214), .B1(G237), .B2(G902), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n313), .B(KEYINPUT86), .ZN(new_n314));
  OAI21_X1  g128(.A(G210), .B1(G237), .B2(G902), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT90), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n230), .A2(G125), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n319), .B1(G125), .B2(new_n266), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n195), .A2(G224), .ZN(new_n321));
  XOR2_X1   g135(.A(new_n321), .B(KEYINPUT89), .Z(new_n322));
  XNOR2_X1  g136(.A(new_n320), .B(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G119), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G116), .ZN(new_n325));
  INV_X1    g139(.A(G116), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G119), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT2), .B(G113), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n328), .B(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n232), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n331), .B1(new_n272), .B2(new_n214), .ZN(new_n332));
  OR2_X1    g146(.A1(new_n328), .A2(new_n329), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n325), .A2(new_n327), .A3(KEYINPUT5), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT87), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT5), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(new_n324), .A3(G116), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n334), .A2(new_n335), .A3(G113), .A4(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n334), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(G113), .ZN(new_n340));
  OAI21_X1  g154(.A(KEYINPUT87), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AND4_X1   g155(.A1(new_n333), .A2(new_n280), .A3(new_n338), .A4(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(G110), .B(G122), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NOR3_X1   g158(.A1(new_n332), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT6), .ZN(new_n346));
  INV_X1    g160(.A(new_n331), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n342), .B1(new_n215), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n344), .A2(KEYINPUT88), .ZN(new_n349));
  OAI22_X1  g163(.A1(new_n345), .A2(new_n346), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n349), .ZN(new_n351));
  OAI211_X1 g165(.A(KEYINPUT6), .B(new_n351), .C1(new_n332), .C2(new_n342), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n323), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n320), .A2(KEYINPUT7), .A3(new_n321), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n333), .B1(new_n339), .B2(new_n340), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n280), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n341), .A2(new_n333), .A3(new_n249), .A4(new_n338), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n343), .B(KEYINPUT8), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n321), .A2(KEYINPUT7), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n319), .B(new_n360), .C1(G125), .C2(new_n266), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n354), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n191), .B1(new_n362), .B2(new_n345), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n318), .B1(new_n353), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n346), .B1(new_n348), .B2(new_n343), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n348), .A2(new_n349), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n352), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n323), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n363), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n317), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n314), .B1(new_n364), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT97), .ZN(new_n373));
  XNOR2_X1  g187(.A(G113), .B(G122), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n374), .B(new_n199), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT16), .ZN(new_n377));
  INV_X1    g191(.A(G140), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(G125), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(G125), .ZN(new_n380));
  INV_X1    g194(.A(G125), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G140), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  OAI211_X1 g197(.A(G146), .B(new_n379), .C1(new_n383), .C2(new_n377), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT77), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n380), .A2(new_n382), .A3(KEYINPUT77), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT19), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n383), .A2(KEYINPUT19), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n384), .B1(new_n391), .B2(G146), .ZN(new_n392));
  XOR2_X1   g206(.A(KEYINPUT65), .B(G131), .Z(new_n393));
  INV_X1    g207(.A(G237), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT70), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT70), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G237), .ZN(new_n397));
  AOI21_X1  g211(.A(G953), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(KEYINPUT91), .B(G143), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(G214), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n398), .A2(G214), .B1(KEYINPUT91), .B2(G143), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n393), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n398), .A2(G214), .ZN(new_n404));
  NAND2_X1  g218(.A1(KEYINPUT91), .A2(G143), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(new_n242), .A3(new_n400), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n392), .B1(new_n403), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT18), .ZN(new_n409));
  INV_X1    g223(.A(G131), .ZN(new_n410));
  NOR3_X1   g224(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT92), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n412), .B1(new_n401), .B2(new_n402), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n406), .A2(new_n411), .A3(new_n400), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n386), .A2(new_n216), .A3(new_n387), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n383), .A2(G146), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n413), .A2(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n376), .B1(new_n408), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n379), .B1(new_n383), .B2(new_n377), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n216), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n384), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n242), .B1(new_n406), .B2(new_n400), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n421), .B1(new_n422), .B2(KEYINPUT17), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT17), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n403), .A2(new_n407), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n417), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n427), .A3(new_n375), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n418), .A2(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(G475), .A2(G902), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT20), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n429), .A2(new_n433), .A3(new_n430), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n426), .A2(new_n427), .A3(new_n375), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n375), .B1(new_n426), .B2(new_n427), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n191), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AOI22_X1  g251(.A1(new_n432), .A2(new_n434), .B1(G475), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n195), .A2(G952), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n439), .B1(G234), .B2(G237), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  XOR2_X1   g255(.A(KEYINPUT21), .B(G898), .Z(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(KEYINPUT96), .ZN(new_n443));
  INV_X1    g257(.A(G234), .ZN(new_n444));
  OAI211_X1 g258(.A(G902), .B(G953), .C1(new_n444), .C2(new_n394), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(KEYINPUT95), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n441), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n218), .A2(G128), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n260), .A2(G143), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n449), .A2(new_n450), .A3(new_n235), .ZN(new_n451));
  XNOR2_X1  g265(.A(G116), .B(G122), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G107), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n202), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n451), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT13), .ZN(new_n457));
  OAI21_X1  g271(.A(KEYINPUT93), .B1(new_n449), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n449), .A2(new_n457), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n450), .A3(new_n459), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n449), .A2(KEYINPUT93), .A3(new_n457), .ZN(new_n461));
  OAI21_X1  g275(.A(G134), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n326), .A2(KEYINPUT14), .A3(G122), .ZN(new_n464));
  OAI211_X1 g278(.A(G107), .B(new_n464), .C1(new_n453), .C2(KEYINPUT14), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n235), .B1(new_n449), .B2(new_n450), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n465), .B(new_n455), .C1(new_n451), .C2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G217), .ZN(new_n468));
  NOR3_X1   g282(.A1(new_n189), .A2(new_n468), .A3(G953), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n463), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n469), .B1(new_n463), .B2(new_n467), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n191), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G478), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n473), .A2(KEYINPUT15), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  OAI221_X1 g289(.A(new_n191), .B1(KEYINPUT15), .B2(new_n473), .C1(new_n470), .C2(new_n471), .ZN(new_n476));
  AOI21_X1  g290(.A(KEYINPUT94), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n475), .A2(new_n476), .A3(KEYINPUT94), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n448), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n373), .B1(new_n438), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n437), .A2(G475), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n433), .B1(new_n429), .B2(new_n430), .ZN(new_n483));
  INV_X1    g297(.A(new_n430), .ZN(new_n484));
  AOI211_X1 g298(.A(KEYINPUT20), .B(new_n484), .C1(new_n418), .C2(new_n428), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n482), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n475), .A2(KEYINPUT94), .A3(new_n476), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n447), .B1(new_n487), .B2(new_n477), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n486), .A2(new_n488), .A3(KEYINPUT97), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n372), .B1(new_n481), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n187), .B1(new_n312), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(KEYINPUT72), .B(KEYINPUT32), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n257), .B1(new_n286), .B2(new_n287), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT68), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n235), .A2(G137), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n237), .A2(G134), .ZN(new_n496));
  OAI21_X1  g310(.A(G131), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n243), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n497), .B1(new_n240), .B2(new_n393), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT68), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n493), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n330), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n230), .A2(new_n244), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT28), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT28), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n501), .A2(new_n506), .A3(new_n502), .A4(new_n503), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n503), .B1(new_n499), .B2(new_n266), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n505), .A2(new_n507), .B1(new_n330), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n398), .A2(G210), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(KEYINPUT27), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT26), .B(G101), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n511), .B(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n501), .A2(KEYINPUT30), .A3(new_n503), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT69), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT69), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n501), .A2(new_n517), .A3(KEYINPUT30), .A4(new_n503), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n499), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n493), .A2(new_n520), .B1(new_n244), .B2(new_n230), .ZN(new_n521));
  OAI21_X1  g335(.A(KEYINPUT67), .B1(new_n521), .B2(KEYINPUT30), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT67), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT30), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n508), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n519), .A2(new_n330), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n527), .A2(new_n513), .A3(new_n504), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT31), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n527), .A2(KEYINPUT31), .A3(new_n513), .A4(new_n504), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n514), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(G472), .A2(G902), .ZN(new_n533));
  XOR2_X1   g347(.A(new_n533), .B(KEYINPUT71), .Z(new_n534));
  OAI21_X1  g348(.A(new_n492), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n514), .ZN(new_n536));
  INV_X1    g350(.A(new_n504), .ZN(new_n537));
  AOI22_X1  g351(.A1(new_n516), .A2(new_n518), .B1(new_n522), .B2(new_n525), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n537), .B1(new_n538), .B2(new_n330), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT31), .B1(new_n539), .B2(new_n513), .ZN(new_n540));
  AND4_X1   g354(.A1(KEYINPUT31), .A2(new_n527), .A3(new_n513), .A4(new_n504), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n536), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n534), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(KEYINPUT32), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n505), .A2(new_n507), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n501), .A2(new_n503), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n330), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n513), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT29), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(G902), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n513), .B1(new_n527), .B2(new_n504), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n508), .A2(new_n330), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n545), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n550), .B1(new_n555), .B2(new_n549), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n552), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT73), .B1(new_n557), .B2(G472), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT73), .ZN(new_n559));
  INV_X1    g373(.A(G472), .ZN(new_n560));
  AOI21_X1  g374(.A(KEYINPUT29), .B1(new_n509), .B2(new_n513), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n561), .B1(new_n539), .B2(new_n513), .ZN(new_n562));
  AOI211_X1 g376(.A(new_n559), .B(new_n560), .C1(new_n562), .C2(new_n552), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n535), .B(new_n544), .C1(new_n558), .C2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT22), .B(G137), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n188), .A2(new_n444), .A3(G953), .ZN(new_n566));
  XOR2_X1   g380(.A(new_n565), .B(new_n566), .Z(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(KEYINPUT23), .B1(new_n260), .B2(G119), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT74), .B1(new_n324), .B2(G128), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n569), .B(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(G110), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT75), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT23), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n574), .B1(new_n324), .B2(G128), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(new_n570), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT75), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n576), .A2(new_n577), .A3(G110), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(G119), .B(G128), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT24), .B(G110), .ZN(new_n582));
  OR2_X1    g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n579), .A2(new_n583), .A3(new_n421), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n582), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT76), .B(G110), .Z(new_n586));
  OAI21_X1  g400(.A(new_n585), .B1(new_n576), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(new_n384), .A3(new_n415), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n568), .B1(new_n584), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n579), .A2(new_n583), .A3(new_n421), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n591), .A2(new_n588), .A3(new_n567), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n590), .A2(new_n592), .A3(new_n191), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT25), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n590), .A2(new_n592), .A3(KEYINPUT25), .A4(new_n191), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n595), .A2(KEYINPUT78), .A3(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT78), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n593), .A2(new_n598), .A3(new_n594), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n468), .B1(G234), .B2(new_n191), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n590), .A2(new_n592), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n600), .A2(G902), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n314), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n353), .A2(new_n318), .A3(new_n363), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n317), .B1(new_n369), .B2(new_n370), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n438), .A2(new_n480), .A3(new_n373), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT97), .B1(new_n486), .B2(new_n488), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n301), .A2(KEYINPUT85), .ZN(new_n615));
  INV_X1    g429(.A(new_n275), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n304), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n617), .A2(new_n306), .A3(new_n191), .ZN(new_n618));
  INV_X1    g432(.A(new_n311), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n192), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n614), .A2(new_n620), .A3(KEYINPUT98), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n491), .A2(new_n564), .A3(new_n607), .A4(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G101), .ZN(G3));
  OAI21_X1  g437(.A(G472), .B1(new_n532), .B2(G902), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n542), .A2(new_n543), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n607), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n353), .A2(new_n316), .A3(new_n363), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n315), .B1(new_n369), .B2(new_n370), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n608), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OR2_X1    g445(.A1(new_n470), .A2(new_n471), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n632), .A2(new_n473), .A3(new_n191), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n473), .A2(new_n191), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n632), .B(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n636), .B1(new_n638), .B2(G478), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n486), .A2(new_n639), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n631), .A2(new_n448), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n628), .A2(new_n620), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  INV_X1    g458(.A(KEYINPUT99), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n482), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n437), .A2(KEYINPUT99), .A3(G475), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n432), .A2(new_n434), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n487), .A2(new_n477), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n648), .A2(new_n649), .A3(new_n650), .A4(new_n447), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n651), .A2(new_n631), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n628), .A2(new_n620), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT35), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n584), .A2(new_n589), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n568), .A2(KEYINPUT36), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  OR2_X1    g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OAI22_X1  g475(.A1(new_n597), .A2(new_n601), .B1(new_n605), .B2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n656), .B1(new_n626), .B2(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n624), .A2(KEYINPUT100), .A3(new_n625), .A4(new_n662), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n491), .A2(new_n621), .A3(new_n664), .A4(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT37), .B(G110), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  NOR2_X1   g482(.A1(new_n446), .A2(G900), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT101), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n441), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n669), .A2(KEYINPUT101), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n648), .A2(new_n649), .A3(new_n650), .A4(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n631), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n564), .A2(new_n620), .A3(new_n662), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  NAND3_X1  g492(.A1(new_n486), .A2(new_n650), .A3(new_n608), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n662), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT104), .ZN(new_n681));
  INV_X1    g495(.A(new_n528), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n513), .B1(new_n547), .B2(new_n504), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT103), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n191), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(G472), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n535), .A2(new_n544), .A3(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n609), .A2(new_n610), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n681), .A2(new_n687), .A3(new_n690), .ZN(new_n691));
  OR2_X1    g505(.A1(new_n691), .A2(KEYINPUT105), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT106), .B(KEYINPUT39), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n673), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n620), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n695), .B(KEYINPUT40), .Z(new_n696));
  NAND2_X1  g510(.A1(new_n691), .A2(KEYINPUT105), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n692), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G143), .ZN(G45));
  NOR3_X1   g513(.A1(new_n631), .A2(new_n640), .A3(new_n673), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n564), .A2(new_n620), .A3(new_n662), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT107), .B(G146), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G48));
  AOI21_X1  g517(.A(new_n306), .B1(new_n617), .B2(new_n191), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n305), .A2(new_n704), .A3(new_n192), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n705), .A2(new_n564), .A3(new_n607), .A4(new_n641), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT41), .B(G113), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G15));
  NAND4_X1  g522(.A1(new_n705), .A2(new_n564), .A3(new_n607), .A4(new_n652), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G116), .ZN(G18));
  NOR4_X1   g524(.A1(new_n305), .A2(new_n704), .A3(new_n631), .A4(new_n192), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n612), .A2(new_n613), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n711), .A2(new_n564), .A3(new_n712), .A4(new_n662), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G119), .ZN(G21));
  OAI22_X1  g528(.A1(new_n540), .A2(new_n541), .B1(new_n513), .B2(new_n548), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n543), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n624), .A2(new_n607), .A3(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n629), .A2(new_n630), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n679), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n717), .A2(new_n705), .A3(new_n447), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G122), .ZN(G24));
  NOR2_X1   g535(.A1(new_n640), .A2(new_n673), .ZN(new_n722));
  AND4_X1   g536(.A1(new_n624), .A2(new_n716), .A3(new_n722), .A4(new_n662), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n711), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n308), .A2(KEYINPUT108), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n728), .B(new_n197), .C1(new_n307), .C2(new_n297), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n727), .A2(new_n309), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n306), .B1(new_n730), .B2(new_n191), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n618), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n192), .A2(new_n314), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n364), .A2(new_n371), .A3(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n726), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  AOI211_X1 g551(.A(KEYINPUT109), .B(new_n735), .C1(new_n618), .C2(new_n732), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT32), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n740), .B1(new_n532), .B2(new_n534), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n741), .B(new_n544), .C1(new_n558), .C2(new_n563), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n607), .A3(new_n722), .ZN(new_n743));
  OAI21_X1  g557(.A(KEYINPUT42), .B1(new_n739), .B2(new_n743), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n535), .A2(new_n544), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n563), .A2(new_n558), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n627), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(G902), .B1(new_n302), .B2(new_n304), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n731), .B1(new_n749), .B2(new_n306), .ZN(new_n750));
  OAI21_X1  g564(.A(KEYINPUT109), .B1(new_n750), .B2(new_n735), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n733), .A2(new_n726), .A3(new_n736), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT42), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n748), .A2(new_n753), .A3(new_n754), .A4(new_n722), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n744), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(new_n410), .ZN(G33));
  INV_X1    g571(.A(new_n675), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n748), .A2(new_n753), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G134), .ZN(G36));
  NAND2_X1  g574(.A1(new_n688), .A2(new_n608), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n438), .A2(new_n639), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT43), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n764), .A2(KEYINPUT111), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n639), .B(KEYINPUT110), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n763), .B1(new_n766), .B2(new_n486), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n764), .A2(KEYINPUT111), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n765), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n769), .A2(new_n626), .A3(new_n662), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT44), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n761), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT45), .B1(new_n308), .B2(new_n309), .ZN(new_n773));
  INV_X1    g587(.A(new_n730), .ZN(new_n774));
  AOI211_X1 g588(.A(new_n306), .B(new_n773), .C1(new_n774), .C2(KEYINPUT45), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n306), .A2(new_n191), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n777), .A2(KEYINPUT46), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(KEYINPUT46), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n618), .A3(new_n779), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n780), .A2(new_n193), .A3(new_n694), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n772), .B(new_n781), .C1(new_n771), .C2(new_n770), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G137), .ZN(G39));
  INV_X1    g597(.A(new_n761), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n627), .A3(new_n722), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(new_n564), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n780), .A2(KEYINPUT47), .A3(new_n193), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT47), .B1(new_n780), .B2(new_n193), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G140), .ZN(G42));
  NAND3_X1  g604(.A1(new_n769), .A2(new_n440), .A3(new_n717), .ZN(new_n791));
  INV_X1    g605(.A(new_n705), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n791), .A2(new_n631), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n439), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n607), .A2(new_n440), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n792), .A2(new_n687), .A3(new_n761), .A4(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(new_n486), .A3(new_n639), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT48), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n798), .A2(KEYINPUT119), .ZN(new_n799));
  AND4_X1   g613(.A1(new_n440), .A2(new_n769), .A3(new_n705), .A4(new_n784), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n742), .A2(new_n607), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n800), .B(new_n801), .C1(KEYINPUT119), .C2(new_n798), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n794), .B(new_n797), .C1(new_n799), .C2(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n803), .B1(new_n799), .B2(new_n802), .ZN(new_n804));
  NOR4_X1   g618(.A1(new_n791), .A2(new_n608), .A3(new_n690), .A4(new_n792), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(KEYINPUT50), .Z(new_n806));
  NOR2_X1   g620(.A1(new_n787), .A2(new_n788), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n305), .A2(new_n704), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n192), .ZN(new_n809));
  AOI211_X1 g623(.A(new_n761), .B(new_n791), .C1(new_n807), .C2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n800), .A2(new_n624), .A3(new_n662), .A4(new_n716), .ZN(new_n811));
  INV_X1    g625(.A(new_n639), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n796), .A2(new_n438), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n806), .A2(new_n810), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n816));
  OR3_X1    g630(.A1(new_n806), .A2(new_n810), .A3(new_n816), .ZN(new_n817));
  XOR2_X1   g631(.A(new_n814), .B(KEYINPUT118), .Z(new_n818));
  OAI221_X1 g632(.A(new_n804), .B1(new_n815), .B2(KEYINPUT51), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT114), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n640), .A2(new_n448), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n628), .A2(new_n620), .A3(new_n372), .A4(new_n821), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n622), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n820), .B1(new_n622), .B2(new_n822), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n475), .A2(new_n476), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n438), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n826), .A2(new_n448), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n628), .A2(new_n620), .A3(new_n372), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n666), .A2(new_n828), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n823), .A2(new_n824), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n753), .A2(new_n723), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n648), .A2(new_n649), .ZN(new_n832));
  NOR4_X1   g646(.A1(new_n761), .A2(new_n832), .A3(new_n825), .A4(new_n673), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n833), .A2(new_n564), .A3(new_n620), .A4(new_n662), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n759), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n713), .A2(new_n706), .A3(new_n709), .A4(new_n720), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n756), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n724), .A2(new_n677), .A3(new_n701), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n662), .A2(new_n192), .A3(new_n673), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n687), .A2(new_n719), .A3(new_n733), .A4(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n838), .A2(KEYINPUT52), .A3(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n724), .A2(new_n677), .A3(new_n701), .A4(new_n840), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n830), .A2(new_n837), .A3(new_n845), .ZN(new_n846));
  XOR2_X1   g660(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n847));
  NOR2_X1   g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT115), .B1(new_n842), .B2(new_n843), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n842), .A2(new_n843), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n842), .A2(KEYINPUT115), .A3(new_n843), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n830), .B(new_n837), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n848), .B1(new_n849), .B2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n744), .A2(new_n755), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n759), .A2(new_n831), .A3(new_n834), .ZN(new_n858));
  INV_X1    g672(.A(new_n836), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n312), .A2(new_n490), .A3(new_n187), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT98), .B1(new_n614), .B2(new_n620), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n535), .A2(new_n544), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n607), .B1(new_n863), .B2(new_n746), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n861), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n822), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT114), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n622), .A2(new_n820), .A3(new_n822), .ZN(new_n868));
  INV_X1    g682(.A(new_n829), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n860), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT115), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n844), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n841), .ZN(new_n874));
  INV_X1    g688(.A(new_n853), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n871), .A2(new_n876), .A3(KEYINPUT53), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n846), .A2(new_n847), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XOR2_X1   g693(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  OAI22_X1  g695(.A1(new_n855), .A2(new_n856), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  OAI22_X1  g696(.A1(new_n819), .A2(new_n882), .B1(G952), .B2(G953), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n808), .B(KEYINPUT49), .Z(new_n884));
  NAND2_X1  g698(.A1(new_n607), .A2(new_n734), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT112), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n762), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n887), .B1(new_n886), .B2(new_n885), .ZN(new_n888));
  NOR4_X1   g702(.A1(new_n884), .A2(new_n888), .A3(new_n687), .A4(new_n690), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT113), .Z(new_n890));
  NAND2_X1  g704(.A1(new_n883), .A2(new_n890), .ZN(G75));
  AOI21_X1  g705(.A(new_n191), .B1(new_n877), .B2(new_n878), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n892), .A2(G210), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(KEYINPUT56), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n367), .B(new_n323), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT55), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n195), .A2(G952), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  XNOR2_X1  g713(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n899), .B1(new_n893), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n897), .A2(new_n902), .ZN(G51));
  XNOR2_X1  g717(.A(new_n879), .B(new_n880), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n776), .B(KEYINPUT57), .Z(new_n905));
  OAI21_X1  g719(.A(new_n617), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n892), .A2(new_n775), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n898), .B1(new_n906), .B2(new_n907), .ZN(G54));
  NAND3_X1  g722(.A1(new_n892), .A2(KEYINPUT58), .A3(G475), .ZN(new_n909));
  INV_X1    g723(.A(new_n429), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n909), .A2(KEYINPUT121), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n899), .B1(new_n909), .B2(new_n910), .ZN(new_n912));
  AOI21_X1  g726(.A(KEYINPUT121), .B1(new_n909), .B2(new_n910), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(G60));
  XNOR2_X1  g728(.A(new_n634), .B(KEYINPUT59), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n904), .A2(new_n638), .A3(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n638), .ZN(new_n917));
  INV_X1    g731(.A(new_n915), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n917), .B1(new_n882), .B2(new_n918), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n916), .A2(new_n919), .A3(new_n898), .ZN(G63));
  INV_X1    g734(.A(KEYINPUT124), .ZN(new_n921));
  NAND2_X1  g735(.A1(G217), .A2(G902), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT60), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n923), .B1(new_n877), .B2(new_n878), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n603), .B(KEYINPUT122), .Z(new_n925));
  OAI21_X1  g739(.A(new_n899), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI211_X1 g740(.A(new_n661), .B(new_n923), .C1(new_n877), .C2(new_n878), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n921), .B1(new_n928), .B2(KEYINPUT61), .ZN(new_n929));
  INV_X1    g743(.A(new_n661), .ZN(new_n930));
  INV_X1    g744(.A(new_n923), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n854), .A2(new_n849), .ZN(new_n932));
  INV_X1    g746(.A(new_n847), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n871), .B2(new_n845), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n930), .B(new_n931), .C1(new_n932), .C2(new_n934), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n935), .B(new_n899), .C1(new_n924), .C2(new_n925), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n936), .A2(KEYINPUT124), .A3(new_n937), .ZN(new_n938));
  OAI211_X1 g752(.A(KEYINPUT123), .B(new_n937), .C1(new_n926), .C2(new_n927), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT123), .B1(new_n936), .B2(new_n937), .ZN(new_n941));
  OAI22_X1  g755(.A1(new_n929), .A2(new_n938), .B1(new_n940), .B2(new_n941), .ZN(G66));
  AOI21_X1  g756(.A(new_n195), .B1(new_n443), .B2(G224), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n830), .A2(new_n859), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT125), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n943), .B1(new_n946), .B2(new_n195), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n350), .B(new_n352), .C1(G898), .C2(new_n195), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n947), .B(new_n948), .Z(G69));
  XOR2_X1   g763(.A(new_n538), .B(new_n391), .Z(new_n950));
  NAND2_X1  g764(.A1(new_n698), .A2(new_n838), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(KEYINPUT62), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n782), .A2(new_n789), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT62), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n698), .A2(new_n954), .A3(new_n838), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n761), .B1(new_n640), .B2(new_n826), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n748), .A2(new_n620), .A3(new_n694), .A4(new_n956), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n952), .A2(new_n953), .A3(new_n955), .A4(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n950), .B1(new_n958), .B2(new_n195), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n959), .A2(KEYINPUT126), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(KEYINPUT126), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n781), .A2(new_n719), .A3(new_n801), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n962), .A2(new_n759), .A3(new_n838), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n953), .A2(new_n857), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n195), .ZN(new_n965));
  INV_X1    g779(.A(new_n950), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n966), .B1(G900), .B2(G953), .ZN(new_n967));
  AOI21_X1  g781(.A(KEYINPUT127), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n960), .A2(new_n961), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n195), .B1(G227), .B2(G900), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n970), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n960), .A2(new_n972), .A3(new_n961), .A4(new_n968), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n971), .A2(new_n973), .ZN(G72));
  NAND2_X1  g788(.A1(G472), .A2(G902), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT63), .Z(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(new_n946), .B2(new_n958), .ZN(new_n977));
  INV_X1    g791(.A(new_n539), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n977), .A2(new_n513), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n945), .A2(new_n964), .ZN(new_n980));
  AOI211_X1 g794(.A(new_n513), .B(new_n978), .C1(new_n980), .C2(new_n976), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n976), .B1(new_n682), .B2(new_n553), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n899), .B1(new_n855), .B2(new_n982), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n979), .A2(new_n981), .A3(new_n983), .ZN(G57));
endmodule


