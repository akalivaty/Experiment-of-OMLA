//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 1 0 1 0 0 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n562, new_n564,
    new_n565, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  XNOR2_X1  g030(.A(G325), .B(KEYINPUT67), .ZN(G261));
  AOI22_X1  g031(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  OR2_X1    g032(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n458));
  NAND2_X1  g033(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  AND3_X1   g039(.A1(new_n462), .A2(new_n464), .A3(KEYINPUT69), .ZN(new_n465));
  AOI21_X1  g040(.A(KEYINPUT69), .B1(new_n462), .B2(new_n464), .ZN(new_n466));
  OAI21_X1  g041(.A(G125), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n460), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n462), .A2(new_n464), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(new_n460), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT70), .ZN(new_n477));
  INV_X1    g052(.A(G101), .ZN(new_n478));
  OAI22_X1  g053(.A1(new_n473), .A2(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n470), .A2(new_n479), .ZN(G160));
  OAI221_X1 g055(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n460), .C2(G112), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT71), .ZN(new_n482));
  OR2_X1    g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n481), .A2(new_n482), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n471), .A2(G2105), .ZN(new_n485));
  AOI22_X1  g060(.A1(new_n483), .A2(new_n484), .B1(G136), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n460), .A2(new_n471), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  AND2_X1   g065(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n491));
  NOR2_X1   g066(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(G138), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(KEYINPUT4), .B1(new_n493), .B2(new_n471), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT72), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n458), .B2(new_n459), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n497), .B(new_n499), .C1(new_n465), .C2(new_n466), .ZN(new_n500));
  OAI211_X1 g075(.A(KEYINPUT72), .B(KEYINPUT4), .C1(new_n493), .C2(new_n471), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n496), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(G114), .A2(G2104), .ZN(new_n503));
  INV_X1    g078(.A(G126), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n471), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n476), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n505), .A2(G2105), .B1(G102), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(KEYINPUT74), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT73), .B(G651), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(G651), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n515), .A2(KEYINPUT73), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(KEYINPUT73), .ZN(new_n517));
  OAI211_X1 g092(.A(KEYINPUT74), .B(KEYINPUT6), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  AND3_X1   g093(.A1(new_n513), .A2(new_n514), .A3(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT5), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT5), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n525), .A2(KEYINPUT75), .A3(G62), .ZN(new_n528));
  NAND2_X1  g103(.A1(G75), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT75), .ZN(new_n530));
  INV_X1    g105(.A(G62), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n524), .B2(new_n531), .ZN(new_n532));
  AND3_X1   g107(.A1(new_n528), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n511), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n526), .A2(new_n527), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n513), .A2(new_n518), .A3(G543), .A4(new_n514), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n537), .A2(G50), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n535), .A2(new_n538), .ZN(G166));
  NAND3_X1  g114(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n540));
  XOR2_X1   g115(.A(new_n540), .B(KEYINPUT76), .Z(new_n541));
  INV_X1    g116(.A(G51), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n542), .B2(new_n536), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n519), .A2(new_n525), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n544), .A2(G89), .ZN(new_n545));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  XOR2_X1   g121(.A(new_n546), .B(KEYINPUT7), .Z(new_n547));
  NOR3_X1   g122(.A1(new_n543), .A2(new_n545), .A3(new_n547), .ZN(G168));
  AOI22_X1  g123(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n534), .ZN(new_n550));
  INV_X1    g125(.A(G52), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n536), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(new_n544), .B2(G90), .ZN(G171));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G56), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n524), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(new_n511), .ZN(new_n557));
  INV_X1    g132(.A(G43), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n536), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n559), .B1(new_n544), .B2(G81), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(G188));
  INV_X1    g141(.A(KEYINPUT77), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n567), .B(new_n568), .C1(new_n536), .C2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n519), .A2(G91), .A3(new_n525), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n525), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n572), .A2(new_n515), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n570), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n537), .A2(KEYINPUT77), .A3(G53), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n567), .B1(new_n536), .B2(new_n569), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n576), .A2(KEYINPUT9), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n575), .A2(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  INV_X1    g155(.A(G168), .ZN(G286));
  OR2_X1    g156(.A1(new_n535), .A2(new_n538), .ZN(G303));
  NAND2_X1  g157(.A1(new_n537), .A2(G49), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n584));
  INV_X1    g159(.A(G87), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n583), .B(new_n584), .C1(new_n585), .C2(new_n526), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT78), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G288));
  INV_X1    g163(.A(G86), .ZN(new_n589));
  INV_X1    g164(.A(G48), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n526), .A2(new_n589), .B1(new_n590), .B2(new_n536), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G61), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n524), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(new_n511), .ZN(new_n595));
  XOR2_X1   g170(.A(new_n595), .B(KEYINPUT79), .Z(new_n596));
  NOR2_X1   g171(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G305));
  AND3_X1   g173(.A1(new_n519), .A2(G85), .A3(new_n525), .ZN(new_n599));
  INV_X1    g174(.A(G47), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  OAI22_X1  g176(.A1(new_n536), .A2(new_n600), .B1(new_n601), .B2(new_n534), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n537), .A2(G54), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n524), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G651), .ZN(new_n610));
  AOI21_X1  g185(.A(KEYINPUT10), .B1(new_n544), .B2(G92), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  NOR3_X1   g188(.A1(new_n526), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n606), .B(new_n610), .C1(new_n611), .C2(new_n614), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT80), .Z(new_n616));
  OAI21_X1  g191(.A(new_n605), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n605), .B1(new_n616), .B2(G868), .ZN(G321));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(G299), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G168), .B2(new_n619), .ZN(G297));
  OAI21_X1  g196(.A(new_n620), .B1(G168), .B2(new_n619), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n616), .B1(new_n623), .B2(G860), .ZN(G148));
  NOR2_X1   g199(.A1(new_n560), .A2(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n616), .A2(new_n623), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G868), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT81), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g204(.A(new_n477), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(new_n466), .B2(new_n465), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(KEYINPUT13), .B(G2100), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n487), .A2(G123), .ZN(new_n636));
  OAI221_X1 g211(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n460), .C2(G111), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n485), .A2(G135), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n635), .A2(new_n640), .ZN(G156));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XOR2_X1   g218(.A(G2443), .B(G2446), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2427), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2430), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT15), .B(G2435), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT14), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n647), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(G14), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(G401));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2067), .B(G2678), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2072), .B(G2078), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT83), .Z(new_n662));
  XOR2_X1   g237(.A(new_n660), .B(KEYINPUT17), .Z(new_n663));
  OAI21_X1  g238(.A(new_n662), .B1(new_n658), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n659), .A2(new_n660), .A3(new_n656), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT18), .Z(new_n666));
  NAND3_X1  g241(.A1(new_n663), .A2(new_n656), .A3(new_n658), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n664), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2096), .B(G2100), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G227));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1956), .B(G2474), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT84), .ZN(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n672), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n674), .A2(new_n675), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n681), .A2(new_n678), .A3(new_n676), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n676), .A2(new_n672), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n683), .A2(new_n680), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n679), .B(new_n682), .C1(new_n684), .C2(new_n678), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1991), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1981), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1986), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n686), .B(new_n690), .ZN(G229));
  INV_X1    g266(.A(G16), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G23), .ZN(new_n693));
  INV_X1    g268(.A(new_n586), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n693), .B1(new_n694), .B2(new_n692), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT33), .ZN(new_n696));
  INV_X1    g271(.A(G1976), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n692), .A2(G6), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(new_n597), .B2(new_n692), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT32), .B(G1981), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n692), .A2(G22), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G166), .B2(new_n692), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT86), .B(G1971), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n696), .A2(new_n697), .ZN(new_n707));
  NAND4_X1  g282(.A1(new_n698), .A2(new_n702), .A3(new_n706), .A4(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n708), .A2(KEYINPUT34), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n692), .A2(G24), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(new_n603), .B2(new_n692), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(G1986), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n487), .A2(G119), .ZN(new_n714));
  OAI221_X1 g289(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n460), .C2(G107), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n485), .A2(G131), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  MUX2_X1   g292(.A(G25), .B(new_n717), .S(G29), .Z(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT35), .B(G1991), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT85), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n718), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n708), .A2(KEYINPUT34), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT87), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(KEYINPUT87), .B1(new_n708), .B2(KEYINPUT34), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n713), .B(new_n721), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT88), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT36), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT89), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G29), .B2(G33), .ZN(new_n733));
  OR3_X1    g308(.A1(new_n732), .A2(G29), .A3(G33), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT25), .Z(new_n736));
  NAND2_X1  g311(.A1(new_n485), .A2(G139), .ZN(new_n737));
  OAI21_X1  g312(.A(G127), .B1(new_n465), .B2(new_n466), .ZN(new_n738));
  NAND2_X1  g313(.A1(G115), .A2(G2104), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n736), .B(new_n737), .C1(new_n460), .C2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G29), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n733), .B(new_n734), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G2072), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT90), .Z(new_n746));
  NOR2_X1   g321(.A1(new_n743), .A2(new_n744), .ZN(new_n747));
  AND2_X1   g322(.A1(KEYINPUT24), .A2(G34), .ZN(new_n748));
  NOR2_X1   g323(.A1(KEYINPUT24), .A2(G34), .ZN(new_n749));
  NOR3_X1   g324(.A1(new_n748), .A2(new_n749), .A3(G29), .ZN(new_n750));
  INV_X1    g325(.A(G160), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(G29), .ZN(new_n752));
  INV_X1    g327(.A(G2084), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n747), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(G29), .A2(G32), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n630), .A2(G105), .B1(G129), .B2(new_n487), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n485), .A2(G141), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g334(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT91), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT26), .Z(new_n762));
  NOR2_X1   g337(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n756), .B1(new_n763), .B2(G29), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT27), .B(G1996), .Z(new_n765));
  OAI211_X1 g340(.A(new_n746), .B(new_n755), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT92), .Z(new_n767));
  AND2_X1   g342(.A1(new_n742), .A2(G26), .ZN(new_n768));
  AOI22_X1  g343(.A1(G128), .A2(new_n487), .B1(new_n485), .B2(G140), .ZN(new_n769));
  OAI221_X1 g344(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n460), .C2(G116), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n768), .B1(new_n771), .B2(G29), .ZN(new_n772));
  MUX2_X1   g347(.A(new_n768), .B(new_n772), .S(KEYINPUT28), .Z(new_n773));
  INV_X1    g348(.A(G2067), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n764), .A2(new_n765), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n639), .A2(new_n742), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT93), .ZN(new_n778));
  INV_X1    g353(.A(G28), .ZN(new_n779));
  NOR3_X1   g354(.A1(new_n779), .A2(KEYINPUT94), .A3(KEYINPUT30), .ZN(new_n780));
  OAI21_X1  g355(.A(KEYINPUT94), .B1(new_n779), .B2(KEYINPUT30), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(new_n742), .ZN(new_n782));
  AOI211_X1 g357(.A(new_n780), .B(new_n782), .C1(KEYINPUT30), .C2(new_n779), .ZN(new_n783));
  NOR4_X1   g358(.A1(new_n775), .A2(new_n776), .A3(new_n778), .A4(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(KEYINPUT95), .B1(G5), .B2(G16), .ZN(new_n785));
  OR3_X1    g360(.A1(KEYINPUT95), .A2(G5), .A3(G16), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n785), .B(new_n786), .C1(G301), .C2(new_n692), .ZN(new_n787));
  INV_X1    g362(.A(G1961), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n742), .A2(G35), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G162), .B2(new_n742), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT29), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(G2090), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n784), .A2(new_n789), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n692), .A2(G21), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G168), .B2(new_n692), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G1966), .ZN(new_n797));
  NOR2_X1   g372(.A1(G27), .A2(G29), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G164), .B2(G29), .ZN(new_n799));
  INV_X1    g374(.A(G2078), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n792), .B2(G2090), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n794), .A2(new_n797), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n692), .A2(G19), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n560), .B2(new_n692), .ZN(new_n805));
  OAI22_X1  g380(.A1(new_n787), .A2(new_n788), .B1(new_n805), .B2(G1341), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n752), .A2(new_n753), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT96), .Z(new_n808));
  AOI211_X1 g383(.A(new_n806), .B(new_n808), .C1(G1341), .C2(new_n805), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n767), .A2(new_n803), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n692), .A2(G20), .ZN(new_n811));
  AND3_X1   g386(.A1(new_n576), .A2(KEYINPUT9), .A3(new_n577), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n812), .A2(new_n574), .ZN(new_n813));
  OAI211_X1 g388(.A(KEYINPUT23), .B(new_n811), .C1(new_n813), .C2(new_n692), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(KEYINPUT23), .B2(new_n811), .ZN(new_n815));
  INV_X1    g390(.A(G1956), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(G4), .A2(G16), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(new_n616), .B2(G16), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(G1348), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n810), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT31), .B(G11), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n727), .A2(new_n728), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n726), .A2(new_n730), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n731), .A2(new_n821), .A3(new_n822), .A4(new_n824), .ZN(G150));
  INV_X1    g400(.A(G150), .ZN(G311));
  NAND2_X1  g401(.A1(new_n616), .A2(G559), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT38), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT97), .B(G93), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n526), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(G55), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n525), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n832));
  OAI22_X1  g407(.A1(new_n536), .A2(new_n831), .B1(new_n832), .B2(new_n534), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(G81), .ZN(new_n835));
  OAI221_X1 g410(.A(new_n557), .B1(new_n558), .B2(new_n536), .C1(new_n526), .C2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n834), .A2(new_n836), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n828), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(KEYINPUT39), .ZN(new_n843));
  AOI21_X1  g418(.A(G860), .B1(new_n843), .B2(KEYINPUT98), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n842), .A2(KEYINPUT39), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n844), .B(new_n845), .C1(KEYINPUT98), .C2(new_n843), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n830), .A2(new_n833), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(G860), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(KEYINPUT37), .Z(new_n849));
  NAND2_X1  g424(.A1(new_n846), .A2(new_n849), .ZN(G145));
  XNOR2_X1  g425(.A(new_n489), .B(new_n751), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n508), .B(new_n771), .ZN(new_n853));
  AOI22_X1  g428(.A1(G130), .A2(new_n487), .B1(new_n485), .B2(G142), .ZN(new_n854));
  OAI221_X1 g429(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n460), .C2(G118), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT99), .Z(new_n857));
  XNOR2_X1  g432(.A(new_n853), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n741), .B(new_n717), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n860), .A2(new_n763), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n633), .B(new_n639), .Z(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n763), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n862), .B1(new_n861), .B2(new_n863), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n852), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n866), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n868), .A2(new_n851), .A3(new_n864), .ZN(new_n869));
  INV_X1    g444(.A(G37), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n867), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g447(.A(new_n626), .B(new_n840), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n544), .A2(KEYINPUT10), .A3(G92), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n612), .B1(new_n526), .B2(new_n613), .ZN(new_n875));
  AOI22_X1  g450(.A1(new_n874), .A2(new_n875), .B1(G651), .B2(new_n609), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n813), .A2(new_n876), .A3(new_n606), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n615), .A2(G299), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(KEYINPUT100), .B(KEYINPUT41), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT41), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n877), .A2(new_n878), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n880), .B1(new_n873), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT42), .ZN(new_n887));
  OR3_X1    g462(.A1(new_n599), .A2(KEYINPUT101), .A3(new_n602), .ZN(new_n888));
  OAI21_X1  g463(.A(KEYINPUT101), .B1(new_n599), .B2(new_n602), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n888), .A2(new_n586), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n586), .B1(new_n888), .B2(new_n889), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(G305), .A2(G166), .ZN(new_n893));
  NAND2_X1  g468(.A1(G303), .A2(new_n597), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n893), .A2(new_n894), .A3(KEYINPUT102), .ZN(new_n895));
  AOI21_X1  g470(.A(KEYINPUT102), .B1(new_n893), .B2(new_n894), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n892), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n893), .A2(new_n894), .ZN(new_n898));
  OAI22_X1  g473(.A1(new_n898), .A2(KEYINPUT102), .B1(new_n891), .B2(new_n890), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT42), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n880), .B(new_n901), .C1(new_n873), .C2(new_n885), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n887), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n900), .B1(new_n887), .B2(new_n902), .ZN(new_n904));
  OAI21_X1  g479(.A(G868), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n847), .A2(new_n619), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(G295));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n906), .ZN(G331));
  NAND2_X1  g483(.A1(new_n847), .A2(new_n560), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n909), .A2(G301), .A3(new_n837), .ZN(new_n910));
  AOI21_X1  g485(.A(G301), .B1(new_n909), .B2(new_n837), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n910), .A2(new_n911), .A3(G286), .ZN(new_n912));
  OAI21_X1  g487(.A(G171), .B1(new_n838), .B2(new_n839), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n909), .A2(G301), .A3(new_n837), .ZN(new_n914));
  AOI21_X1  g489(.A(G168), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n884), .ZN(new_n916));
  INV_X1    g491(.A(new_n881), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n917), .B1(new_n877), .B2(new_n878), .ZN(new_n918));
  OAI22_X1  g493(.A1(new_n912), .A2(new_n915), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n897), .A2(new_n899), .ZN(new_n920));
  OAI21_X1  g495(.A(G286), .B1(new_n910), .B2(new_n911), .ZN(new_n921));
  INV_X1    g496(.A(new_n879), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n913), .A2(G168), .A3(new_n914), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n919), .A2(new_n920), .A3(new_n924), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n925), .A2(new_n870), .ZN(new_n926));
  INV_X1    g501(.A(new_n924), .ZN(new_n927));
  AOI22_X1  g502(.A1(new_n921), .A2(new_n923), .B1(new_n882), .B2(new_n884), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n900), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n924), .B(KEYINPUT103), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n879), .A2(new_n917), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n933), .B1(new_n883), .B2(new_n879), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n921), .A2(new_n923), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n926), .B1(new_n936), .B2(new_n920), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n931), .B1(new_n937), .B2(KEYINPUT43), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT104), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n926), .A2(new_n941), .A3(new_n942), .A4(new_n929), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n929), .A2(new_n942), .A3(new_n870), .A4(new_n925), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT104), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n939), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT105), .ZN(new_n947));
  XOR2_X1   g522(.A(new_n924), .B(KEYINPUT103), .Z(new_n948));
  NAND2_X1  g523(.A1(new_n934), .A2(new_n935), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n920), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n926), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT43), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n946), .A2(new_n947), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n947), .B1(new_n946), .B2(new_n952), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n940), .B1(new_n953), .B2(new_n954), .ZN(G397));
  XOR2_X1   g530(.A(KEYINPUT106), .B(G1384), .Z(new_n956));
  NAND2_X1  g531(.A1(new_n508), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT107), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n957), .B(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT45), .ZN(new_n960));
  INV_X1    g535(.A(G40), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n470), .A2(new_n479), .A3(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n959), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n963), .B(KEYINPUT108), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n771), .B(new_n774), .ZN(new_n965));
  INV_X1    g540(.A(G1996), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n965), .B1(new_n966), .B2(new_n763), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n717), .B(new_n719), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n969), .B(KEYINPUT109), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n964), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n963), .A2(G1996), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n763), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n968), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  OR2_X1    g549(.A1(G290), .A2(G1986), .ZN(new_n975));
  NAND2_X1  g550(.A1(G290), .A2(G1986), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n963), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G1966), .ZN(new_n979));
  AOI21_X1  g554(.A(G1384), .B1(new_n502), .B2(new_n507), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n962), .B1(new_n980), .B2(KEYINPUT45), .ZN(new_n981));
  AOI211_X1 g556(.A(new_n960), .B(G1384), .C1(new_n502), .C2(new_n507), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G1384), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n508), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT50), .ZN(new_n986));
  XNOR2_X1  g561(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n980), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n986), .A2(new_n753), .A3(new_n962), .A4(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n983), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT119), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT119), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n983), .A2(new_n990), .A3(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n992), .A2(G168), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(G8), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT51), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n983), .A2(new_n990), .A3(new_n993), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n993), .B1(new_n983), .B2(new_n990), .ZN(new_n999));
  OAI211_X1 g574(.A(G8), .B(G286), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n983), .A2(new_n990), .A3(G168), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(new_n1002), .A3(G8), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT120), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n997), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1002), .B1(new_n995), .B2(G8), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT120), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g585(.A(KEYINPUT121), .B(KEYINPUT54), .Z(new_n1011));
  NAND3_X1  g586(.A1(new_n986), .A2(new_n962), .A3(new_n989), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(new_n788), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT122), .ZN(new_n1014));
  INV_X1    g589(.A(new_n981), .ZN(new_n1015));
  INV_X1    g590(.A(new_n982), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1015), .A2(KEYINPUT53), .A3(new_n800), .A4(new_n1016), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n1013), .A2(new_n1014), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1014), .B1(new_n1013), .B2(new_n1017), .ZN(new_n1019));
  OR2_X1    g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT123), .ZN(new_n1022));
  OR2_X1    g597(.A1(new_n1021), .A2(KEYINPUT123), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n508), .A2(KEYINPUT45), .A3(new_n956), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1024), .B(new_n962), .C1(KEYINPUT45), .C2(new_n980), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1022), .B(new_n1023), .C1(new_n1025), .C2(G2078), .ZN(new_n1026));
  AOI21_X1  g601(.A(G301), .B1(new_n1020), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n959), .A2(new_n960), .ZN(new_n1028));
  INV_X1    g603(.A(new_n470), .ZN(new_n1029));
  INV_X1    g604(.A(new_n479), .ZN(new_n1030));
  OAI21_X1  g605(.A(G40), .B1(new_n1030), .B2(KEYINPUT124), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1031), .B1(KEYINPUT124), .B2(new_n1030), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1028), .A2(new_n1029), .A3(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1024), .A2(KEYINPUT53), .A3(new_n800), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1026), .B(new_n1013), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1035), .A2(G171), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1011), .B1(new_n1027), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(G305), .A2(G1981), .ZN(new_n1038));
  INV_X1    g613(.A(G1981), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n597), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT49), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n980), .A2(new_n962), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1038), .A2(KEYINPUT49), .A3(new_n1040), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1043), .A2(G8), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(G8), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1047), .B1(G1976), .B2(new_n694), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n1049));
  OR2_X1    g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1048), .B(new_n1049), .C1(new_n587), .C2(G1976), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n1046), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G8), .ZN(new_n1053));
  NOR2_X1   g628(.A1(G166), .A2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1054), .B(KEYINPUT55), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT112), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n1058));
  AND4_X1   g633(.A1(new_n1057), .A2(new_n508), .A3(new_n1058), .A4(new_n984), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n962), .B1(new_n980), .B2(new_n988), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1057), .B1(new_n980), .B2(new_n1058), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT111), .B(G2090), .Z(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G1971), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n1062), .A2(new_n1064), .B1(new_n1065), .B2(new_n1025), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1056), .B1(new_n1066), .B2(new_n1053), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n1012), .A2(new_n1063), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1025), .A2(new_n1065), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1053), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n1055), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1052), .A2(new_n1067), .A3(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1020), .A2(G301), .A3(new_n1026), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1035), .A2(G171), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1073), .A2(KEYINPUT54), .A3(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1010), .A2(new_n1037), .A3(new_n1072), .A4(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT56), .B(G2072), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1015), .A2(new_n1024), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1079), .B1(new_n812), .B2(new_n574), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n575), .A2(KEYINPUT57), .A3(new_n578), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1078), .B(new_n1082), .C1(new_n1062), .C2(G1956), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1082), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1029), .A2(G40), .A3(new_n1030), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1088), .B1(new_n985), .B2(new_n987), .ZN(new_n1089));
  AOI21_X1  g664(.A(G1956), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1077), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1025), .A2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1086), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n508), .A2(new_n1058), .A3(new_n984), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT112), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n980), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n816), .B1(new_n1097), .B2(new_n1060), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1098), .A2(KEYINPUT113), .A3(new_n1082), .A4(new_n1078), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1085), .A2(new_n1093), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT61), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT114), .B1(new_n1025), .B2(G1996), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT114), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1015), .A2(new_n1103), .A3(new_n966), .A4(new_n1024), .ZN(new_n1104));
  XOR2_X1   g679(.A(KEYINPUT58), .B(G1341), .Z(new_n1105));
  NAND2_X1  g680(.A1(new_n1044), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1102), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n560), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1109), .A2(KEYINPUT115), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1107), .B(new_n560), .C1(KEYINPUT115), .C2(new_n1109), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1100), .A2(new_n1101), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1101), .B1(new_n1083), .B2(KEYINPUT116), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT116), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1098), .A2(new_n1115), .A3(new_n1082), .A4(new_n1078), .ZN(new_n1116));
  AND4_X1   g691(.A1(KEYINPUT117), .A2(new_n1114), .A3(new_n1093), .A4(new_n1116), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1093), .A2(new_n1116), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT117), .B1(new_n1118), .B2(new_n1114), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1113), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT118), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(G1348), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1044), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1012), .A2(new_n1123), .B1(new_n774), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT60), .ZN(new_n1126));
  XOR2_X1   g701(.A(new_n1126), .B(new_n615), .Z(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(KEYINPUT60), .B2(new_n1125), .ZN(new_n1128));
  OAI211_X1 g703(.A(KEYINPUT118), .B(new_n1113), .C1(new_n1117), .C2(new_n1119), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1122), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1093), .B1(new_n615), .B2(new_n1125), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1131), .A2(new_n1085), .A3(new_n1099), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1076), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1005), .B1(new_n997), .B2(new_n1004), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1007), .A2(new_n1008), .A3(KEYINPUT120), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT62), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT62), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1006), .A2(new_n1009), .A3(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1136), .A2(new_n1072), .A3(new_n1027), .A4(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1052), .A2(new_n1055), .A3(new_n1070), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1141), .A2(new_n697), .A3(new_n587), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1047), .B1(new_n1142), .B2(new_n1040), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n991), .A2(G8), .A3(G168), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1052), .A2(new_n1067), .A3(new_n1071), .A4(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT63), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1070), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1146), .B1(new_n1148), .B2(new_n1056), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1052), .A2(new_n1149), .A3(new_n1071), .A4(new_n1144), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1143), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1139), .A2(new_n1140), .A3(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n978), .B1(new_n1133), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n968), .A2(new_n973), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1154), .A2(new_n717), .A3(new_n719), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n771), .A2(G2067), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n964), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n974), .A2(KEYINPUT126), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n974), .A2(KEYINPUT126), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT48), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1160), .B1(new_n963), .B2(new_n975), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1158), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n963), .A2(new_n1160), .A3(new_n975), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1157), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  XOR2_X1   g739(.A(new_n972), .B(KEYINPUT46), .Z(new_n1165));
  NAND2_X1  g740(.A1(new_n965), .A2(new_n763), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n964), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n1168), .A2(KEYINPUT125), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(KEYINPUT125), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(KEYINPUT47), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT47), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1169), .A2(new_n1173), .A3(new_n1170), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1164), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1153), .A2(new_n1175), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g751(.A1(new_n654), .A2(new_n670), .A3(G319), .ZN(new_n1178));
  INV_X1    g752(.A(KEYINPUT127), .ZN(new_n1179));
  AND2_X1   g753(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1181));
  NOR3_X1   g755(.A1(new_n1180), .A2(new_n1181), .A3(G229), .ZN(new_n1182));
  NAND3_X1  g756(.A1(new_n938), .A2(new_n871), .A3(new_n1182), .ZN(G225));
  INV_X1    g757(.A(G225), .ZN(G308));
endmodule


