//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 1 1 0 1 0 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n509, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n545,
    new_n546, new_n547, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n591, new_n592, new_n593, new_n594, new_n597,
    new_n599, new_n600, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1203, new_n1204, new_n1205, new_n1206;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(G125), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI211_X1 g038(.A(G137), .B(new_n458), .C1(new_n459), .C2(new_n460), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n463), .A2(new_n468), .ZN(G160));
  NOR2_X1   g044(.A1(new_n459), .A2(new_n460), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G136), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n470), .A2(new_n458), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G124), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n458), .A2(G112), .ZN(new_n475));
  OAI21_X1  g050(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n472), .B(new_n474), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT65), .ZN(G162));
  NAND2_X1  g053(.A1(KEYINPUT4), .A2(G138), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(new_n465), .ZN(new_n481));
  NAND2_X1  g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n479), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AND2_X1   g058(.A1(G102), .A2(G2104), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n458), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G126), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n486), .B1(new_n481), .B2(new_n482), .ZN(new_n487));
  AND2_X1   g062(.A1(G114), .A2(G2104), .ZN(new_n488));
  OAI21_X1  g063(.A(G2105), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI211_X1 g064(.A(G138), .B(new_n458), .C1(new_n459), .C2(new_n460), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n485), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G164));
  INV_X1    g069(.A(G50), .ZN(new_n495));
  AND2_X1   g070(.A1(KEYINPUT6), .A2(G651), .ZN(new_n496));
  NOR2_X1   g071(.A1(KEYINPUT6), .A2(G651), .ZN(new_n497));
  OR2_X1    g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G543), .ZN(new_n499));
  XNOR2_X1  g074(.A(KEYINPUT5), .B(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G88), .ZN(new_n502));
  OAI22_X1  g077(.A1(new_n495), .A2(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n500), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OR2_X1    g081(.A1(new_n503), .A2(new_n506), .ZN(G303));
  INV_X1    g082(.A(G303), .ZN(G166));
  NAND3_X1  g083(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n509));
  XNOR2_X1  g084(.A(new_n509), .B(KEYINPUT7), .ZN(new_n510));
  INV_X1    g085(.A(G51), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n499), .B2(new_n511), .ZN(new_n512));
  XOR2_X1   g087(.A(KEYINPUT5), .B(G543), .Z(new_n513));
  NAND2_X1  g088(.A1(new_n498), .A2(G89), .ZN(new_n514));
  NAND2_X1  g089(.A1(G63), .A2(G651), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n512), .A2(new_n516), .ZN(G168));
  NAND2_X1  g092(.A1(G77), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G64), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n513), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT66), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n505), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n522), .B1(new_n521), .B2(new_n520), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n496), .A2(new_n497), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n513), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n525), .A2(G90), .B1(new_n527), .B2(G52), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n523), .A2(new_n528), .ZN(G301));
  INV_X1    g104(.A(G301), .ZN(G171));
  INV_X1    g105(.A(G43), .ZN(new_n531));
  INV_X1    g106(.A(G81), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n531), .A2(new_n499), .B1(new_n501), .B2(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n500), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n505), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(KEYINPUT67), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n527), .A2(G43), .ZN(new_n538));
  OAI221_X1 g113(.A(new_n538), .B1(new_n501), .B2(new_n532), .C1(new_n505), .C2(new_n534), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT67), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  NAND4_X1  g118(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT68), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g122(.A1(G319), .A2(G483), .A3(G661), .A4(new_n547), .ZN(G188));
  AOI22_X1  g123(.A1(new_n500), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G91), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n505), .A2(new_n549), .B1(new_n501), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  OAI211_X1 g127(.A(G53), .B(G543), .C1(new_n496), .C2(new_n497), .ZN(new_n553));
  NAND2_X1  g128(.A1(KEYINPUT69), .A2(KEYINPUT9), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(KEYINPUT69), .A2(KEYINPUT9), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n553), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n552), .A2(new_n559), .ZN(G299));
  INV_X1    g135(.A(G168), .ZN(G286));
  NAND2_X1  g136(.A1(new_n525), .A2(G87), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n500), .B2(G74), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n527), .A2(G49), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(G288));
  NAND2_X1  g140(.A1(new_n525), .A2(G86), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n527), .A2(G48), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n500), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n569), .A2(new_n505), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G305));
  AOI22_X1  g147(.A1(new_n525), .A2(G85), .B1(new_n527), .B2(G47), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n500), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n505), .B2(new_n574), .ZN(G290));
  NAND2_X1  g150(.A1(G301), .A2(G868), .ZN(new_n576));
  NAND2_X1  g151(.A1(G79), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G66), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n513), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G651), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT70), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n527), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g158(.A(G54), .B1(new_n527), .B2(new_n581), .ZN(new_n584));
  AND3_X1   g159(.A1(new_n525), .A2(KEYINPUT10), .A3(G92), .ZN(new_n585));
  AOI21_X1  g160(.A(KEYINPUT10), .B1(new_n525), .B2(G92), .ZN(new_n586));
  OAI221_X1 g161(.A(new_n580), .B1(new_n583), .B2(new_n584), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n576), .B1(new_n588), .B2(G868), .ZN(G284));
  OAI21_X1  g164(.A(new_n576), .B1(new_n588), .B2(G868), .ZN(G321));
  INV_X1    g165(.A(KEYINPUT71), .ZN(new_n591));
  INV_X1    g166(.A(G868), .ZN(new_n592));
  NOR2_X1   g167(.A1(G168), .A2(new_n592), .ZN(new_n593));
  AOI211_X1 g168(.A(new_n591), .B(new_n593), .C1(new_n592), .C2(G299), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n594), .B1(new_n591), .B2(new_n593), .ZN(G280));
  XNOR2_X1  g170(.A(G280), .B(KEYINPUT72), .ZN(G297));
  INV_X1    g171(.A(G559), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n588), .B1(new_n597), .B2(G860), .ZN(G148));
  NAND2_X1  g173(.A1(new_n588), .A2(new_n597), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(G868), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(G868), .B2(new_n542), .ZN(G323));
  XNOR2_X1  g176(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g177(.A1(new_n481), .A2(new_n482), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(new_n466), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT12), .Z(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT13), .Z(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(G2100), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n471), .A2(G135), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n473), .A2(G123), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n458), .A2(G111), .ZN(new_n610));
  OAI21_X1  g185(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n611));
  OAI211_X1 g186(.A(new_n608), .B(new_n609), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT73), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(G2096), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n607), .A2(new_n614), .ZN(G156));
  XOR2_X1   g190(.A(KEYINPUT15), .B(G2435), .Z(new_n616));
  XOR2_X1   g191(.A(KEYINPUT74), .B(G2438), .Z(new_n617));
  XOR2_X1   g192(.A(new_n616), .B(new_n617), .Z(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(G2427), .B(G2430), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(KEYINPUT14), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT75), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n619), .A2(new_n621), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(G2443), .B(G2446), .Z(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G1341), .B(G1348), .Z(new_n628));
  INV_X1    g203(.A(new_n626), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n623), .A2(new_n624), .A3(new_n629), .ZN(new_n630));
  AND3_X1   g205(.A1(new_n627), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n628), .B1(new_n627), .B2(new_n630), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(G14), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(new_n633), .B2(new_n635), .ZN(new_n638));
  AND2_X1   g213(.A1(new_n636), .A2(new_n638), .ZN(G401));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  XNOR2_X1  g215(.A(G2067), .B(G2678), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT18), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(KEYINPUT17), .ZN(new_n646));
  INV_X1    g221(.A(new_n640), .ZN(new_n647));
  INV_X1    g222(.A(new_n641), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n647), .A2(new_n643), .A3(new_n648), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(new_n642), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n645), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2096), .B(G2100), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(G227));
  XNOR2_X1  g229(.A(G1971), .B(G1976), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT19), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G1956), .B(G2474), .Z(new_n658));
  XOR2_X1   g233(.A(G1961), .B(G1966), .Z(new_n659));
  AND2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT20), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n658), .A2(new_n659), .ZN(new_n663));
  NOR3_X1   g238(.A1(new_n657), .A2(new_n660), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n657), .B2(new_n663), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G1991), .B(G1996), .Z(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1981), .B(G1986), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n668), .A2(new_n670), .ZN(new_n673));
  AND3_X1   g248(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n672), .B1(new_n671), .B2(new_n673), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(G229));
  NOR2_X1   g251(.A1(G29), .A2(G35), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(G162), .B2(G29), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT29), .Z(new_n679));
  INV_X1    g254(.A(G2090), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT93), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n679), .A2(new_n680), .ZN(new_n683));
  INV_X1    g258(.A(G16), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G19), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(new_n542), .B2(new_n684), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT85), .B(G1341), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n684), .A2(G20), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT23), .ZN(new_n690));
  INV_X1    g265(.A(G299), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(new_n684), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT94), .B(G1956), .Z(new_n694));
  OR2_X1    g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g270(.A(KEYINPUT86), .B1(G104), .B2(G2105), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NOR3_X1   g272(.A1(KEYINPUT86), .A2(G104), .A3(G2105), .ZN(new_n698));
  OAI221_X1 g273(.A(G2104), .B1(G116), .B2(new_n458), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n603), .A2(G140), .A3(new_n458), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n603), .A2(G128), .A3(G2105), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G29), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n704));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G26), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n704), .B(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G2067), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n693), .A2(new_n694), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n695), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n684), .A2(G4), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(new_n588), .B2(new_n684), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G1348), .ZN(new_n715));
  NOR4_X1   g290(.A1(new_n683), .A2(new_n688), .A3(new_n712), .A4(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n682), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(G27), .A2(G29), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G164), .B2(G29), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n719), .A2(G2078), .ZN(new_n720));
  NAND2_X1  g295(.A1(G115), .A2(G2104), .ZN(new_n721));
  INV_X1    g296(.A(G127), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n470), .B2(new_n722), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n723), .A2(G2105), .B1(new_n471), .B2(G139), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n725), .A2(KEYINPUT88), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(KEYINPUT88), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n726), .A2(KEYINPUT25), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT25), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AND3_X1   g306(.A1(new_n724), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n732), .A2(new_n705), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n705), .B2(G33), .ZN(new_n734));
  INV_X1    g309(.A(G2072), .ZN(new_n735));
  OAI22_X1  g310(.A1(new_n734), .A2(new_n735), .B1(new_n719), .B2(G2078), .ZN(new_n736));
  AOI211_X1 g311(.A(new_n720), .B(new_n736), .C1(new_n735), .C2(new_n734), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n705), .A2(G32), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n471), .A2(G141), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n466), .A2(G105), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n603), .A2(G129), .A3(G2105), .ZN(new_n741));
  NAND3_X1  g316(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT26), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n739), .A2(new_n740), .A3(new_n741), .A4(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n738), .B1(new_n746), .B2(new_n705), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT27), .B(G1996), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n684), .A2(G21), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G168), .B2(new_n684), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G1966), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT31), .B(G11), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT30), .B(G28), .Z(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(new_n754), .B2(G29), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n612), .A2(new_n705), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT90), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n757), .B2(new_n756), .ZN(new_n759));
  NAND2_X1  g334(.A1(G160), .A2(G29), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G34), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n760), .B1(G29), .B2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G2084), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NOR4_X1   g340(.A1(new_n749), .A2(new_n752), .A3(new_n759), .A4(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(G5), .A2(G16), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT91), .Z(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G301), .B2(new_n684), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1961), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n737), .A2(new_n766), .A3(new_n770), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n771), .A2(KEYINPUT92), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(KEYINPUT92), .ZN(new_n773));
  NOR3_X1   g348(.A1(new_n717), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  OR2_X1    g349(.A1(G288), .A2(KEYINPUT80), .ZN(new_n775));
  NAND2_X1  g350(.A1(G288), .A2(KEYINPUT80), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(G16), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n684), .A2(G23), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT33), .B(G1976), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT81), .Z(new_n783));
  AND2_X1   g358(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n781), .A2(new_n783), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(G303), .A2(G16), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n684), .A2(G22), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(KEYINPUT82), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT82), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n787), .A2(new_n791), .A3(new_n788), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(G1971), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n790), .A2(G1971), .A3(new_n792), .ZN(new_n796));
  NOR2_X1   g371(.A1(G6), .A2(G16), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n571), .B2(G16), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT32), .B(G1981), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n795), .A2(new_n796), .A3(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n786), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(KEYINPUT84), .B1(new_n802), .B2(KEYINPUT34), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT83), .ZN(new_n805));
  MUX2_X1   g380(.A(G24), .B(G290), .S(G16), .Z(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT79), .Z(new_n807));
  INV_X1    g382(.A(G1986), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n705), .A2(G25), .ZN(new_n812));
  OAI21_X1  g387(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n813));
  INV_X1    g388(.A(G107), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(G2105), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n473), .B2(G119), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n603), .A2(G131), .A3(new_n458), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n817), .A2(KEYINPUT76), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n817), .A2(KEYINPUT76), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n816), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT77), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n812), .B1(new_n822), .B2(new_n705), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT35), .B(G1991), .Z(new_n824));
  OR2_X1    g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n825), .A2(KEYINPUT78), .A3(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT78), .ZN(new_n828));
  INV_X1    g403(.A(new_n826), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n823), .A2(new_n824), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n811), .A2(new_n827), .A3(new_n831), .ZN(new_n832));
  NOR3_X1   g407(.A1(new_n786), .A2(new_n801), .A3(KEYINPUT34), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n805), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(KEYINPUT78), .B1(new_n825), .B2(new_n826), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(new_n809), .B2(new_n810), .ZN(new_n836));
  OR3_X1    g411(.A1(new_n786), .A2(new_n801), .A3(KEYINPUT34), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n836), .A2(new_n837), .A3(KEYINPUT83), .A4(new_n827), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n804), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n774), .B1(new_n839), .B2(KEYINPUT36), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT36), .ZN(new_n841));
  AOI211_X1 g416(.A(new_n841), .B(new_n804), .C1(new_n838), .C2(new_n834), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n840), .A2(new_n842), .ZN(G311));
  AND2_X1   g418(.A1(new_n834), .A2(new_n838), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n841), .B1(new_n844), .B2(new_n804), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n839), .A2(KEYINPUT36), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n845), .A2(new_n846), .A3(new_n774), .ZN(G150));
  INV_X1    g422(.A(G55), .ZN(new_n848));
  INV_X1    g423(.A(G93), .ZN(new_n849));
  OAI22_X1  g424(.A1(new_n848), .A2(new_n499), .B1(new_n501), .B2(new_n849), .ZN(new_n850));
  AOI22_X1  g425(.A1(new_n500), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n851), .A2(new_n505), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(G860), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT37), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n536), .A2(KEYINPUT67), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n539), .A2(new_n540), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n853), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n853), .A2(new_n536), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT38), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n588), .A2(G559), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n865), .A2(KEYINPUT39), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n866), .A2(KEYINPUT96), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(KEYINPUT96), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n867), .A2(new_n854), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n865), .A2(KEYINPUT39), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT95), .Z(new_n871));
  OAI21_X1  g446(.A(new_n856), .B1(new_n869), .B2(new_n871), .ZN(G145));
  XNOR2_X1  g447(.A(new_n612), .B(G160), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(G162), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n493), .B(KEYINPUT97), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n745), .A2(new_n702), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n700), .A2(new_n701), .ZN(new_n877));
  AOI22_X1  g452(.A1(new_n471), .A2(G141), .B1(G105), .B2(new_n466), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n741), .A2(new_n744), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .A4(new_n699), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n724), .A2(new_n728), .A3(new_n731), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n876), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n881), .B1(new_n876), .B2(new_n880), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n875), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n876), .A2(new_n880), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n732), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n493), .B(KEYINPUT97), .Z(new_n887));
  NAND3_X1  g462(.A1(new_n876), .A2(new_n880), .A3(new_n881), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n473), .A2(G130), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n471), .A2(G142), .ZN(new_n892));
  OR3_X1    g467(.A1(new_n458), .A2(KEYINPUT98), .A3(G118), .ZN(new_n893));
  OAI21_X1  g468(.A(KEYINPUT98), .B1(new_n458), .B2(G118), .ZN(new_n894));
  OR2_X1    g469(.A1(G106), .A2(G2105), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n893), .A2(G2104), .A3(new_n894), .A4(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n891), .A2(new_n892), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT99), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n820), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n817), .B(KEYINPUT76), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n900), .A2(KEYINPUT99), .A3(new_n816), .ZN(new_n901));
  INV_X1    g476(.A(new_n605), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n902), .B1(new_n899), .B2(new_n901), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n897), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n905), .ZN(new_n907));
  INV_X1    g482(.A(new_n897), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(new_n908), .A3(new_n903), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n890), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT100), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT101), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n890), .A2(new_n906), .A3(new_n909), .A4(KEYINPUT100), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n906), .A2(new_n909), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n916), .A2(new_n889), .A3(new_n884), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n913), .B1(new_n912), .B2(new_n914), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n874), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT103), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n922));
  AOI22_X1  g497(.A1(new_n890), .A2(new_n922), .B1(new_n906), .B2(new_n909), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n884), .A2(new_n889), .A3(KEYINPUT102), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n874), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n912), .A2(new_n914), .ZN(new_n926));
  AOI21_X1  g501(.A(G37), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n920), .A2(new_n921), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n921), .B1(new_n920), .B2(new_n927), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT40), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n920), .A2(new_n927), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT103), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT40), .B1(new_n934), .B2(new_n928), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n932), .A2(new_n935), .ZN(G395));
  XNOR2_X1  g511(.A(G303), .B(G290), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n777), .A2(new_n571), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n777), .A2(new_n571), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n938), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n941), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n943), .A2(new_n937), .A3(new_n939), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT105), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT42), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n862), .B(new_n599), .ZN(new_n949));
  NAND2_X1  g524(.A1(G299), .A2(KEYINPUT104), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT104), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n552), .A2(new_n951), .A3(new_n559), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n588), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n587), .A2(KEYINPUT104), .A3(G299), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT41), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n953), .A2(new_n954), .A3(KEYINPUT41), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n949), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n955), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n960), .B1(new_n949), .B2(new_n961), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n948), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n948), .A2(new_n962), .ZN(new_n964));
  OAI21_X1  g539(.A(G868), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(G868), .B2(new_n853), .ZN(G295));
  OAI21_X1  g541(.A(new_n965), .B1(G868), .B2(new_n853), .ZN(G331));
  INV_X1    g542(.A(new_n853), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(new_n537), .B2(new_n541), .ZN(new_n969));
  AOI21_X1  g544(.A(G168), .B1(new_n523), .B2(new_n528), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n523), .A2(G168), .A3(new_n528), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n969), .A2(new_n860), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n972), .ZN(new_n974));
  OAI22_X1  g549(.A1(new_n859), .A2(new_n861), .B1(new_n974), .B2(new_n970), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT107), .B1(new_n976), .B2(new_n955), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n961), .A2(new_n978), .A3(new_n975), .A4(new_n973), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT106), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n973), .A2(new_n975), .A3(new_n981), .ZN(new_n982));
  OAI221_X1 g557(.A(KEYINPUT106), .B1(new_n974), .B2(new_n970), .C1(new_n859), .C2(new_n861), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n982), .A2(new_n957), .A3(new_n958), .A4(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n945), .B1(new_n980), .B2(new_n984), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n984), .A2(new_n977), .A3(new_n945), .A4(new_n979), .ZN(new_n986));
  INV_X1    g561(.A(G37), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OR3_X1    g563(.A1(new_n985), .A2(new_n988), .A3(KEYINPUT43), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT43), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n976), .A2(new_n957), .A3(new_n958), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n982), .A2(new_n983), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n991), .B1(new_n992), .B2(new_n955), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n988), .B1(new_n993), .B2(new_n946), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n989), .B(KEYINPUT44), .C1(new_n990), .C2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT43), .B1(new_n985), .B2(new_n988), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n993), .A2(new_n946), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n997), .A2(new_n990), .A3(new_n987), .A4(new_n986), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT108), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT108), .ZN(new_n1002));
  AOI211_X1 g577(.A(new_n1002), .B(KEYINPUT44), .C1(new_n996), .C2(new_n998), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n995), .B1(new_n1001), .B2(new_n1003), .ZN(G397));
  INV_X1    g579(.A(G1384), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n493), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT45), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(new_n1007), .B2(new_n1006), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n461), .A2(new_n462), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(G2105), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1011), .A2(G40), .A3(new_n467), .A4(new_n464), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(G290), .A2(G1986), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n1015), .A2(KEYINPUT48), .ZN(new_n1016));
  INV_X1    g591(.A(G1996), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n745), .B(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n702), .B(new_n709), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g595(.A(new_n820), .B(new_n824), .Z(new_n1021));
  OAI21_X1  g596(.A(new_n1013), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1015), .A2(KEYINPUT48), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1016), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n822), .A2(new_n824), .ZN(new_n1025));
  OAI22_X1  g600(.A1(new_n1025), .A2(new_n1020), .B1(G2067), .B2(new_n702), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(new_n1013), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1013), .A2(new_n1017), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT46), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1019), .A2(new_n746), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n1028), .A2(new_n1029), .B1(new_n1013), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(new_n1029), .B2(new_n1028), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT47), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1024), .B(new_n1027), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1034), .B1(new_n1033), .B2(new_n1032), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT112), .ZN(new_n1037));
  NAND3_X1  g612(.A1(G303), .A2(G8), .A3(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1036), .A2(KEYINPUT112), .ZN(new_n1039));
  XNOR2_X1  g614(.A(new_n1039), .B(KEYINPUT113), .ZN(new_n1040));
  XNOR2_X1  g615(.A(new_n1038), .B(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1012), .B1(new_n1006), .B2(KEYINPUT50), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT50), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n493), .A2(new_n1043), .A3(new_n1005), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT45), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1046), .A2(G1384), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n493), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G40), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n463), .A2(new_n468), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT45), .B1(new_n493), .B2(new_n1005), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  OAI22_X1  g628(.A1(new_n1045), .A2(G2090), .B1(new_n1053), .B2(G1971), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1041), .A2(new_n1054), .A3(G8), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT114), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1041), .A2(new_n1054), .A3(KEYINPUT114), .A4(G8), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1050), .A2(new_n493), .A3(new_n1005), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(G8), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1060), .A2(KEYINPUT115), .A3(G8), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(G1981), .B1(new_n568), .B2(new_n570), .ZN(new_n1066));
  INV_X1    g641(.A(new_n570), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT116), .B(G1981), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1067), .A2(new_n566), .A3(new_n567), .A4(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT117), .B1(new_n1066), .B2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1071), .A2(KEYINPUT49), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT49), .ZN(new_n1073));
  AOI211_X1 g648(.A(KEYINPUT117), .B(new_n1073), .C1(new_n1066), .C2(new_n1070), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1065), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n775), .A2(G1976), .A3(new_n776), .ZN(new_n1076));
  INV_X1    g651(.A(G1976), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT52), .B1(G288), .B2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1065), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1065), .A2(new_n1076), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1075), .B(new_n1079), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1059), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G288), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1075), .A2(new_n1077), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n1070), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1083), .B1(new_n1065), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1041), .B1(new_n1054), .B2(G8), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1082), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G1966), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g668(.A(KEYINPUT118), .B(new_n1090), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1042), .A2(new_n764), .A3(new_n1044), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1096), .A2(G8), .A3(G168), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1089), .A2(new_n1059), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT63), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1087), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT57), .B1(new_n559), .B2(KEYINPUT119), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n551), .A2(new_n1106), .ZN(new_n1107));
  OAI221_X1 g682(.A(KEYINPUT120), .B1(new_n501), .B2(new_n550), .C1(new_n505), .C2(new_n549), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n556), .A2(new_n1109), .A3(new_n558), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1107), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1103), .B1(new_n1105), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G1956), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1045), .A2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT56), .B(G2072), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1053), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1113), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(G1348), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1060), .A2(G2067), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1121), .A2(new_n587), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1113), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1118), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1113), .A2(new_n1115), .A3(new_n1125), .A4(new_n1117), .ZN(new_n1126));
  AOI21_X1  g701(.A(G1956), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1012), .B1(new_n493), .B2(new_n1047), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1006), .A2(new_n1046), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1128), .A2(new_n1129), .A3(new_n1116), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1112), .B(new_n1125), .C1(new_n1127), .C2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT61), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1126), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1132), .B1(new_n1126), .B2(new_n1131), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1121), .A2(KEYINPUT60), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT60), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1136), .A2(new_n588), .A3(new_n1138), .ZN(new_n1139));
  XOR2_X1   g714(.A(KEYINPUT58), .B(G1341), .Z(new_n1140));
  NAND2_X1  g715(.A1(new_n1060), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT121), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1060), .A2(KEYINPUT121), .A3(new_n1140), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1143), .B(new_n1144), .C1(new_n1145), .C2(G1996), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n542), .ZN(new_n1147));
  XNOR2_X1  g722(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1121), .A2(KEYINPUT60), .A3(new_n587), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1146), .A2(new_n1151), .A3(KEYINPUT59), .A4(new_n542), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1139), .A2(new_n1149), .A3(new_n1150), .A4(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1124), .B1(new_n1135), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT51), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1155), .B1(new_n1096), .B2(G286), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1093), .A2(G168), .A3(new_n1095), .A4(new_n1094), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(G8), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1155), .B1(new_n1157), .B2(G8), .ZN(new_n1160));
  OAI21_X1  g735(.A(KEYINPUT124), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(KEYINPUT126), .B(G2078), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1009), .A2(KEYINPUT53), .A3(new_n1128), .A4(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(G1961), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1045), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT53), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1166), .B1(new_n1145), .B2(G2078), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1163), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(KEYINPUT127), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT127), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1163), .A2(new_n1167), .A3(new_n1165), .A4(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1169), .A2(G171), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(G2078), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1053), .A2(KEYINPUT125), .A3(KEYINPUT53), .A4(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(KEYINPUT125), .A2(KEYINPUT53), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1175), .B1(new_n1145), .B2(G2078), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1174), .A2(new_n1176), .A3(new_n1165), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1177), .A2(G171), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT54), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1177), .A2(G171), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1181), .B1(G171), .B2(new_n1168), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n1172), .A2(new_n1180), .B1(new_n1182), .B2(new_n1179), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1158), .A2(KEYINPUT51), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT124), .ZN(new_n1185));
  OAI211_X1 g760(.A(new_n1184), .B(new_n1185), .C1(new_n1158), .C2(new_n1156), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1154), .A2(new_n1161), .A3(new_n1183), .A4(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1161), .A2(KEYINPUT62), .A3(new_n1186), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1181), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(KEYINPUT62), .B1(new_n1161), .B2(new_n1186), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1187), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  AND2_X1   g767(.A1(new_n1089), .A2(new_n1059), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1102), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(KEYINPUT110), .B1(G290), .B2(G1986), .ZN(new_n1195));
  NAND2_X1  g770(.A1(G290), .A2(G1986), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n1195), .B(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1197), .A2(new_n1013), .ZN(new_n1198));
  XNOR2_X1  g773(.A(new_n1198), .B(KEYINPUT111), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(new_n1022), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1035), .B1(new_n1194), .B2(new_n1200), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g776(.A(G319), .ZN(new_n1203));
  NOR2_X1   g777(.A1(G227), .A2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g778(.A(new_n1204), .B1(new_n674), .B2(new_n675), .ZN(new_n1205));
  AOI21_X1  g779(.A(new_n1205), .B1(new_n636), .B2(new_n638), .ZN(new_n1206));
  OAI211_X1 g780(.A(new_n1206), .B(new_n999), .C1(new_n929), .C2(new_n930), .ZN(G225));
  INV_X1    g781(.A(G225), .ZN(G308));
endmodule


