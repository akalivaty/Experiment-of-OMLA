//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 1 0 0 1 0 1 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n865, new_n866, new_n867, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988;
  INV_X1    g000(.A(KEYINPUT73), .ZN(new_n202));
  NOR2_X1   g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT66), .B1(new_n203), .B2(KEYINPUT23), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT66), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n205), .B(new_n206), .C1(G169gat), .C2(G176gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT67), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n212));
  AOI22_X1  g011(.A1(new_n211), .A2(new_n212), .B1(KEYINPUT23), .B2(new_n203), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n208), .A2(new_n213), .A3(KEYINPUT65), .ZN(new_n214));
  NAND2_X1  g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT24), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n218));
  INV_X1    g017(.A(G183gat), .ZN(new_n219));
  INV_X1    g018(.A(G190gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n217), .A2(new_n218), .A3(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n208), .A2(new_n213), .A3(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT25), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n214), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n223), .B1(new_n224), .B2(new_n214), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT68), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G169gat), .ZN(new_n228));
  INV_X1    g027(.A(G176gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n228), .A2(new_n229), .A3(KEYINPUT23), .ZN(new_n230));
  AND3_X1   g029(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n233), .B1(new_n204), .B2(new_n207), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n234), .B(new_n222), .C1(KEYINPUT65), .C2(KEYINPUT25), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n214), .A2(new_n223), .A3(new_n224), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT27), .B(G183gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(new_n220), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT28), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n203), .B(KEYINPUT26), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n243), .B1(new_n232), .B2(new_n231), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n242), .A2(new_n215), .A3(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n238), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G113gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n247), .A2(KEYINPUT70), .A3(G120gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT70), .ZN(new_n249));
  INV_X1    g048(.A(G120gat), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n249), .B1(G113gat), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(G113gat), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n248), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT71), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT71), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n255), .B(new_n248), .C1(new_n251), .C2(new_n252), .ZN(new_n256));
  INV_X1    g055(.A(G127gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G134gat), .ZN(new_n258));
  INV_X1    g057(.A(G134gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G127gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n254), .A2(new_n256), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n250), .A2(G113gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n247), .A2(G120gat), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT1), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n257), .A2(G134gat), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n268), .B1(KEYINPUT69), .B2(new_n258), .ZN(new_n269));
  OR2_X1    g068(.A1(new_n258), .A2(KEYINPUT69), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n267), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n264), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n246), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n235), .A2(new_n237), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n244), .A2(new_n215), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n275), .A2(KEYINPUT68), .B1(new_n242), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n262), .B1(new_n253), .B2(KEYINPUT71), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n271), .B1(new_n278), .B2(new_n256), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n279), .A3(new_n238), .ZN(new_n280));
  NAND2_X1  g079(.A1(G227gat), .A2(G233gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n274), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT34), .ZN(new_n283));
  XOR2_X1   g082(.A(new_n281), .B(KEYINPUT64), .Z(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n285), .A2(KEYINPUT34), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n274), .A2(new_n280), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT72), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT72), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n274), .A2(new_n280), .A3(new_n289), .A4(new_n286), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n283), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G15gat), .B(G43gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(G71gat), .B(G99gat), .ZN(new_n293));
  XOR2_X1   g092(.A(new_n292), .B(new_n293), .Z(new_n294));
  AOI21_X1  g093(.A(new_n284), .B1(new_n274), .B2(new_n280), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n294), .B1(new_n295), .B2(KEYINPUT33), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT32), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n274), .A2(new_n280), .ZN(new_n300));
  AOI221_X4 g099(.A(new_n297), .B1(KEYINPUT33), .B2(new_n294), .C1(new_n300), .C2(new_n285), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n291), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  AND3_X1   g101(.A1(new_n283), .A2(new_n288), .A3(new_n290), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n279), .B1(new_n277), .B2(new_n238), .ZN(new_n304));
  AND4_X1   g103(.A1(new_n279), .A2(new_n227), .A3(new_n238), .A4(new_n245), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n285), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT32), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT33), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n307), .A2(new_n309), .A3(new_n294), .ZN(new_n310));
  INV_X1    g109(.A(new_n294), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n306), .B(KEYINPUT32), .C1(new_n308), .C2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n303), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n202), .B1(new_n302), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n299), .A2(new_n301), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT73), .B1(new_n315), .B2(new_n303), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  XOR2_X1   g116(.A(G8gat), .B(G36gat), .Z(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G64gat), .B(G92gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n320), .B(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G211gat), .B(G218gat), .ZN(new_n324));
  OR2_X1    g123(.A1(G197gat), .A2(G204gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(G197gat), .A2(G204gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT22), .ZN(new_n327));
  NAND2_X1  g126(.A1(G211gat), .A2(G218gat), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n325), .A2(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT74), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n324), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n331), .B1(new_n330), .B2(new_n329), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT75), .ZN(new_n333));
  XNOR2_X1  g132(.A(G197gat), .B(G204gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n328), .A2(new_n327), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n324), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n333), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n329), .A2(KEYINPUT75), .A3(new_n324), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n332), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(G226gat), .A2(G233gat), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  AND3_X1   g142(.A1(new_n275), .A2(new_n245), .A3(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(KEYINPUT29), .ZN(new_n345));
  AOI211_X1 g144(.A(new_n341), .B(new_n344), .C1(new_n246), .C2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n341), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n227), .A2(new_n238), .A3(new_n245), .A4(new_n343), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n275), .A2(new_n245), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n345), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n347), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n323), .B1(new_n346), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n246), .A2(new_n345), .ZN(new_n353));
  INV_X1    g152(.A(new_n344), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n353), .A2(new_n347), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n348), .A2(new_n350), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n341), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n355), .A2(new_n357), .A3(new_n322), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n352), .A2(KEYINPUT30), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n344), .B1(new_n246), .B2(new_n345), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n351), .B1(new_n347), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT30), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(new_n362), .A3(new_n322), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT89), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n359), .A2(KEYINPUT89), .A3(new_n363), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT4), .ZN(new_n369));
  XNOR2_X1  g168(.A(G141gat), .B(G148gat), .ZN(new_n370));
  OR2_X1    g169(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(G155gat), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n370), .B1(new_n373), .B2(KEYINPUT2), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n375));
  NAND2_X1  g174(.A1(G155gat), .A2(G162gat), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(G155gat), .A2(G162gat), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n375), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OR2_X1    g178(.A1(G155gat), .A2(G162gat), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n380), .A2(KEYINPUT78), .A3(new_n376), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  XOR2_X1   g181(.A(G141gat), .B(G148gat), .Z(new_n383));
  INV_X1    g182(.A(KEYINPUT2), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n377), .A2(new_n378), .ZN(new_n386));
  AOI22_X1  g185(.A1(new_n374), .A2(new_n382), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n279), .A2(new_n369), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n369), .B1(new_n279), .B2(new_n387), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n388), .B1(new_n389), .B2(KEYINPUT83), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n382), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n385), .A2(new_n386), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n273), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT83), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n394), .A2(new_n395), .A3(new_n369), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT80), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT3), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n397), .B1(new_n387), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n387), .A2(new_n398), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n399), .A2(new_n273), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n393), .A2(KEYINPUT80), .A3(KEYINPUT3), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n390), .A2(new_n396), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(G225gat), .A2(G233gat), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n405), .A2(KEYINPUT5), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n402), .A2(new_n399), .A3(new_n273), .A4(new_n400), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n404), .ZN(new_n409));
  AOI211_X1 g208(.A(KEYINPUT81), .B(new_n369), .C1(new_n279), .C2(new_n387), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT81), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n388), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n413), .B1(new_n369), .B2(new_n394), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n409), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT82), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n416), .B1(new_n279), .B2(new_n387), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n273), .A2(new_n393), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n273), .A2(new_n416), .A3(new_n393), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n419), .A2(new_n405), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT5), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n407), .B1(new_n415), .B2(new_n422), .ZN(new_n423));
  XOR2_X1   g222(.A(G1gat), .B(G29gat), .Z(new_n424));
  XNOR2_X1  g223(.A(new_n424), .B(G85gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT0), .B(G57gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  NAND3_X1  g226(.A1(new_n423), .A2(KEYINPUT6), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n421), .A2(KEYINPUT5), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n389), .B1(new_n412), .B2(new_n388), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n404), .B(new_n408), .C1(new_n431), .C2(new_n410), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n430), .A2(new_n432), .B1(new_n403), .B2(new_n406), .ZN(new_n433));
  INV_X1    g232(.A(new_n427), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n429), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n407), .B(new_n434), .C1(new_n415), .C2(new_n422), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n428), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT35), .ZN(new_n439));
  XNOR2_X1  g238(.A(G78gat), .B(G106gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT31), .B(G50gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n440), .B(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n442), .B(KEYINPUT85), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n338), .A2(new_n339), .B1(new_n337), .B2(new_n336), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n398), .B1(new_n444), .B2(KEYINPUT29), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n393), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT29), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n400), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n347), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(G228gat), .A2(G233gat), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT29), .B1(new_n332), .B2(new_n340), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n393), .B1(new_n452), .B2(KEYINPUT3), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n451), .B1(new_n448), .B2(new_n347), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n450), .A2(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  XOR2_X1   g254(.A(KEYINPUT86), .B(G22gat), .Z(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n454), .A2(new_n453), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n446), .A2(new_n449), .B1(G228gat), .B2(G233gat), .ZN(new_n460));
  NOR3_X1   g259(.A1(new_n459), .A2(new_n460), .A3(new_n456), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n443), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  NOR4_X1   g261(.A1(new_n459), .A2(new_n460), .A3(KEYINPUT88), .A4(new_n456), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT88), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n464), .B1(new_n455), .B2(new_n457), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT87), .ZN(new_n467));
  INV_X1    g266(.A(G22gat), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n467), .B1(new_n455), .B2(new_n468), .ZN(new_n469));
  OAI211_X1 g268(.A(KEYINPUT87), .B(G22gat), .C1(new_n459), .C2(new_n460), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(new_n442), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n462), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n438), .A2(new_n439), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n317), .A2(new_n368), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n423), .A2(new_n427), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT84), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n475), .A2(new_n476), .A3(new_n429), .A4(new_n436), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n428), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT6), .B1(new_n423), .B2(new_n427), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n476), .B1(new_n479), .B2(new_n436), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n364), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n302), .A2(new_n472), .A3(new_n313), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT35), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n474), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT36), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n485), .B1(new_n314), .B2(new_n316), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n299), .A2(new_n291), .A3(new_n301), .ZN(new_n487));
  AOI22_X1  g286(.A1(KEYINPUT72), .A2(new_n287), .B1(new_n282), .B2(KEYINPUT34), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n310), .A2(new_n312), .B1(new_n290), .B2(new_n488), .ZN(new_n489));
  NOR3_X1   g288(.A1(new_n487), .A2(new_n489), .A3(new_n485), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT39), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n419), .A2(new_n420), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n494), .B1(new_n495), .B2(new_n404), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n496), .B1(new_n403), .B2(new_n404), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n390), .A2(new_n396), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n408), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(new_n494), .A3(new_n405), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(new_n500), .A3(new_n434), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT90), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n502), .A2(KEYINPUT40), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n503), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n497), .A2(new_n500), .A3(new_n434), .A4(new_n505), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n504), .A2(new_n475), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n507), .A2(new_n366), .A3(new_n367), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n322), .B1(new_n355), .B2(new_n357), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT37), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n322), .A2(new_n510), .ZN(new_n511));
  OAI22_X1  g310(.A1(new_n509), .A2(new_n511), .B1(new_n361), .B2(new_n510), .ZN(new_n512));
  AOI22_X1  g311(.A1(new_n512), .A2(KEYINPUT38), .B1(new_n361), .B2(new_n322), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n479), .A2(new_n436), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n510), .B1(new_n356), .B2(new_n347), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n360), .A2(new_n341), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT91), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n322), .B1(new_n361), .B2(new_n510), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT38), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT91), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n518), .A2(new_n519), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n513), .A2(new_n514), .A3(new_n522), .A4(new_n428), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n508), .A2(new_n472), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n472), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n481), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n484), .B1(new_n493), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G64gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(G57gat), .ZN(new_n530));
  XOR2_X1   g329(.A(KEYINPUT95), .B(G57gat), .Z(new_n531));
  OAI21_X1  g330(.A(new_n530), .B1(new_n531), .B2(new_n529), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT96), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g333(.A(KEYINPUT96), .B(new_n530), .C1(new_n531), .C2(new_n529), .ZN(new_n535));
  NOR2_X1   g334(.A1(G71gat), .A2(G78gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT9), .ZN(new_n537));
  NAND2_X1  g336(.A1(G71gat), .A2(G78gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n534), .A2(new_n535), .A3(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(G57gat), .B(G64gat), .Z(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT9), .ZN(new_n542));
  INV_X1    g341(.A(new_n538), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n543), .A2(new_n536), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT7), .ZN(new_n547));
  NAND2_X1  g346(.A1(G85gat), .A2(G92gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(G99gat), .A2(G106gat), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n547), .A2(new_n548), .B1(new_n549), .B2(KEYINPUT8), .ZN(new_n550));
  XNOR2_X1  g349(.A(KEYINPUT99), .B(G85gat), .ZN(new_n551));
  OAI221_X1 g350(.A(new_n550), .B1(new_n547), .B2(new_n548), .C1(G92gat), .C2(new_n551), .ZN(new_n552));
  XOR2_X1   g351(.A(G99gat), .B(G106gat), .Z(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT102), .B1(new_n546), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT10), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT102), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n552), .A2(new_n553), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n552), .A2(new_n553), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n545), .ZN(new_n562));
  AOI22_X1  g361(.A1(new_n532), .A2(new_n533), .B1(new_n538), .B2(new_n537), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n562), .B1(new_n563), .B2(new_n535), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n558), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT10), .ZN(new_n566));
  NAND2_X1  g365(.A1(G230gat), .A2(G233gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n546), .A2(new_n554), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n557), .A2(new_n566), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n554), .B(new_n564), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n569), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G120gat), .B(G148gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(G176gat), .B(G204gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n571), .A2(new_n574), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G15gat), .B(G22gat), .ZN(new_n578));
  INV_X1    g377(.A(G1gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT16), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n581), .B1(G1gat), .B2(new_n578), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(G8gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT14), .ZN(new_n585));
  INV_X1    g384(.A(G29gat), .ZN(new_n586));
  INV_X1    g385(.A(G36gat), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n590), .A2(KEYINPUT94), .ZN(new_n591));
  XNOR2_X1  g390(.A(G43gat), .B(G50gat), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT15), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n592), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n590), .A2(KEYINPUT94), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n591), .A2(new_n595), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n593), .A2(new_n594), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT93), .ZN(new_n600));
  OAI22_X1  g399(.A1(new_n590), .A2(new_n600), .B1(new_n586), .B2(new_n587), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT93), .B1(new_n588), .B2(new_n589), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n599), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT17), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n598), .A2(new_n603), .A3(KEYINPUT17), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n584), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G229gat), .A2(G233gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n583), .A2(new_n604), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT18), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n608), .A2(KEYINPUT18), .A3(new_n609), .A4(new_n610), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n609), .B(KEYINPUT13), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n610), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n583), .A2(new_n604), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n613), .A2(new_n614), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G113gat), .B(G141gat), .Z(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT92), .B(G197gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(KEYINPUT11), .B(G169gat), .Z(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n620), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n613), .A2(new_n626), .A3(new_n614), .A4(new_n619), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n577), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n583), .B1(new_n564), .B2(KEYINPUT21), .ZN(new_n633));
  XOR2_X1   g432(.A(KEYINPUT97), .B(KEYINPUT19), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(G127gat), .B(G155gat), .Z(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT20), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n635), .B(new_n637), .Z(new_n638));
  OR2_X1    g437(.A1(new_n564), .A2(KEYINPUT21), .ZN(new_n639));
  NAND2_X1  g438(.A1(G231gat), .A2(G233gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(new_n219), .ZN(new_n641));
  INV_X1    g440(.A(G211gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n639), .B(new_n643), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n638), .B(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n606), .A2(new_n607), .A3(new_n554), .ZN(new_n646));
  NAND2_X1  g445(.A1(G232gat), .A2(G233gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT98), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT41), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n650), .B1(new_n561), .B2(new_n604), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g451(.A(G190gat), .B(G218gat), .Z(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(KEYINPUT100), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n655), .B1(new_n654), .B2(new_n652), .ZN(new_n656));
  INV_X1    g455(.A(new_n652), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n657), .A2(KEYINPUT100), .A3(new_n653), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n648), .A2(new_n649), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(new_n259), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(G162gat), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n652), .A2(new_n654), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n662), .B1(new_n663), .B2(KEYINPUT101), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n659), .B(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n645), .A2(new_n666), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n528), .A2(new_n632), .A3(new_n667), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n478), .A2(new_n480), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(G1gat), .ZN(G1324gat));
  INV_X1    g471(.A(new_n368), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n668), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(G8gat), .ZN(new_n675));
  OAI21_X1  g474(.A(KEYINPUT42), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT103), .B(KEYINPUT16), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(new_n675), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  MUX2_X1   g478(.A(KEYINPUT42), .B(new_n676), .S(new_n679), .Z(G1325gat));
  AOI21_X1  g479(.A(G15gat), .B1(new_n668), .B2(new_n317), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT104), .ZN(new_n682));
  OAI21_X1  g481(.A(KEYINPUT73), .B1(new_n487), .B2(new_n489), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n313), .A2(new_n202), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT36), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n682), .B1(new_n685), .B2(new_n490), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n486), .A2(KEYINPUT104), .A3(new_n491), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n689), .A2(G15gat), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n681), .B1(new_n668), .B2(new_n690), .ZN(new_n691));
  XOR2_X1   g490(.A(new_n691), .B(KEYINPUT105), .Z(G1326gat));
  NAND2_X1  g491(.A1(new_n668), .A2(new_n525), .ZN(new_n693));
  XNOR2_X1  g492(.A(KEYINPUT43), .B(G22gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1327gat));
  NAND2_X1  g494(.A1(new_n355), .A2(new_n357), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n520), .B(new_n323), .C1(new_n696), .C2(KEYINPUT37), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT91), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n697), .A2(new_n517), .A3(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n438), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n525), .B1(new_n700), .B2(new_n513), .ZN(new_n701));
  AOI22_X1  g500(.A1(new_n701), .A2(new_n508), .B1(new_n481), .B2(new_n525), .ZN(new_n702));
  AOI22_X1  g501(.A1(new_n702), .A2(new_n492), .B1(new_n483), .B2(new_n474), .ZN(new_n703));
  INV_X1    g502(.A(new_n666), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n645), .A2(new_n632), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n706), .A2(new_n586), .A3(new_n670), .ZN(new_n707));
  XOR2_X1   g506(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n527), .B1(new_n686), .B2(new_n687), .ZN(new_n711));
  INV_X1    g510(.A(new_n484), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n710), .B(new_n666), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT44), .B1(new_n703), .B2(new_n704), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n705), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(G29gat), .B1(new_n717), .B2(new_n669), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n709), .A2(new_n718), .ZN(G1328gat));
  NAND3_X1  g518(.A1(new_n706), .A2(new_n587), .A3(new_n673), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT46), .Z(new_n721));
  OAI21_X1  g520(.A(G36gat), .B1(new_n717), .B2(new_n368), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(G1329gat));
  NAND3_X1  g522(.A1(new_n715), .A2(new_n689), .A3(new_n716), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(G43gat), .ZN(new_n725));
  INV_X1    g524(.A(new_n317), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(G43gat), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n528), .A2(new_n666), .A3(new_n716), .A4(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n725), .A2(KEYINPUT47), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(KEYINPUT107), .ZN(new_n730));
  AOI211_X1 g529(.A(KEYINPUT108), .B(KEYINPUT47), .C1(new_n725), .C2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n732));
  AOI211_X1 g531(.A(new_n688), .B(new_n705), .C1(new_n713), .C2(new_n714), .ZN(new_n733));
  INV_X1    g532(.A(G43gat), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n730), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n732), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n729), .B1(new_n731), .B2(new_n737), .ZN(G1330gat));
  INV_X1    g537(.A(G50gat), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n706), .A2(new_n739), .A3(new_n525), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n717), .A2(new_n472), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n741), .B2(new_n739), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT48), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI211_X1 g543(.A(KEYINPUT48), .B(new_n740), .C1(new_n741), .C2(new_n739), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(G1331gat));
  AND3_X1   g545(.A1(new_n486), .A2(KEYINPUT104), .A3(new_n491), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT104), .B1(new_n486), .B2(new_n491), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n702), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n484), .ZN(new_n750));
  AND4_X1   g549(.A1(new_n631), .A2(new_n750), .A3(new_n577), .A4(new_n667), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n670), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(new_n531), .ZN(G1332gat));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n673), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n755));
  XOR2_X1   g554(.A(KEYINPUT49), .B(G64gat), .Z(new_n756));
  OAI21_X1  g555(.A(new_n755), .B1(new_n754), .B2(new_n756), .ZN(G1333gat));
  NAND2_X1  g556(.A1(new_n751), .A2(new_n689), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(G71gat), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n760));
  INV_X1    g559(.A(G71gat), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n317), .B(KEYINPUT109), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n751), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n759), .A2(new_n760), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n760), .B1(new_n759), .B2(new_n763), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n764), .A2(new_n765), .ZN(G1334gat));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n525), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g567(.A1(new_n645), .A2(new_n631), .ZN(new_n769));
  INV_X1    g568(.A(new_n577), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n772), .B1(new_n713), .B2(new_n714), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n551), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n774), .A2(new_n669), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n769), .B1(KEYINPUT110), .B2(new_n777), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n666), .B(new_n778), .C1(new_n711), .C2(new_n712), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n777), .A2(KEYINPUT110), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n780), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n750), .A2(new_n666), .A3(new_n782), .A4(new_n778), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n781), .A2(new_n783), .A3(new_n577), .ZN(new_n784));
  OR2_X1    g583(.A1(new_n784), .A2(new_n669), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n776), .B1(new_n785), .B2(new_n775), .ZN(G1336gat));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n368), .A2(G92gat), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n781), .A2(new_n783), .A3(new_n577), .A4(new_n788), .ZN(new_n789));
  AOI211_X1 g588(.A(new_n368), .B(new_n772), .C1(new_n713), .C2(new_n714), .ZN(new_n790));
  OAI21_X1  g589(.A(G92gat), .B1(new_n790), .B2(KEYINPUT112), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n715), .A2(new_n673), .A3(new_n771), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n787), .B(new_n789), .C1(new_n791), .C2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n792), .A2(G92gat), .ZN(new_n797));
  AOI211_X1 g596(.A(new_n796), .B(new_n787), .C1(new_n797), .C2(new_n789), .ZN(new_n798));
  INV_X1    g597(.A(G92gat), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n789), .B1(new_n790), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT111), .B1(new_n800), .B2(KEYINPUT52), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n795), .B1(new_n798), .B2(new_n801), .ZN(G1337gat));
  OAI21_X1  g601(.A(G99gat), .B1(new_n774), .B2(new_n688), .ZN(new_n803));
  OR2_X1    g602(.A1(new_n726), .A2(G99gat), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n803), .B1(new_n784), .B2(new_n804), .ZN(G1338gat));
  INV_X1    g604(.A(G106gat), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n806), .B1(new_n784), .B2(new_n472), .ZN(new_n807));
  NAND2_X1  g606(.A1(KEYINPUT113), .A2(KEYINPUT53), .ZN(new_n808));
  NOR2_X1   g607(.A1(KEYINPUT113), .A2(KEYINPUT53), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n472), .A2(new_n806), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n809), .B1(new_n773), .B2(new_n810), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n807), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n808), .B1(new_n807), .B2(new_n811), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n812), .A2(new_n813), .ZN(G1339gat));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n569), .A2(KEYINPUT54), .ZN(new_n816));
  INV_X1    g615(.A(new_n568), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n817), .B1(new_n555), .B2(new_n556), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n567), .B1(new_n818), .B2(new_n566), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n818), .A2(new_n821), .A3(new_n567), .A4(new_n566), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n574), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n815), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n568), .B1(new_n565), .B2(KEYINPUT10), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n555), .A2(new_n556), .ZN(new_n826));
  OAI211_X1 g625(.A(G230gat), .B(G233gat), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n827), .A2(KEYINPUT54), .A3(new_n569), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n828), .A2(KEYINPUT55), .A3(new_n574), .A4(new_n822), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n824), .A2(new_n630), .A3(new_n575), .A4(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n609), .B1(new_n608), .B2(new_n610), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n617), .A2(new_n618), .A3(new_n616), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n625), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n629), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n577), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n830), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n704), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n659), .A2(new_n665), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n664), .B1(new_n656), .B2(new_n658), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n834), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n824), .A2(new_n575), .A3(new_n829), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n837), .A2(KEYINPUT114), .A3(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT114), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n666), .B1(new_n830), .B2(new_n835), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n840), .A2(new_n841), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n843), .A2(new_n645), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n667), .A2(new_n631), .A3(new_n770), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n472), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT115), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n850), .A2(new_n853), .A3(new_n472), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n855), .A2(new_n670), .A3(new_n317), .A4(new_n368), .ZN(new_n856));
  OAI21_X1  g655(.A(G113gat), .B1(new_n856), .B2(new_n631), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n670), .A2(new_n368), .ZN(new_n858));
  AOI211_X1 g657(.A(new_n482), .B(new_n858), .C1(new_n848), .C2(new_n849), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n247), .A3(new_n630), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n857), .A2(new_n860), .ZN(G1340gat));
  OAI21_X1  g660(.A(G120gat), .B1(new_n856), .B2(new_n770), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n859), .A2(new_n250), .A3(new_n577), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(G1341gat));
  NOR3_X1   g663(.A1(new_n856), .A2(new_n257), .A3(new_n645), .ZN(new_n865));
  INV_X1    g664(.A(new_n645), .ZN(new_n866));
  AOI21_X1  g665(.A(G127gat), .B1(new_n859), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n865), .A2(new_n867), .ZN(G1342gat));
  NAND3_X1  g667(.A1(new_n859), .A2(new_n259), .A3(new_n666), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n869), .A2(KEYINPUT56), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n870), .A2(KEYINPUT116), .ZN(new_n871));
  OAI21_X1  g670(.A(G134gat), .B1(new_n856), .B2(new_n704), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n869), .A2(KEYINPUT56), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n870), .A2(KEYINPUT116), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n871), .A2(new_n872), .A3(new_n873), .A4(new_n874), .ZN(G1343gat));
  NAND3_X1  g674(.A1(new_n688), .A2(new_n670), .A3(new_n368), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n472), .B1(new_n848), .B2(new_n849), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n631), .A2(G141gat), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT119), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT58), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n645), .B1(new_n845), .B2(new_n846), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n849), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(KEYINPUT57), .A3(new_n525), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT117), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n886), .A2(KEYINPUT117), .A3(KEYINPUT57), .A4(new_n525), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT57), .B1(new_n850), .B2(new_n525), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n630), .B(new_n877), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT120), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(G141gat), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n893), .A2(KEYINPUT120), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n882), .B(new_n884), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n893), .A2(KEYINPUT118), .A3(G141gat), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT118), .B1(new_n893), .B2(G141gat), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n898), .A2(new_n899), .A3(new_n881), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT58), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n897), .B1(new_n900), .B2(new_n901), .ZN(G1344gat));
  NAND2_X1  g701(.A1(new_n877), .A2(new_n878), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(G148gat), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(new_n905), .A3(new_n577), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n891), .A2(new_n892), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n907), .A2(new_n689), .A3(new_n858), .ZN(new_n908));
  AOI211_X1 g707(.A(KEYINPUT59), .B(new_n905), .C1(new_n908), .C2(new_n577), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT59), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n876), .B(KEYINPUT121), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n850), .A2(KEYINPUT57), .A3(new_n525), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n472), .B1(new_n885), .B2(new_n849), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n913), .A2(KEYINPUT57), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n911), .A2(new_n577), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n910), .B1(new_n916), .B2(G148gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n906), .B1(new_n909), .B2(new_n917), .ZN(G1345gat));
  AOI21_X1  g717(.A(G155gat), .B1(new_n904), .B2(new_n866), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n866), .A2(G155gat), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n919), .B1(new_n908), .B2(new_n920), .ZN(G1346gat));
  NAND2_X1  g720(.A1(new_n371), .A2(new_n372), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n704), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n904), .A2(new_n666), .ZN(new_n924));
  AOI22_X1  g723(.A1(new_n908), .A2(new_n923), .B1(new_n924), .B2(new_n922), .ZN(G1347gat));
  AOI21_X1  g724(.A(new_n670), .B1(new_n848), .B2(new_n849), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n368), .A2(new_n482), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT122), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(new_n228), .A3(new_n630), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n670), .A2(new_n368), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n762), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n933), .B1(new_n852), .B2(new_n854), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n934), .A2(new_n630), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n931), .B1(new_n935), .B2(new_n228), .ZN(G1348gat));
  AOI21_X1  g735(.A(G176gat), .B1(new_n930), .B2(new_n577), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n770), .A2(new_n229), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n937), .B1(new_n934), .B2(new_n938), .ZN(G1349gat));
  AND3_X1   g738(.A1(new_n930), .A2(new_n239), .A3(new_n866), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n934), .A2(new_n866), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n941), .B2(G183gat), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT60), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n942), .B(new_n943), .ZN(G1350gat));
  NAND3_X1  g743(.A1(new_n930), .A2(new_n220), .A3(new_n666), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n934), .A2(new_n666), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n946), .B1(new_n947), .B2(G190gat), .ZN(new_n948));
  AOI211_X1 g747(.A(KEYINPUT61), .B(new_n220), .C1(new_n934), .C2(new_n666), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(G1351gat));
  NAND2_X1  g749(.A1(new_n850), .A2(new_n669), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT123), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n688), .A2(new_n525), .A3(new_n673), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n953), .A2(new_n952), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n631), .A2(G197gat), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  XOR2_X1   g756(.A(new_n957), .B(KEYINPUT124), .Z(new_n958));
  AND3_X1   g757(.A1(new_n688), .A2(KEYINPUT125), .A3(new_n932), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT125), .B1(new_n688), .B2(new_n932), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n961), .A2(new_n630), .A3(new_n915), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(G197gat), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n958), .A2(new_n963), .ZN(G1352gat));
  AND2_X1   g763(.A1(new_n954), .A2(new_n955), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n770), .A2(G204gat), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OR2_X1    g766(.A1(new_n967), .A2(KEYINPUT62), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n961), .A2(new_n577), .A3(new_n915), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(G204gat), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n967), .A2(KEYINPUT62), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n968), .A2(new_n970), .A3(new_n971), .ZN(G1353gat));
  NAND3_X1  g771(.A1(new_n965), .A2(new_n642), .A3(new_n866), .ZN(new_n973));
  OAI211_X1 g772(.A(new_n915), .B(new_n866), .C1(new_n960), .C2(new_n959), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(KEYINPUT126), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n961), .A2(new_n976), .A3(new_n866), .A4(new_n915), .ZN(new_n977));
  AND4_X1   g776(.A1(KEYINPUT63), .A2(new_n975), .A3(new_n977), .A4(G211gat), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n642), .B1(new_n974), .B2(KEYINPUT126), .ZN(new_n979));
  AOI21_X1  g778(.A(KEYINPUT63), .B1(new_n979), .B2(new_n977), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n973), .B1(new_n978), .B2(new_n980), .ZN(G1354gat));
  NOR2_X1   g780(.A1(new_n704), .A2(G218gat), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n965), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n961), .A2(new_n666), .A3(new_n915), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(G218gat), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT127), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n983), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n986), .B1(new_n983), .B2(new_n985), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n987), .A2(new_n988), .ZN(G1355gat));
endmodule


