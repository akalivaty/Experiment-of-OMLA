//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 0 1 0 0 0 1 1 1 0 0 0 0 0 0 1 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n805, new_n806, new_n807, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XOR2_X1   g002(.A(KEYINPUT2), .B(G113), .Z(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G116), .ZN(new_n191));
  INV_X1    g005(.A(G116), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G119), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n189), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(new_n193), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT2), .B(G113), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G101), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT75), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n200), .A2(KEYINPUT75), .ZN(new_n202));
  INV_X1    g016(.A(G107), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G104), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n201), .B1(new_n202), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G104), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G107), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n200), .A2(new_n203), .A3(KEYINPUT75), .A4(G104), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n199), .B1(new_n209), .B2(KEYINPUT76), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT76), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n205), .A2(new_n211), .A3(new_n207), .A4(new_n208), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n205), .A2(new_n199), .A3(new_n207), .A4(new_n208), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n210), .A2(new_n212), .B1(KEYINPUT4), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT75), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(KEYINPUT3), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n206), .A2(G107), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(KEYINPUT3), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n208), .A2(new_n207), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT76), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n221), .A2(new_n212), .A3(KEYINPUT4), .A4(G101), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n198), .B1(new_n214), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n204), .A2(new_n207), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G101), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n213), .A2(new_n226), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT5), .ZN(new_n228));
  OAI21_X1  g042(.A(G113), .B1(new_n191), .B2(KEYINPUT5), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n194), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(G110), .B(G122), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n224), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n233), .ZN(new_n235));
  INV_X1    g049(.A(new_n198), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n221), .A2(G101), .A3(new_n212), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n213), .A2(KEYINPUT4), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n236), .B1(new_n239), .B2(new_n222), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n235), .B1(new_n240), .B2(new_n231), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n234), .A2(new_n241), .A3(KEYINPUT6), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT6), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n243), .B(new_n235), .C1(new_n240), .C2(new_n231), .ZN(new_n244));
  INV_X1    g058(.A(G146), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G143), .ZN(new_n246));
  INV_X1    g060(.A(G143), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G146), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  AND2_X1   g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  OR2_X1    g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT64), .ZN(new_n254));
  XNOR2_X1  g068(.A(G143), .B(G146), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n254), .B1(new_n255), .B2(new_n250), .ZN(new_n256));
  AND4_X1   g070(.A1(new_n254), .A2(new_n246), .A3(new_n248), .A4(new_n250), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n253), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G125), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT1), .ZN(new_n260));
  OAI22_X1  g074(.A1(new_n255), .A2(G128), .B1(new_n260), .B2(new_n248), .ZN(new_n261));
  INV_X1    g075(.A(G128), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(KEYINPUT1), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(new_n246), .A3(new_n248), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G125), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n259), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G224), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n270), .A2(G953), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n269), .B(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n242), .A2(new_n244), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n271), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT7), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n246), .A2(new_n248), .A3(new_n250), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT64), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n255), .A2(new_n254), .A3(new_n250), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n267), .B1(new_n279), .B2(new_n253), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n247), .A2(KEYINPUT1), .A3(G146), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n281), .B1(new_n249), .B2(new_n262), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n264), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(G125), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n275), .B1(new_n280), .B2(new_n284), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n259), .A2(new_n268), .A3(KEYINPUT7), .A4(new_n274), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT80), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n230), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n227), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n194), .B(KEYINPUT80), .C1(new_n228), .C2(new_n229), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n289), .A2(new_n290), .A3(KEYINPUT81), .A4(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n233), .B(KEYINPUT8), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT81), .B1(new_n227), .B2(new_n230), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n287), .B1(new_n294), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(G902), .B1(new_n298), .B2(new_n234), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n273), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G210), .B1(G237), .B2(G902), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n273), .A2(new_n299), .A3(new_n301), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n188), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(G237), .A2(G953), .ZN(new_n306));
  AOI21_X1  g120(.A(G143), .B1(new_n306), .B2(G214), .ZN(new_n307));
  NAND2_X1  g121(.A1(G143), .A2(G214), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n308), .A2(G237), .A3(G953), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(KEYINPUT18), .A2(G131), .ZN(new_n311));
  INV_X1    g125(.A(G140), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G125), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n267), .A2(G140), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G146), .ZN(new_n316));
  XNOR2_X1  g130(.A(G125), .B(G140), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n245), .ZN(new_n318));
  AOI22_X1  g132(.A1(new_n310), .A2(new_n311), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  OAI211_X1 g133(.A(KEYINPUT18), .B(G131), .C1(new_n307), .C2(new_n309), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT82), .ZN(new_n322));
  INV_X1    g136(.A(G131), .ZN(new_n323));
  INV_X1    g137(.A(G237), .ZN(new_n324));
  INV_X1    g138(.A(G953), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n323), .B1(new_n326), .B2(new_n308), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n322), .B1(new_n327), .B2(new_n307), .ZN(new_n328));
  INV_X1    g142(.A(G214), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n247), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  AND2_X1   g144(.A1(G143), .A2(G214), .ZN(new_n331));
  AOI21_X1  g145(.A(G131), .B1(new_n331), .B2(new_n306), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n330), .A2(KEYINPUT82), .A3(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(G131), .B1(new_n307), .B2(new_n309), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT17), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n328), .A2(new_n333), .A3(new_n334), .A4(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT84), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n267), .A2(KEYINPUT16), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n245), .B1(new_n338), .B2(new_n312), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT16), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT71), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n339), .A2(KEYINPUT71), .A3(new_n340), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n338), .A2(new_n312), .ZN(new_n345));
  AOI21_X1  g159(.A(G146), .B1(new_n340), .B2(new_n345), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n343), .A2(new_n344), .B1(KEYINPUT72), .B2(new_n346), .ZN(new_n347));
  OR2_X1    g161(.A1(new_n346), .A2(KEYINPUT72), .ZN(new_n348));
  OR2_X1    g162(.A1(new_n334), .A2(new_n335), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n337), .A2(new_n347), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n336), .A2(KEYINPUT84), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n321), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(G113), .B(G122), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n353), .B(new_n206), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n354), .B(new_n321), .C1(new_n350), .C2(new_n351), .ZN(new_n357));
  AOI21_X1  g171(.A(G902), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G475), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT19), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n315), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n317), .A2(KEYINPUT19), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n364), .A2(new_n245), .B1(new_n340), .B2(new_n339), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n328), .A2(new_n333), .A3(new_n334), .ZN(new_n366));
  AOI22_X1  g180(.A1(new_n365), .A2(new_n366), .B1(new_n319), .B2(new_n320), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT83), .B1(new_n367), .B2(new_n354), .ZN(new_n368));
  INV_X1    g182(.A(new_n366), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n315), .A2(new_n361), .ZN(new_n370));
  AOI21_X1  g184(.A(KEYINPUT19), .B1(new_n313), .B2(new_n314), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n245), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n341), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n321), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT83), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n375), .A3(new_n355), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n368), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n357), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT85), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(G475), .A2(G902), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n377), .A2(new_n357), .A3(KEYINPUT85), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT20), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT20), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n378), .A2(new_n385), .A3(new_n381), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n360), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G952), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n388), .A2(G953), .ZN(new_n389));
  INV_X1    g203(.A(G234), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n389), .B1(new_n390), .B2(new_n324), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  OAI211_X1 g206(.A(G902), .B(G953), .C1(new_n390), .C2(new_n324), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(KEYINPUT92), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT21), .B(G898), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n392), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G478), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(KEYINPUT15), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT86), .B1(new_n192), .B2(G122), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT86), .ZN(new_n402));
  INV_X1    g216(.A(G122), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(G116), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT87), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n406), .B1(new_n403), .B2(G116), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n192), .A2(KEYINPUT87), .A3(G122), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT88), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n405), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n410), .B1(new_n405), .B2(new_n409), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n203), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT90), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n247), .A2(G128), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n262), .A2(G143), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n415), .A2(new_n416), .A3(new_n414), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(G134), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G134), .ZN(new_n421));
  INV_X1    g235(.A(new_n419), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n421), .B1(new_n422), .B2(new_n417), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n409), .A2(KEYINPUT14), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n405), .B1(new_n409), .B2(KEYINPUT14), .ZN(new_n426));
  OAI21_X1  g240(.A(G107), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n413), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT89), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n247), .A2(G128), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT13), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n429), .B(new_n415), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n262), .A2(G143), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n433), .B1(KEYINPUT13), .B2(new_n416), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT89), .B1(new_n415), .B2(new_n431), .ZN(new_n435));
  OAI211_X1 g249(.A(G134), .B(new_n432), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n423), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n405), .A2(new_n409), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT88), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n405), .A2(new_n409), .A3(new_n410), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(G107), .A3(new_n440), .ZN(new_n441));
  AOI211_X1 g255(.A(KEYINPUT91), .B(new_n437), .C1(new_n441), .C2(new_n413), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT91), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n413), .A2(new_n441), .ZN(new_n444));
  INV_X1    g258(.A(new_n437), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n428), .B1(new_n442), .B2(new_n446), .ZN(new_n447));
  XOR2_X1   g261(.A(KEYINPUT9), .B(G234), .Z(new_n448));
  XNOR2_X1  g262(.A(new_n448), .B(KEYINPUT74), .ZN(new_n449));
  XOR2_X1   g263(.A(KEYINPUT70), .B(G217), .Z(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n325), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n447), .A2(new_n452), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n411), .A2(new_n412), .A3(new_n203), .ZN(new_n454));
  AOI21_X1  g268(.A(G107), .B1(new_n439), .B2(new_n440), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n445), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT91), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n444), .A2(new_n443), .A3(new_n445), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n452), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n428), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n453), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G902), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n400), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AOI211_X1 g278(.A(G902), .B(new_n399), .C1(new_n453), .C2(new_n461), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n305), .A2(new_n387), .A3(new_n397), .A4(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT79), .ZN(new_n468));
  XNOR2_X1  g282(.A(G110), .B(G140), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n325), .A2(G227), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n469), .B(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G137), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT65), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT65), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G137), .ZN(new_n476));
  AND2_X1   g290(.A1(KEYINPUT11), .A2(G134), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(KEYINPUT11), .A2(G134), .ZN(new_n479));
  NOR2_X1   g293(.A1(KEYINPUT11), .A2(G134), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n479), .B1(new_n480), .B2(G137), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n478), .A2(new_n323), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n323), .B1(new_n478), .B2(new_n481), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n227), .A2(new_n266), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n264), .A2(KEYINPUT77), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT77), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n255), .A2(new_n487), .A3(new_n263), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n282), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(new_n213), .A3(new_n226), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n484), .B1(new_n485), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(KEYINPUT12), .ZN(new_n492));
  INV_X1    g306(.A(new_n258), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(new_n214), .B2(new_n223), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT10), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n266), .A2(new_n495), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n495), .A2(new_n490), .B1(new_n496), .B2(new_n290), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n494), .A2(new_n484), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n472), .B1(new_n492), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n484), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n258), .B1(new_n239), .B2(new_n222), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n282), .A2(new_n486), .A3(new_n488), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n495), .B1(new_n502), .B2(new_n227), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n283), .A2(KEYINPUT10), .A3(new_n213), .A4(new_n226), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n500), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n498), .A2(new_n506), .A3(new_n472), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n463), .B1(new_n499), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n484), .B1(new_n494), .B2(new_n497), .ZN(new_n509));
  NOR3_X1   g323(.A1(new_n501), .A2(new_n505), .A3(new_n500), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n471), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT12), .ZN(new_n512));
  OR2_X1    g326(.A1(new_n491), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n491), .A2(new_n512), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n498), .A2(new_n513), .A3(new_n514), .A4(new_n472), .ZN(new_n515));
  AOI21_X1  g329(.A(G902), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT78), .B(G469), .ZN(new_n517));
  AOI22_X1  g331(.A1(G469), .A2(new_n508), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(G221), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n519), .B1(new_n449), .B2(new_n463), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n468), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n520), .ZN(new_n522));
  INV_X1    g336(.A(G469), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n498), .A2(new_n513), .A3(new_n514), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n471), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n498), .A2(new_n506), .A3(new_n472), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n523), .B1(new_n527), .B2(new_n463), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n511), .A2(new_n515), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n529), .A2(new_n463), .A3(new_n517), .ZN(new_n530));
  OAI211_X1 g344(.A(KEYINPUT79), .B(new_n522), .C1(new_n528), .C2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n467), .B1(new_n521), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT68), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT32), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n279), .B(new_n253), .C1(new_n482), .C2(new_n483), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT30), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n478), .A2(new_n323), .A3(new_n481), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n474), .A2(new_n476), .A3(new_n421), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n323), .B1(G134), .B2(G137), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n537), .B(new_n540), .C1(new_n261), .C2(new_n265), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n535), .A2(new_n536), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n536), .B1(new_n535), .B2(new_n541), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n198), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n535), .A2(new_n236), .A3(new_n541), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n306), .A2(G210), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(KEYINPUT27), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT26), .B(G101), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n547), .B(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n544), .A2(new_n545), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT31), .ZN(new_n551));
  INV_X1    g365(.A(new_n549), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n535), .A2(new_n236), .A3(new_n541), .ZN(new_n553));
  NOR2_X1   g367(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n541), .B1(new_n484), .B2(new_n258), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n198), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT67), .B1(new_n557), .B2(new_n545), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT28), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n552), .B(new_n555), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n551), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT31), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n544), .A2(new_n562), .A3(new_n545), .A4(new_n549), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT66), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n556), .A2(KEYINPUT30), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n535), .A2(new_n536), .A3(new_n541), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n553), .B1(new_n568), .B2(new_n198), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n569), .A2(KEYINPUT66), .A3(new_n562), .A4(new_n549), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n561), .B1(new_n565), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(G472), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n463), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n533), .B(new_n534), .C1(new_n571), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n570), .A2(new_n565), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT67), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n236), .B1(new_n535), .B2(new_n541), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n576), .B1(new_n553), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n578), .A2(KEYINPUT28), .B1(new_n553), .B2(new_n554), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n579), .A2(new_n552), .B1(new_n550), .B2(KEYINPUT31), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n573), .B1(new_n575), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT29), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n552), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT69), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n557), .A2(new_n584), .A3(new_n545), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n577), .A2(KEYINPUT69), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n559), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n545), .A2(KEYINPUT28), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n583), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n582), .B1(new_n569), .B2(new_n549), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n578), .A2(KEYINPUT28), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n552), .B1(new_n591), .B2(new_n555), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n589), .B(new_n463), .C1(new_n590), .C2(new_n592), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n581), .A2(KEYINPUT32), .B1(G472), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(KEYINPUT68), .B1(new_n581), .B2(KEYINPUT32), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n574), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n347), .A2(new_n348), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n190), .A2(G128), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n262), .A2(KEYINPUT23), .A3(G119), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n190), .A2(G128), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n598), .B(new_n599), .C1(new_n600), .C2(KEYINPUT23), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT24), .B(G110), .Z(new_n602));
  XNOR2_X1  g416(.A(G119), .B(G128), .ZN(new_n603));
  AOI22_X1  g417(.A1(new_n601), .A2(G110), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n597), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(KEYINPUT73), .B(G110), .ZN(new_n606));
  OAI22_X1  g420(.A1(new_n601), .A2(new_n606), .B1(new_n602), .B2(new_n603), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(new_n341), .A3(new_n318), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT22), .B(G137), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n519), .A2(new_n390), .A3(G953), .ZN(new_n611));
  XOR2_X1   g425(.A(new_n610), .B(new_n611), .Z(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n605), .A2(new_n608), .A3(new_n612), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n614), .A2(new_n463), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT25), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n450), .B1(G234), .B2(new_n463), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n614), .A2(new_n615), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n619), .A2(G902), .ZN(new_n621));
  AOI22_X1  g435(.A1(new_n618), .A2(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n596), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n532), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G101), .ZN(G3));
  NOR2_X1   g439(.A1(new_n571), .A2(G902), .ZN(new_n626));
  NAND2_X1  g440(.A1(KEYINPUT93), .A2(G472), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n575), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n463), .B1(new_n629), .B2(new_n561), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n630), .A2(KEYINPUT93), .A3(G472), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n628), .A2(new_n631), .A3(new_n622), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n521), .A2(new_n531), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT96), .B(G478), .Z(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n462), .B2(new_n463), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n460), .B1(new_n459), .B2(new_n428), .ZN(new_n637));
  INV_X1    g451(.A(new_n428), .ZN(new_n638));
  AOI211_X1 g452(.A(new_n638), .B(new_n452), .C1(new_n457), .C2(new_n458), .ZN(new_n639));
  OAI21_X1  g453(.A(KEYINPUT33), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT33), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n453), .A2(new_n461), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n398), .A2(G902), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n636), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n387), .A2(new_n645), .A3(new_n396), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT95), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n273), .A2(new_n299), .A3(new_n301), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n301), .B1(new_n273), .B2(new_n299), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT94), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n300), .A2(new_n650), .A3(new_n302), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n187), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n647), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n303), .A2(KEYINPUT94), .A3(new_n304), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n188), .B1(new_n649), .B2(new_n650), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n655), .A2(KEYINPUT95), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n646), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n634), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT34), .B(G104), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G6));
  NAND2_X1  g475(.A1(new_n462), .A2(new_n463), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n399), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n462), .A2(new_n463), .A3(new_n400), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n360), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n380), .A2(new_n385), .A3(new_n381), .A4(new_n382), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n384), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT97), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n384), .A2(KEYINPUT97), .A3(new_n668), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n667), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT98), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n673), .A2(new_n674), .A3(new_n397), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n655), .A2(KEYINPUT95), .A3(new_n656), .ZN(new_n676));
  AOI21_X1  g490(.A(KEYINPUT95), .B1(new_n655), .B2(new_n656), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n360), .B1(new_n663), .B2(new_n664), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n384), .A2(KEYINPUT97), .A3(new_n668), .ZN(new_n680));
  AOI21_X1  g494(.A(KEYINPUT97), .B1(new_n384), .B2(new_n668), .ZN(new_n681));
  OAI211_X1 g495(.A(new_n397), .B(new_n679), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(KEYINPUT98), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n675), .A2(new_n678), .A3(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n634), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT35), .B(G107), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G9));
  NAND2_X1  g501(.A1(new_n618), .A2(new_n619), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n613), .A2(KEYINPUT36), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n609), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n621), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n628), .A2(new_n631), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n532), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT37), .B(G110), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G12));
  AND3_X1   g510(.A1(new_n633), .A2(new_n596), .A3(new_n692), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT99), .B(G900), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n394), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n391), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n679), .B(new_n700), .C1(new_n680), .C2(new_n681), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n701), .A2(new_n676), .A3(new_n677), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G128), .ZN(G30));
  NOR2_X1   g518(.A1(new_n648), .A2(new_n649), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT38), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n384), .A2(new_n386), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n666), .ZN(new_n708));
  INV_X1    g522(.A(new_n692), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n708), .A2(new_n665), .A3(new_n709), .A4(new_n187), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n700), .B(KEYINPUT39), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n633), .A2(new_n711), .ZN(new_n712));
  AOI211_X1 g526(.A(new_n706), .B(new_n710), .C1(new_n712), .C2(KEYINPUT40), .ZN(new_n713));
  INV_X1    g527(.A(new_n569), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n549), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n585), .A2(new_n586), .ZN(new_n716));
  AOI21_X1  g530(.A(G902), .B1(new_n716), .B2(new_n552), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n572), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n718), .B1(new_n581), .B2(KEYINPUT32), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n574), .A2(new_n595), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(KEYINPUT100), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT100), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n574), .A2(new_n595), .A3(new_n719), .A4(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n713), .B(new_n724), .C1(KEYINPUT40), .C2(new_n712), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G143), .ZN(G45));
  INV_X1    g540(.A(KEYINPUT101), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n453), .A2(new_n461), .A3(new_n641), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n641), .B1(new_n453), .B2(new_n461), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n644), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n636), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n386), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n733), .B1(new_n383), .B2(KEYINPUT20), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n732), .B(new_n700), .C1(new_n360), .C2(new_n734), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n676), .A2(new_n735), .A3(new_n677), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n697), .A2(new_n727), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n633), .A2(new_n596), .A3(new_n692), .ZN(new_n738));
  INV_X1    g552(.A(new_n700), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n387), .A2(new_n645), .A3(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n654), .A3(new_n657), .ZN(new_n741));
  OAI21_X1  g555(.A(KEYINPUT101), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n737), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G146), .ZN(G48));
  INV_X1    g558(.A(new_n658), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n516), .A2(new_n523), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n516), .A2(new_n517), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n522), .A3(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n596), .A2(new_n622), .A3(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n745), .A2(new_n750), .A3(KEYINPUT102), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT102), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n596), .A2(new_n622), .A3(new_n749), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n752), .B1(new_n658), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(KEYINPUT41), .B(G113), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(G15));
  NAND4_X1  g571(.A1(new_n750), .A2(new_n675), .A3(new_n678), .A4(new_n683), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G116), .ZN(G18));
  NOR4_X1   g573(.A1(new_n665), .A2(new_n734), .A3(new_n360), .A4(new_n396), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n596), .A2(new_n760), .A3(new_n692), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n676), .A2(new_n677), .A3(new_n748), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G119), .ZN(G21));
  OAI21_X1  g578(.A(new_n665), .B1(new_n360), .B2(new_n734), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n676), .A2(new_n677), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n587), .A2(new_n588), .ZN(new_n767));
  AOI22_X1  g581(.A1(new_n767), .A2(new_n552), .B1(KEYINPUT31), .B2(new_n550), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n573), .B1(new_n768), .B2(new_n575), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n770), .B(new_n622), .C1(new_n626), .C2(new_n572), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n746), .A2(new_n522), .A3(new_n747), .A4(new_n397), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n766), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G122), .ZN(G24));
  AOI21_X1  g589(.A(new_n769), .B1(new_n630), .B2(G472), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n692), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n735), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n762), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G125), .ZN(G27));
  NAND2_X1  g594(.A1(G469), .A2(G902), .ZN(new_n781));
  XOR2_X1   g595(.A(new_n781), .B(KEYINPUT103), .Z(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n747), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT104), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n491), .B(new_n512), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n785), .B(new_n471), .C1(new_n786), .C2(new_n510), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n526), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n785), .B1(new_n524), .B2(new_n471), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n788), .A2(new_n523), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n522), .B1(new_n784), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n303), .A2(new_n187), .A3(new_n304), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n793), .A2(new_n596), .A3(new_n622), .A4(new_n740), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT42), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n791), .A2(new_n795), .A3(new_n792), .ZN(new_n797));
  OAI211_X1 g611(.A(KEYINPUT105), .B(new_n534), .C1(new_n571), .C2(new_n573), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT105), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n799), .B1(new_n581), .B2(KEYINPUT32), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n798), .A2(new_n594), .A3(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n797), .A2(new_n622), .A3(new_n740), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n796), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G131), .ZN(G33));
  NAND3_X1  g618(.A1(new_n673), .A2(KEYINPUT106), .A3(new_n700), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT106), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n701), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n805), .A2(new_n623), .A3(new_n793), .A4(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G134), .ZN(G36));
  NOR2_X1   g623(.A1(new_n708), .A2(new_n645), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT43), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n709), .B1(new_n628), .B2(new_n631), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(KEYINPUT44), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n792), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n815), .A2(KEYINPUT107), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(KEYINPUT107), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT44), .B1(new_n811), .B2(new_n812), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT45), .B1(new_n525), .B2(new_n526), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n788), .A2(new_n789), .ZN(new_n820));
  AOI211_X1 g634(.A(new_n523), .B(new_n819), .C1(new_n820), .C2(KEYINPUT45), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n782), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n822), .A2(KEYINPUT46), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n747), .B1(new_n822), .B2(KEYINPUT46), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n522), .B(new_n711), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n818), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n816), .A2(new_n817), .A3(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G137), .ZN(G39));
  OAI21_X1  g642(.A(new_n522), .B1(new_n823), .B2(new_n824), .ZN(new_n829));
  XNOR2_X1  g643(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n522), .B(new_n830), .C1(new_n823), .C2(new_n824), .ZN(new_n833));
  NOR4_X1   g647(.A1(new_n596), .A2(new_n735), .A3(new_n622), .A4(new_n792), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(G140), .ZN(G42));
  NAND3_X1  g650(.A1(new_n622), .A2(new_n522), .A3(new_n187), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n746), .A2(new_n747), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n837), .B1(KEYINPUT49), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n810), .ZN(new_n840));
  XOR2_X1   g654(.A(new_n840), .B(KEYINPUT109), .Z(new_n841));
  INV_X1    g655(.A(new_n724), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n838), .A2(KEYINPUT49), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT110), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n841), .A2(new_n842), .A3(new_n706), .A4(new_n844), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n762), .A2(new_n761), .B1(new_n766), .B2(new_n773), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT102), .B1(new_n745), .B2(new_n750), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n658), .A2(new_n753), .A3(new_n752), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n846), .B(new_n758), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT111), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT111), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n755), .A2(new_n851), .A3(new_n758), .A4(new_n846), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n803), .A2(new_n808), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n532), .B1(new_n623), .B2(new_n693), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n596), .A2(new_n692), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT112), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n680), .A2(new_n681), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n360), .A2(new_n739), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n705), .A2(new_n466), .A3(new_n187), .A4(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n856), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n671), .A2(new_n672), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n466), .A2(new_n858), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n861), .A2(KEYINPUT112), .A3(new_n814), .A4(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n855), .A2(new_n633), .A3(new_n860), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n387), .A2(new_n665), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n865), .B1(new_n387), .B2(new_n645), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n305), .A2(new_n397), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n632), .A2(new_n633), .A3(new_n866), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n778), .A2(new_n793), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n854), .A2(new_n864), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n853), .A2(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n850), .A2(new_n852), .A3(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n874));
  AOI22_X1  g688(.A1(new_n697), .A2(new_n702), .B1(new_n762), .B2(new_n778), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(KEYINPUT113), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n727), .B1(new_n697), .B2(new_n736), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n738), .A2(new_n741), .A3(KEYINPUT101), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n875), .A2(KEYINPUT113), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n791), .A2(new_n692), .A3(new_n739), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n724), .A2(new_n766), .A3(new_n882), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n883), .A2(KEYINPUT52), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n880), .A2(new_n881), .A3(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  XOR2_X1   g700(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n887));
  INV_X1    g701(.A(KEYINPUT114), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n883), .A2(new_n703), .A3(new_n779), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n888), .B1(new_n879), .B2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n743), .A2(KEYINPUT114), .A3(new_n875), .A4(new_n883), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n887), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n873), .B(new_n874), .C1(new_n886), .C2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT52), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n890), .A2(new_n894), .A3(new_n891), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n894), .B1(new_n890), .B2(new_n891), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n850), .A2(new_n872), .A3(new_n852), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n893), .B(KEYINPUT54), .C1(new_n898), .C2(new_n874), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT54), .ZN(new_n900));
  NOR4_X1   g714(.A1(new_n849), .A2(new_n853), .A3(new_n871), .A4(new_n874), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n901), .B1(new_n886), .B2(new_n892), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n900), .B(new_n902), .C1(new_n898), .C2(KEYINPUT53), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n811), .A2(new_n392), .ZN(new_n904));
  INV_X1    g718(.A(new_n771), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n904), .A2(new_n762), .A3(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n748), .A2(new_n792), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n907), .A2(new_n622), .A3(new_n392), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n842), .A2(new_n708), .A3(new_n732), .A4(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n906), .A2(new_n389), .A3(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT48), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n801), .A2(new_n622), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n904), .A2(new_n911), .A3(new_n913), .A4(new_n907), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n904), .A2(new_n913), .A3(new_n907), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(KEYINPUT48), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n910), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n777), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n904), .A2(new_n918), .A3(new_n907), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n842), .A2(new_n387), .A3(new_n645), .A4(new_n908), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n706), .A2(new_n188), .A3(new_n749), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n904), .A2(KEYINPUT50), .A3(new_n905), .A4(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT50), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n811), .A2(new_n392), .A3(new_n905), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n925), .B1(new_n926), .B2(new_n922), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n921), .A2(KEYINPUT51), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n746), .A2(new_n520), .A3(new_n747), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n931), .B1(new_n832), .B2(new_n833), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n904), .A2(new_n905), .A3(new_n814), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n917), .B1(new_n929), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT117), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n924), .A2(new_n936), .A3(new_n927), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n921), .A2(new_n937), .ZN(new_n938));
  OR3_X1    g752(.A1(new_n932), .A2(KEYINPUT116), .A3(new_n933), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n928), .A2(KEYINPUT117), .ZN(new_n940));
  OAI21_X1  g754(.A(KEYINPUT116), .B1(new_n932), .B2(new_n933), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n938), .A2(new_n939), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT51), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n935), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n899), .A2(new_n903), .A3(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT118), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n388), .A2(new_n325), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT119), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(new_n945), .B2(new_n946), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n845), .B1(new_n947), .B2(new_n950), .ZN(G75));
  NOR2_X1   g765(.A1(new_n325), .A2(G952), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n883), .A2(new_n703), .A3(new_n779), .ZN(new_n954));
  AOI21_X1  g768(.A(KEYINPUT114), .B1(new_n954), .B2(new_n743), .ZN(new_n955));
  INV_X1    g769(.A(new_n891), .ZN(new_n956));
  OAI21_X1  g770(.A(KEYINPUT52), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n890), .A2(new_n894), .A3(new_n891), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n957), .A2(new_n873), .A3(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n887), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(new_n955), .B2(new_n956), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n885), .ZN(new_n962));
  AOI22_X1  g776(.A1(new_n959), .A2(new_n874), .B1(new_n962), .B2(new_n901), .ZN(new_n963));
  INV_X1    g777(.A(G210), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n963), .A2(new_n964), .A3(new_n463), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n242), .A2(new_n244), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(new_n272), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT55), .Z(new_n968));
  OR2_X1    g782(.A1(new_n968), .A2(KEYINPUT56), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n953), .B1(new_n965), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n902), .B1(new_n898), .B2(KEYINPUT53), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n971), .A2(G210), .A3(G902), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(KEYINPUT120), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT56), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT120), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n971), .A2(new_n975), .A3(G210), .A4(G902), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n973), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n970), .B1(new_n977), .B2(new_n968), .ZN(G51));
  XNOR2_X1  g792(.A(new_n782), .B(KEYINPUT57), .ZN(new_n979));
  INV_X1    g793(.A(new_n903), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n959), .A2(new_n874), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n900), .B1(new_n981), .B2(new_n902), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n979), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n529), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n971), .A2(G902), .A3(new_n821), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n952), .B1(new_n984), .B2(new_n985), .ZN(G54));
  NAND2_X1  g800(.A1(KEYINPUT58), .A2(G475), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT121), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n971), .A2(G902), .A3(new_n988), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n380), .A2(new_n382), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n953), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n989), .A2(new_n991), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(KEYINPUT122), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT122), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n989), .A2(new_n995), .A3(new_n991), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n992), .B1(new_n994), .B2(new_n996), .ZN(G60));
  NAND2_X1  g811(.A1(new_n899), .A2(new_n903), .ZN(new_n998));
  NAND2_X1  g812(.A1(G478), .A2(G902), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT59), .Z(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n643), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n643), .A2(new_n1001), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n971), .A2(KEYINPUT54), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1003), .B1(new_n1004), .B2(new_n903), .ZN(new_n1005));
  NOR3_X1   g819(.A1(new_n1002), .A2(new_n1005), .A3(new_n952), .ZN(G63));
  INV_X1    g820(.A(new_n620), .ZN(new_n1007));
  XNOR2_X1  g821(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n1008));
  NAND2_X1  g822(.A1(G217), .A2(G902), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1008), .B(new_n1009), .Z(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1007), .B1(new_n963), .B2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n971), .A2(new_n690), .A3(new_n1010), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1012), .A2(new_n953), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT61), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n1012), .A2(new_n1013), .A3(KEYINPUT61), .A4(new_n953), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(new_n1017), .ZN(G66));
  NAND4_X1  g832(.A1(new_n850), .A2(new_n852), .A3(new_n869), .A4(new_n854), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n325), .ZN(new_n1020));
  OAI21_X1  g834(.A(G953), .B1(new_n395), .B2(new_n270), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n966), .B1(G898), .B2(new_n325), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(KEYINPUT124), .Z(new_n1024));
  XNOR2_X1  g838(.A(new_n1022), .B(new_n1024), .ZN(G69));
  INV_X1    g839(.A(new_n825), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1026), .A2(new_n766), .A3(new_n913), .ZN(new_n1027));
  AND4_X1   g841(.A1(new_n803), .A2(new_n1027), .A3(new_n835), .A4(new_n808), .ZN(new_n1028));
  AND2_X1   g842(.A1(new_n880), .A2(new_n881), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n827), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  OR2_X1    g844(.A1(new_n1030), .A2(G953), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n568), .B(KEYINPUT125), .Z(new_n1032));
  XNOR2_X1  g846(.A(new_n1032), .B(new_n364), .ZN(new_n1033));
  INV_X1    g847(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1034), .B1(G900), .B2(G953), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n325), .B1(G227), .B2(G900), .ZN(new_n1036));
  AOI22_X1  g850(.A1(new_n1031), .A2(new_n1035), .B1(KEYINPUT127), .B2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g851(.A1(new_n1036), .A2(KEYINPUT127), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1029), .A2(new_n725), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1040), .A2(KEYINPUT62), .ZN(new_n1041));
  INV_X1    g855(.A(KEYINPUT62), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n1029), .A2(new_n1042), .A3(new_n725), .ZN(new_n1043));
  NOR2_X1   g857(.A1(new_n712), .A2(new_n792), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n1044), .A2(new_n623), .A3(new_n866), .ZN(new_n1045));
  AND2_X1   g859(.A1(new_n835), .A2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g860(.A1(new_n1041), .A2(new_n827), .A3(new_n1043), .A4(new_n1046), .ZN(new_n1047));
  AND2_X1   g861(.A1(new_n1047), .A2(new_n325), .ZN(new_n1048));
  XNOR2_X1  g862(.A(new_n1033), .B(KEYINPUT126), .ZN(new_n1049));
  OAI211_X1 g863(.A(new_n1037), .B(new_n1039), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  INV_X1    g864(.A(KEYINPUT127), .ZN(new_n1051));
  INV_X1    g865(.A(new_n1036), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n1049), .B1(new_n1047), .B2(new_n325), .ZN(new_n1053));
  NOR2_X1   g867(.A1(new_n1030), .A2(G953), .ZN(new_n1054));
  INV_X1    g868(.A(new_n1035), .ZN(new_n1055));
  NOR2_X1   g869(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g870(.A(new_n1051), .B(new_n1052), .C1(new_n1053), .C2(new_n1056), .ZN(new_n1057));
  AND2_X1   g871(.A1(new_n1050), .A2(new_n1057), .ZN(G72));
  NAND2_X1  g872(.A1(G472), .A2(G902), .ZN(new_n1059));
  XOR2_X1   g873(.A(new_n1059), .B(KEYINPUT63), .Z(new_n1060));
  OAI21_X1  g874(.A(new_n1060), .B1(new_n1047), .B2(new_n1019), .ZN(new_n1061));
  NAND3_X1  g875(.A1(new_n1061), .A2(new_n714), .A3(new_n549), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n715), .A2(new_n1060), .ZN(new_n1063));
  NOR2_X1   g877(.A1(new_n714), .A2(new_n549), .ZN(new_n1064));
  NOR2_X1   g878(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g879(.A(new_n893), .B(new_n1065), .C1(new_n898), .C2(new_n874), .ZN(new_n1066));
  OAI21_X1  g880(.A(new_n1060), .B1(new_n1030), .B2(new_n1019), .ZN(new_n1067));
  AOI21_X1  g881(.A(new_n952), .B1(new_n1067), .B2(new_n1064), .ZN(new_n1068));
  AND3_X1   g882(.A1(new_n1062), .A2(new_n1066), .A3(new_n1068), .ZN(G57));
endmodule


