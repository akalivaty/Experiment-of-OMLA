//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 1 1 1 1 1 0 1 0 0 0 1 0 0 0 0 1 0 1 1 0 0 1 1 1 1 0 1 0 0 0 0 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n448, new_n450, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n571, new_n572,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n601, new_n602, new_n603,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n637,
    new_n638, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1222, new_n1223, new_n1224;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT66), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  NAND2_X1  g022(.A1(G94), .A2(G452), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT67), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n455), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OR2_X1    g036(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  XNOR2_X1  g041(.A(new_n466), .B(KEYINPUT69), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND3_X1  g043(.A1(KEYINPUT68), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(KEYINPUT3), .B1(KEYINPUT68), .B2(G2104), .ZN(new_n471));
  OR2_X1    g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(G137), .A3(new_n465), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n475), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(new_n465), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n474), .A2(new_n477), .ZN(G160));
  OR3_X1    g053(.A1(new_n470), .A2(KEYINPUT70), .A3(new_n471), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n472), .A2(KEYINPUT70), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n479), .A2(new_n465), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  AND3_X1   g058(.A1(new_n479), .A2(G2105), .A3(new_n480), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  OAI211_X1 g064(.A(G138), .B(new_n465), .C1(new_n470), .C2(new_n471), .ZN(new_n490));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR3_X1   g066(.A1(new_n491), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n492));
  AOI22_X1  g067(.A1(new_n490), .A2(KEYINPUT4), .B1(new_n475), .B2(new_n492), .ZN(new_n493));
  AND2_X1   g068(.A1(G126), .A2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n494), .B1(new_n470), .B2(new_n471), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT71), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G114), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n465), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n495), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n493), .A2(new_n502), .ZN(G164));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n504), .A2(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(G543), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n504), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OR2_X1    g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n504), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G50), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n510), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n513), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  NAND2_X1  g098(.A1(new_n508), .A2(new_n509), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n507), .A2(G543), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n524), .A2(G89), .A3(new_n525), .A4(new_n518), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(KEYINPUT74), .A2(KEYINPUT7), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(KEYINPUT74), .A2(KEYINPUT7), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n531), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n533), .A2(new_n527), .A3(new_n529), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n526), .A2(new_n535), .ZN(new_n536));
  AND2_X1   g111(.A1(G63), .A2(G651), .ZN(new_n537));
  AND3_X1   g112(.A1(new_n504), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n538));
  AOI21_X1  g113(.A(KEYINPUT72), .B1(new_n504), .B2(KEYINPUT5), .ZN(new_n539));
  OAI211_X1 g114(.A(new_n525), .B(new_n537), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n518), .A2(G51), .A3(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(KEYINPUT73), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n540), .A2(new_n544), .A3(new_n541), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n536), .B1(new_n543), .B2(new_n545), .ZN(G168));
  OAI211_X1 g121(.A(G64), .B(new_n525), .C1(new_n538), .C2(new_n539), .ZN(new_n547));
  NAND2_X1  g122(.A1(G77), .A2(G543), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n512), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g124(.A1(KEYINPUT75), .A2(G90), .ZN(new_n550));
  NOR2_X1   g125(.A1(KEYINPUT75), .A2(G90), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n524), .A2(new_n525), .A3(new_n518), .A4(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n516), .A2(G52), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n549), .A2(new_n555), .ZN(G171));
  AND2_X1   g131(.A1(new_n510), .A2(new_n518), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n557), .A2(G81), .B1(G43), .B2(new_n516), .ZN(new_n558));
  NAND2_X1  g133(.A1(G68), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n560), .B1(new_n510), .B2(G56), .ZN(new_n561));
  OAI21_X1  g136(.A(G651), .B1(new_n561), .B2(KEYINPUT76), .ZN(new_n562));
  OAI211_X1 g137(.A(G56), .B(new_n525), .C1(new_n538), .C2(new_n539), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n563), .A2(KEYINPUT76), .A3(new_n559), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n558), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT77), .ZN(G153));
  NAND4_X1  g144(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND4_X1  g147(.A1(G319), .A2(G483), .A3(G661), .A4(new_n572), .ZN(G188));
  AND2_X1   g148(.A1(KEYINPUT6), .A2(G651), .ZN(new_n574));
  NOR2_X1   g149(.A1(KEYINPUT6), .A2(G651), .ZN(new_n575));
  OAI211_X1 g150(.A(G53), .B(G543), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT9), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT9), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n516), .A2(new_n578), .A3(G53), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n557), .A2(G91), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n524), .A2(G65), .A3(new_n525), .ZN(new_n581));
  NAND2_X1  g156(.A1(G78), .A2(G543), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n512), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g159(.A(KEYINPUT78), .B1(new_n580), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n510), .A2(G91), .A3(new_n518), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n578), .B1(new_n516), .B2(G53), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n576), .A2(KEYINPUT9), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT78), .ZN(new_n590));
  NOR3_X1   g165(.A1(new_n589), .A2(new_n583), .A3(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n585), .A2(new_n591), .ZN(G299));
  NAND2_X1  g167(.A1(new_n547), .A2(new_n548), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G651), .ZN(new_n594));
  AND2_X1   g169(.A1(new_n553), .A2(new_n554), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n594), .A2(new_n595), .A3(KEYINPUT79), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT79), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(new_n549), .B2(new_n555), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G301));
  AND2_X1   g175(.A1(new_n526), .A2(new_n535), .ZN(new_n601));
  AND3_X1   g176(.A1(new_n540), .A2(new_n544), .A3(new_n541), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n544), .B1(new_n540), .B2(new_n541), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(G286));
  NAND2_X1  g179(.A1(new_n516), .A2(G49), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT80), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n557), .A2(G87), .ZN(new_n607));
  OAI21_X1  g182(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(G288));
  AOI22_X1  g184(.A1(new_n510), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n610), .A2(new_n512), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n516), .A2(G48), .ZN(new_n612));
  INV_X1    g187(.A(G86), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n519), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(G305));
  AOI22_X1  g191(.A1(new_n557), .A2(G85), .B1(G47), .B2(new_n516), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n512), .B2(new_n618), .ZN(G290));
  NAND2_X1  g194(.A1(new_n510), .A2(G66), .ZN(new_n620));
  NAND2_X1  g195(.A1(G79), .A2(G543), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n518), .A2(G543), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n623), .A2(KEYINPUT81), .ZN(new_n624));
  INV_X1    g199(.A(G54), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n625), .B1(new_n623), .B2(KEYINPUT81), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n622), .A2(G651), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT10), .ZN(new_n628));
  INV_X1    g203(.A(G92), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n519), .B2(new_n629), .ZN(new_n630));
  NAND4_X1  g205(.A1(new_n510), .A2(KEYINPUT10), .A3(G92), .A4(new_n518), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n633), .A2(G868), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n634), .B1(G868), .B2(new_n599), .ZN(G284));
  AOI21_X1  g210(.A(new_n634), .B1(G868), .B2(new_n599), .ZN(G321));
  NAND2_X1  g211(.A1(G286), .A2(G868), .ZN(new_n637));
  INV_X1    g212(.A(G299), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(G868), .ZN(G297));
  OAI21_X1  g214(.A(new_n637), .B1(new_n638), .B2(G868), .ZN(G280));
  INV_X1    g215(.A(new_n633), .ZN(new_n641));
  INV_X1    g216(.A(G559), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n641), .B1(new_n642), .B2(G860), .ZN(G148));
  INV_X1    g218(.A(G868), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n566), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n633), .A2(G559), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n645), .B1(new_n646), .B2(new_n644), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT82), .Z(G323));
  XNOR2_X1  g223(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g224(.A1(new_n482), .A2(G135), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT84), .Z(new_n651));
  NAND2_X1  g226(.A1(new_n484), .A2(G123), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT85), .Z(new_n653));
  OR2_X1    g228(.A1(G99), .A2(G2105), .ZN(new_n654));
  OAI211_X1 g229(.A(new_n654), .B(G2104), .C1(G111), .C2(new_n465), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n651), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n656), .A2(G2096), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n467), .A2(new_n475), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT12), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT13), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n660), .B1(KEYINPUT83), .B2(G2100), .ZN(new_n661));
  NAND2_X1  g236(.A1(KEYINPUT83), .A2(G2100), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n656), .A2(G2096), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n660), .A2(KEYINPUT83), .A3(G2100), .ZN(new_n665));
  NAND4_X1  g240(.A1(new_n657), .A2(new_n663), .A3(new_n664), .A4(new_n665), .ZN(G156));
  XNOR2_X1  g241(.A(G2427), .B(G2438), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2430), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT15), .B(G2435), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(KEYINPUT14), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2451), .B(G2454), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT16), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n672), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2443), .B(G2446), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1341), .B(G1348), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT86), .ZN(new_n680));
  OAI21_X1  g255(.A(G14), .B1(new_n677), .B2(new_n678), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(G401));
  XOR2_X1   g257(.A(G2084), .B(G2090), .Z(new_n683));
  XNOR2_X1  g258(.A(G2067), .B(G2678), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT87), .Z(new_n685));
  NOR2_X1   g260(.A1(G2072), .A2(G2078), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n444), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n683), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(KEYINPUT17), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n688), .B1(new_n685), .B2(new_n689), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n683), .B(new_n684), .C1(new_n444), .C2(new_n686), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT18), .Z(new_n692));
  NAND3_X1  g267(.A1(new_n689), .A2(new_n685), .A3(new_n683), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n690), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G2096), .B(G2100), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(G227));
  XOR2_X1   g271(.A(G1971), .B(G1976), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT19), .ZN(new_n698));
  XOR2_X1   g273(.A(G1956), .B(G2474), .Z(new_n699));
  XOR2_X1   g274(.A(G1961), .B(G1966), .Z(new_n700));
  AND2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT20), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n699), .A2(new_n700), .ZN(new_n704));
  NOR3_X1   g279(.A1(new_n698), .A2(new_n701), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n698), .B2(new_n704), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(G1991), .B(G1996), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(G1981), .B(G1986), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(G229));
  INV_X1    g288(.A(KEYINPUT90), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT88), .B(G16), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n715), .A2(G24), .ZN(new_n716));
  INV_X1    g291(.A(new_n715), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n716), .B1(G290), .B2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G1986), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n714), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(G25), .A2(G29), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n482), .A2(G131), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n484), .A2(G119), .ZN(new_n723));
  OR2_X1    g298(.A1(G95), .A2(G2105), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n724), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n721), .B1(new_n727), .B2(G29), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT35), .B(G1991), .Z(new_n729));
  XOR2_X1   g304(.A(new_n728), .B(new_n729), .Z(new_n730));
  AOI211_X1 g305(.A(new_n720), .B(new_n730), .C1(new_n719), .C2(new_n718), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n717), .A2(G22), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G166), .B2(new_n717), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(G1971), .Z(new_n734));
  INV_X1    g309(.A(G288), .ZN(new_n735));
  INV_X1    g310(.A(G16), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n736), .B2(G23), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT33), .B(G1976), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n615), .A2(G16), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G6), .B2(G16), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT32), .B(G1981), .Z(new_n743));
  AOI22_X1  g318(.A1(new_n738), .A2(new_n739), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n734), .A2(new_n740), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n746), .A2(KEYINPUT89), .A3(KEYINPUT34), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(KEYINPUT89), .B1(new_n746), .B2(KEYINPUT34), .ZN(new_n749));
  OAI221_X1 g324(.A(new_n731), .B1(KEYINPUT34), .B2(new_n746), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT36), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  INV_X1    g328(.A(G29), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G35), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G162), .B2(new_n754), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT29), .Z(new_n757));
  INV_X1    g332(.A(G2090), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT99), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n736), .A2(G21), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G168), .B2(new_n736), .ZN(new_n762));
  INV_X1    g337(.A(G1966), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n754), .A2(G27), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT97), .Z(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G164), .B2(new_n754), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(new_n443), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT98), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n764), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n754), .A2(G26), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT28), .Z(new_n772));
  NAND2_X1  g347(.A1(new_n482), .A2(G140), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n484), .A2(G128), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n465), .A2(G116), .ZN(new_n775));
  OAI21_X1  g350(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n773), .B(new_n774), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n772), .B1(new_n777), .B2(G29), .ZN(new_n778));
  INV_X1    g353(.A(G2067), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  AOI211_X1 g355(.A(new_n770), .B(new_n780), .C1(new_n769), .C2(new_n768), .ZN(new_n781));
  NAND2_X1  g356(.A1(G160), .A2(G29), .ZN(new_n782));
  INV_X1    g357(.A(G34), .ZN(new_n783));
  AOI21_X1  g358(.A(G29), .B1(new_n783), .B2(KEYINPUT24), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n784), .A2(KEYINPUT93), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(KEYINPUT93), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(KEYINPUT24), .B2(new_n783), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n782), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(G2084), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n736), .A2(G5), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G171), .B2(new_n736), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n754), .A2(G32), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n482), .A2(G141), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n484), .A2(G129), .ZN(new_n795));
  NAND3_X1  g370(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT26), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n467), .A2(G105), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n794), .A2(new_n795), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n793), .B1(new_n801), .B2(G29), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT27), .B(G1996), .ZN(new_n803));
  OAI221_X1 g378(.A(new_n790), .B1(G1961), .B2(new_n792), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT96), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n802), .A2(new_n803), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n656), .B2(new_n754), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n788), .A2(new_n789), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT31), .B(G11), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT94), .B(G28), .Z(new_n811));
  AOI21_X1  g386(.A(G29), .B1(new_n811), .B2(KEYINPUT30), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT95), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(KEYINPUT30), .B2(new_n811), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n812), .A2(new_n813), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n810), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n809), .A2(new_n817), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n754), .A2(G33), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT25), .Z(new_n821));
  AOI22_X1  g396(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n822));
  INV_X1    g397(.A(G139), .ZN(new_n823));
  OAI221_X1 g398(.A(new_n821), .B1(new_n465), .B2(new_n822), .C1(new_n481), .C2(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n819), .B1(new_n824), .B2(G29), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n825), .A2(new_n442), .B1(G1961), .B2(new_n792), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n818), .B(new_n826), .C1(new_n442), .C2(new_n825), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n806), .A2(new_n808), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(G4), .A2(G16), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT91), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n633), .B2(new_n736), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT92), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(G1348), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n781), .A2(new_n828), .A3(new_n833), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n757), .A2(new_n758), .B1(new_n804), .B2(new_n805), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n717), .A2(G19), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(new_n567), .B2(new_n717), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(G1341), .Z(new_n838));
  NAND2_X1  g413(.A1(new_n715), .A2(G20), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT23), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n638), .B2(new_n736), .ZN(new_n841));
  INV_X1    g416(.A(G1956), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n835), .A2(new_n838), .A3(new_n843), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n760), .A2(new_n834), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n752), .A2(new_n753), .A3(new_n845), .ZN(G150));
  INV_X1    g421(.A(G150), .ZN(G311));
  INV_X1    g422(.A(KEYINPUT101), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n524), .A2(G67), .A3(new_n525), .ZN(new_n849));
  NAND2_X1  g424(.A1(G80), .A2(G543), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(G651), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n524), .A2(G93), .A3(new_n525), .A4(new_n518), .ZN(new_n853));
  XNOR2_X1  g428(.A(KEYINPUT100), .B(G55), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n516), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n848), .B1(new_n852), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n512), .B1(new_n849), .B2(new_n850), .ZN(new_n859));
  NOR3_X1   g434(.A1(new_n859), .A2(new_n856), .A3(KEYINPUT101), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n566), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n563), .A2(new_n559), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT76), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n864), .A2(G651), .A3(new_n564), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n859), .A2(new_n856), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(new_n558), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n861), .A2(new_n867), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT38), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n641), .A2(G559), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n871), .A2(KEYINPUT39), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(KEYINPUT39), .ZN(new_n873));
  NOR3_X1   g448(.A1(new_n872), .A2(new_n873), .A3(G860), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n852), .A2(new_n857), .A3(new_n848), .ZN(new_n875));
  OAI21_X1  g450(.A(KEYINPUT101), .B1(new_n859), .B2(new_n856), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(G860), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT37), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n874), .A2(new_n879), .ZN(G145));
  INV_X1    g455(.A(new_n493), .ZN(new_n881));
  INV_X1    g456(.A(new_n501), .ZN(new_n882));
  XNOR2_X1  g457(.A(KEYINPUT71), .B(G114), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n882), .B1(new_n883), .B2(new_n465), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n885), .A3(new_n495), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n885), .B1(new_n884), .B2(new_n495), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n881), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT103), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n502), .A2(KEYINPUT102), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n493), .B1(new_n892), .B2(new_n886), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT103), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n777), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n727), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n482), .A2(G142), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n484), .A2(G130), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n465), .A2(G118), .ZN(new_n900));
  OAI21_X1  g475(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n898), .B(new_n899), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(new_n659), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n801), .B(new_n824), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n903), .B(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n897), .B(new_n905), .ZN(new_n906));
  XOR2_X1   g481(.A(new_n488), .B(G160), .Z(new_n907));
  XNOR2_X1  g482(.A(new_n656), .B(new_n907), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n906), .A2(new_n908), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n909), .A2(new_n910), .A3(G37), .ZN(new_n911));
  XNOR2_X1  g486(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n911), .B(new_n912), .ZN(G395));
  NAND2_X1  g488(.A1(new_n877), .A2(new_n644), .ZN(new_n914));
  XNOR2_X1  g489(.A(G305), .B(G288), .ZN(new_n915));
  XNOR2_X1  g490(.A(G303), .B(G290), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n915), .B(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n917), .A2(KEYINPUT42), .ZN(new_n918));
  XOR2_X1   g493(.A(new_n918), .B(KEYINPUT107), .Z(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(KEYINPUT42), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(KEYINPUT106), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n868), .B(new_n646), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n633), .B1(new_n585), .B2(new_n591), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n580), .A2(new_n584), .A3(KEYINPUT78), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n590), .B1(new_n589), .B2(new_n583), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n925), .A2(new_n926), .A3(new_n632), .A4(new_n627), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n923), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT41), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n924), .A2(new_n927), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n930), .B1(new_n923), .B2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n922), .B(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n914), .B1(new_n938), .B2(new_n644), .ZN(G295));
  OAI21_X1  g514(.A(new_n914), .B1(new_n938), .B2(new_n644), .ZN(G331));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n941));
  XNOR2_X1  g516(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n942));
  AOI22_X1  g517(.A1(new_n875), .A2(new_n876), .B1(new_n865), .B2(new_n558), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n865), .A2(new_n558), .A3(new_n866), .ZN(new_n944));
  AOI21_X1  g519(.A(G286), .B1(new_n598), .B2(new_n596), .ZN(new_n945));
  NOR2_X1   g520(.A1(G168), .A2(G171), .ZN(new_n946));
  OAI22_X1  g521(.A1(new_n943), .A2(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT79), .B1(new_n594), .B2(new_n595), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n549), .A2(new_n555), .A3(new_n597), .ZN(new_n949));
  OAI21_X1  g524(.A(G168), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(G286), .B1(new_n549), .B2(new_n555), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n861), .A2(new_n950), .A3(new_n867), .A4(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n947), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n868), .B(KEYINPUT110), .C1(new_n945), .C2(new_n946), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n928), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n945), .A2(new_n946), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n958), .A2(new_n959), .A3(new_n861), .A4(new_n867), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n947), .A2(new_n952), .A3(KEYINPUT109), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n936), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n957), .A2(new_n917), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G37), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n917), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n936), .A2(new_n960), .A3(new_n961), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n929), .B1(new_n954), .B2(new_n955), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n942), .B1(new_n966), .B2(new_n970), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n924), .A2(new_n931), .A3(new_n927), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n933), .B1(new_n924), .B2(new_n927), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n974), .A2(new_n955), .A3(new_n954), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n929), .B1(new_n961), .B2(new_n960), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n967), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n977), .A2(new_n964), .A3(new_n963), .ZN(new_n978));
  INV_X1    g553(.A(new_n942), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n941), .B1(new_n971), .B2(new_n980), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n978), .A2(KEYINPUT112), .A3(KEYINPUT43), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT112), .B1(new_n978), .B2(KEYINPUT43), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT44), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n970), .A2(new_n964), .A3(new_n963), .A4(new_n942), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n986), .B(new_n987), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n984), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n976), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n974), .A2(new_n955), .A3(new_n954), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n917), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT43), .B1(new_n965), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n978), .A2(KEYINPUT112), .A3(KEYINPUT43), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n941), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n986), .B(KEYINPUT111), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT113), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n981), .B1(new_n989), .B2(new_n999), .ZN(G397));
  INV_X1    g575(.A(G40), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n474), .A2(new_n1001), .A3(new_n477), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  XOR2_X1   g578(.A(KEYINPUT115), .B(KEYINPUT45), .Z(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1384), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n895), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT114), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT114), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n895), .A2(new_n1009), .A3(new_n1006), .ZN(new_n1010));
  AOI211_X1 g585(.A(new_n1003), .B(new_n1005), .C1(new_n1008), .C2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n777), .B(new_n779), .ZN(new_n1012));
  INV_X1    g587(.A(G1996), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n801), .B(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n727), .A2(new_n729), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n727), .A2(new_n729), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(G290), .B(G1986), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1011), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G164), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1020), .A2(new_n1006), .A3(new_n1005), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n892), .A2(new_n886), .ZN(new_n1022));
  AOI21_X1  g597(.A(G1384), .B1(new_n1022), .B2(new_n881), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1021), .B(new_n1002), .C1(new_n1023), .C2(KEYINPUT45), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n763), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1026), .B1(new_n893), .B2(G1384), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1020), .A2(KEYINPUT50), .A3(new_n1006), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1003), .A2(G2084), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1025), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1032), .A2(G8), .A3(G286), .ZN(new_n1033));
  NAND2_X1  g608(.A1(G286), .A2(G8), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1034), .B(KEYINPUT123), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n1024), .A2(new_n763), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1036));
  INV_X1    g611(.A(G8), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1035), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1033), .A2(new_n1038), .A3(KEYINPUT51), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT124), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT51), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1041), .B(new_n1034), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n1039), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1040), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT62), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1037), .B1(new_n1025), .B2(new_n1031), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1035), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT51), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n1036), .A2(new_n1037), .A3(G168), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1042), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT124), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT62), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1039), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(G303), .A2(G8), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n1055), .B(KEYINPUT55), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1006), .A2(KEYINPUT45), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n891), .A2(new_n894), .A3(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1004), .B1(G164), .B2(G1384), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1058), .A2(new_n1002), .A3(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT116), .B(G1971), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1026), .B(new_n1006), .C1(new_n493), .C2(new_n502), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1002), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n889), .A2(new_n1006), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1064), .B1(KEYINPUT50), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n758), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1062), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1060), .A2(new_n1061), .B1(new_n1066), .B2(new_n758), .ZN(new_n1071));
  OAI21_X1  g646(.A(G8), .B1(new_n1071), .B2(KEYINPUT117), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1056), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1003), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n758), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1037), .B1(new_n1062), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1056), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1079), .B1(new_n1060), .B2(G2078), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n1074), .A2(G1961), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OR3_X1    g657(.A1(new_n1024), .A2(new_n1079), .A3(G2078), .ZN(new_n1083));
  AOI21_X1  g658(.A(G301), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT49), .ZN(new_n1085));
  INV_X1    g660(.A(G1981), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n615), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n615), .A2(new_n1086), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1085), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1089), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1091), .A2(KEYINPUT49), .A3(new_n1087), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1037), .B1(new_n1023), .B2(new_n1002), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1090), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(G1976), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT52), .B1(G288), .B2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1093), .B(new_n1096), .C1(new_n1095), .C2(G288), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1093), .ZN(new_n1098));
  NOR2_X1   g673(.A1(G288), .A2(new_n1095), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT52), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1094), .A2(new_n1097), .A3(new_n1100), .ZN(new_n1101));
  AND4_X1   g676(.A1(new_n1073), .A2(new_n1078), .A3(new_n1084), .A4(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1045), .A2(new_n1054), .A3(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1094), .A2(new_n1095), .A3(new_n735), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1098), .B1(new_n1104), .B2(new_n1087), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1078), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1105), .B1(new_n1106), .B2(new_n1101), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1003), .A2(G1996), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1058), .A2(new_n1108), .A3(new_n1059), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1023), .A2(new_n1002), .ZN(new_n1110));
  XOR2_X1   g685(.A(KEYINPUT58), .B(G1341), .Z(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n567), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT120), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1113), .A2(new_n1117), .A3(new_n567), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1115), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1117), .B1(new_n1113), .B2(new_n567), .ZN(new_n1120));
  AOI211_X1 g695(.A(KEYINPUT120), .B(new_n566), .C1(new_n1109), .C2(new_n1112), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT59), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT56), .B(G2072), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1058), .A2(new_n1002), .A3(new_n1059), .A4(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n842), .B1(new_n1126), .B2(new_n1064), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n580), .A2(new_n584), .ZN(new_n1129));
  XOR2_X1   g704(.A(new_n1129), .B(KEYINPUT57), .Z(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1125), .A2(new_n1127), .A3(new_n1130), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1130), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT61), .B1(new_n1136), .B2(KEYINPUT121), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT61), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1135), .A2(new_n1137), .B1(new_n1139), .B2(new_n1134), .ZN(new_n1140));
  OAI22_X1  g715(.A1(new_n1074), .A2(G1348), .B1(G2067), .B2(new_n1110), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT60), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n641), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(KEYINPUT122), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1110), .A2(G2067), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1029), .A2(new_n1002), .ZN(new_n1147));
  INV_X1    g722(.A(G1348), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(KEYINPUT60), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT122), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1143), .A2(new_n1152), .A3(new_n641), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1145), .A2(new_n1151), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1152), .B1(new_n1143), .B2(new_n641), .ZN(new_n1155));
  AOI211_X1 g730(.A(KEYINPUT122), .B(new_n633), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1150), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1123), .A2(new_n1140), .A3(new_n1154), .A4(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1149), .A2(new_n633), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1134), .B1(new_n1159), .B2(new_n1136), .ZN(new_n1160));
  AND2_X1   g735(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1078), .A2(new_n1101), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1163), .B1(new_n1164), .B2(new_n1056), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT54), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n443), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1167));
  INV_X1    g742(.A(new_n476), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n1168), .A2(KEYINPUT126), .ZN(new_n1169));
  OAI21_X1  g744(.A(G2105), .B1(new_n1168), .B2(KEYINPUT126), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n1171));
  OAI22_X1  g746(.A1(new_n1169), .A2(new_n1170), .B1(new_n1171), .B2(new_n474), .ZN(new_n1172));
  AOI211_X1 g747(.A(new_n1167), .B(new_n1172), .C1(new_n1171), .C2(new_n474), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(new_n1058), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1174), .B1(new_n1175), .B2(new_n1004), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1080), .A2(G301), .A3(new_n1081), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1166), .B1(new_n1178), .B2(new_n1084), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1180));
  OAI21_X1  g755(.A(G171), .B1(new_n1176), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1082), .A2(G301), .A3(new_n1083), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1181), .A2(new_n1182), .A3(KEYINPUT54), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1162), .A2(new_n1165), .A3(new_n1179), .A4(new_n1183), .ZN(new_n1184));
  OAI211_X1 g759(.A(new_n1103), .B(new_n1107), .C1(new_n1161), .C2(new_n1184), .ZN(new_n1185));
  NOR3_X1   g760(.A1(new_n1036), .A2(new_n1037), .A3(G286), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1073), .A2(new_n1078), .A3(new_n1101), .A4(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT118), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT63), .ZN(new_n1189));
  AND3_X1   g764(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1188), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1078), .A2(KEYINPUT63), .A3(new_n1186), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1101), .B1(new_n1077), .B2(new_n1076), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT119), .ZN(new_n1194));
  OR2_X1    g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1192), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NOR3_X1   g772(.A1(new_n1190), .A2(new_n1191), .A3(new_n1197), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1019), .B1(new_n1185), .B2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g774(.A1(G290), .A2(G1986), .ZN(new_n1200));
  AND2_X1   g775(.A1(new_n1011), .A2(new_n1200), .ZN(new_n1201));
  XOR2_X1   g776(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1202));
  OR2_X1    g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1011), .A2(new_n1017), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1207));
  OAI22_X1  g782(.A1(new_n1207), .A2(new_n1015), .B1(G2067), .B2(new_n777), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1208), .A2(new_n1011), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1206), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g785(.A(new_n1012), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1011), .B1(new_n801), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g787(.A(KEYINPUT46), .ZN(new_n1213));
  AND3_X1   g788(.A1(new_n1011), .A2(new_n1213), .A3(new_n1013), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1213), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1212), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  OR2_X1    g791(.A1(new_n1216), .A2(KEYINPUT47), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1216), .A2(KEYINPUT47), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1210), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1199), .A2(new_n1219), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g795(.A1(G227), .A2(new_n463), .ZN(new_n1222));
  OR3_X1    g796(.A1(G401), .A2(G229), .A3(new_n1222), .ZN(new_n1223));
  NOR2_X1   g797(.A1(new_n971), .A2(new_n980), .ZN(new_n1224));
  NOR3_X1   g798(.A1(new_n911), .A2(new_n1223), .A3(new_n1224), .ZN(G308));
  INV_X1    g799(.A(G308), .ZN(G225));
endmodule


