//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 0 0 1 1 1 1 0 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT0), .A2(G128), .ZN(new_n188));
  XNOR2_X1  g002(.A(G143), .B(G146), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(KEYINPUT64), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT0), .B(G128), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n190), .A2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(KEYINPUT75), .B(G125), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  OAI211_X1 g015(.A(KEYINPUT67), .B(KEYINPUT1), .C1(new_n193), .C2(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G128), .ZN(new_n203));
  AOI21_X1  g017(.A(KEYINPUT67), .B1(new_n192), .B2(KEYINPUT1), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n195), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT1), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n189), .A2(new_n206), .A3(G128), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n201), .B1(new_n200), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT7), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT81), .ZN(new_n212));
  INV_X1    g026(.A(G104), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G107), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT81), .A2(G104), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT3), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT82), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(KEYINPUT3), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n221), .A2(KEYINPUT82), .ZN(new_n222));
  OAI211_X1 g036(.A(G104), .B(new_n215), .C1(new_n220), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n214), .A2(new_n216), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G107), .ZN(new_n225));
  INV_X1    g039(.A(G101), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n218), .A2(new_n223), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT84), .B1(new_n215), .B2(G104), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n217), .A2(new_n228), .ZN(new_n229));
  NOR3_X1   g043(.A1(new_n215), .A2(KEYINPUT84), .A3(G104), .ZN(new_n230));
  OAI21_X1  g044(.A(G101), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G113), .ZN(new_n233));
  XNOR2_X1  g047(.A(G116), .B(G119), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n233), .B1(new_n234), .B2(KEYINPUT5), .ZN(new_n235));
  INV_X1    g049(.A(G119), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G116), .ZN(new_n237));
  OR2_X1    g051(.A1(new_n237), .A2(KEYINPUT5), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n233), .A2(KEYINPUT2), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT2), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G113), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  AOI22_X1  g056(.A1(new_n235), .A2(new_n238), .B1(new_n234), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n232), .A2(new_n243), .ZN(new_n244));
  XOR2_X1   g058(.A(new_n244), .B(KEYINPUT89), .Z(new_n245));
  NAND3_X1  g059(.A1(new_n218), .A2(new_n223), .A3(new_n225), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G101), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT83), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT4), .A4(new_n227), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n247), .A2(KEYINPUT4), .A3(new_n227), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n246), .A2(new_n251), .A3(G101), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT83), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n249), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n242), .B1(new_n234), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G116), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G119), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n237), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT2), .B(G113), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n260), .A3(KEYINPUT68), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n254), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT88), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT88), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n254), .A2(new_n265), .A3(new_n262), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n245), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  XOR2_X1   g081(.A(G110), .B(G122), .Z(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n211), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  XOR2_X1   g084(.A(new_n268), .B(KEYINPUT8), .Z(new_n271));
  INV_X1    g085(.A(new_n244), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n232), .A2(new_n243), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G953), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n209), .A2(G224), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n209), .B1(G224), .B2(new_n275), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT7), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n270), .A2(new_n274), .A3(new_n276), .A4(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n244), .B(KEYINPUT89), .ZN(new_n280));
  INV_X1    g094(.A(new_n262), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n247), .A2(KEYINPUT4), .A3(new_n227), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(KEYINPUT83), .A3(new_n252), .ZN(new_n283));
  AOI211_X1 g097(.A(KEYINPUT88), .B(new_n281), .C1(new_n283), .C2(new_n249), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n265), .B1(new_n254), .B2(new_n262), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n280), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n268), .B(KEYINPUT90), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT6), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n269), .B(new_n280), .C1(new_n284), .C2(new_n285), .ZN(new_n289));
  INV_X1    g103(.A(new_n287), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n289), .B1(new_n267), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n288), .B1(new_n291), .B2(KEYINPUT6), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n275), .A2(G224), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n209), .B(new_n293), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n187), .B(new_n279), .C1(new_n292), .C2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(G210), .B1(G237), .B2(G902), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n294), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT6), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n286), .A2(new_n287), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n300), .B1(new_n301), .B2(new_n289), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n299), .B1(new_n302), .B2(new_n288), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n303), .A2(new_n187), .A3(new_n296), .A4(new_n279), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n298), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(G214), .B1(G237), .B2(G902), .ZN(new_n306));
  XOR2_X1   g120(.A(new_n306), .B(KEYINPUT87), .Z(new_n307));
  XOR2_X1   g121(.A(KEYINPUT9), .B(G234), .Z(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(G221), .B1(new_n309), .B2(G902), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  XOR2_X1   g125(.A(G110), .B(G140), .Z(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(KEYINPUT80), .ZN(new_n313));
  INV_X1    g127(.A(G227), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(G953), .ZN(new_n315));
  XOR2_X1   g129(.A(new_n313), .B(new_n315), .Z(new_n316));
  INV_X1    g130(.A(G131), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT11), .ZN(new_n318));
  INV_X1    g132(.A(G134), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT65), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT65), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G134), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(new_n322), .A3(G137), .ZN(new_n323));
  NOR2_X1   g137(.A1(G134), .A2(G137), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n318), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G137), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n320), .A2(new_n322), .A3(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n328), .A2(KEYINPUT11), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n317), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT65), .B(G134), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(new_n318), .A3(new_n327), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n324), .B1(new_n331), .B2(G137), .ZN(new_n333));
  OAI211_X1 g147(.A(G131), .B(new_n332), .C1(new_n333), .C2(new_n318), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n232), .A2(KEYINPUT10), .A3(new_n208), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n199), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n338), .B1(new_n254), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G128), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n341), .B1(new_n192), .B2(KEYINPUT1), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n207), .B1(new_n342), .B2(new_n189), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n227), .A2(new_n231), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT10), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n336), .B1(new_n340), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n199), .B1(new_n283), .B2(new_n249), .ZN(new_n348));
  INV_X1    g162(.A(new_n346), .ZN(new_n349));
  NOR4_X1   g163(.A1(new_n348), .A2(new_n335), .A3(new_n349), .A4(new_n338), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n316), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT86), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n344), .B1(new_n232), .B2(new_n208), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(KEYINPUT12), .A3(new_n335), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT12), .B1(new_n353), .B2(new_n335), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n352), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n356), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(KEYINPUT86), .A3(new_n354), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n254), .A2(new_n339), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n360), .A2(new_n336), .A3(new_n346), .A4(new_n337), .ZN(new_n361));
  INV_X1    g175(.A(new_n316), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n357), .A2(new_n359), .A3(new_n361), .A4(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n351), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(KEYINPUT85), .A2(G469), .ZN(new_n365));
  NOR2_X1   g179(.A1(KEYINPUT85), .A2(G469), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n364), .A2(new_n187), .A3(new_n365), .A4(new_n367), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n348), .A2(new_n349), .A3(new_n338), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n316), .B1(new_n369), .B2(new_n336), .ZN(new_n370));
  INV_X1    g184(.A(new_n347), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n358), .A2(new_n354), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n361), .A2(new_n372), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n370), .A2(new_n371), .B1(new_n373), .B2(new_n316), .ZN(new_n374));
  OAI21_X1  g188(.A(G469), .B1(new_n374), .B2(G902), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n311), .B1(new_n368), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G478), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(KEYINPUT15), .ZN(new_n378));
  INV_X1    g192(.A(G122), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT94), .B1(new_n379), .B2(G116), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT94), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(new_n257), .A3(G122), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n257), .A2(G122), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n383), .A2(new_n215), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n215), .B1(new_n383), .B2(new_n385), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n341), .A2(G143), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n341), .A2(G143), .ZN(new_n391));
  AOI22_X1  g205(.A1(KEYINPUT13), .A2(new_n390), .B1(new_n391), .B2(KEYINPUT95), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n193), .A2(KEYINPUT95), .A3(KEYINPUT13), .A4(G128), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n393), .B1(new_n390), .B2(KEYINPUT13), .ZN(new_n394));
  OAI21_X1  g208(.A(G134), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n331), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n193), .A2(G128), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT96), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n397), .A2(new_n391), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n398), .B1(new_n397), .B2(new_n391), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n396), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n395), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n389), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n383), .A2(KEYINPUT14), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT97), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(new_n405), .A3(new_n385), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT14), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n380), .A2(new_n382), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n407), .B1(new_n380), .B2(new_n382), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT97), .B1(new_n409), .B2(new_n384), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n406), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n387), .B1(new_n411), .B2(G107), .ZN(new_n412));
  OR3_X1    g226(.A1(new_n399), .A2(new_n396), .A3(new_n400), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n401), .ZN(new_n414));
  AOI211_X1 g228(.A(KEYINPUT98), .B(new_n403), .C1(new_n412), .C2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G217), .ZN(new_n416));
  NOR3_X1   g230(.A1(new_n309), .A2(new_n416), .A3(G953), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n411), .A2(G107), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(new_n386), .A3(new_n414), .ZN(new_n420));
  INV_X1    g234(.A(new_n403), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT98), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n403), .B1(new_n412), .B2(new_n414), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT98), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n418), .B1(new_n417), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n378), .B1(new_n428), .B2(G902), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n425), .B1(new_n420), .B2(new_n421), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n417), .B1(new_n415), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n417), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n426), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n378), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n187), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n429), .A2(KEYINPUT99), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(KEYINPUT99), .B1(new_n429), .B2(new_n436), .ZN(new_n439));
  INV_X1    g253(.A(G475), .ZN(new_n440));
  INV_X1    g254(.A(G237), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(new_n275), .A3(G214), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(new_n193), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G131), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n442), .B(G143), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n317), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  OR2_X1    g261(.A1(new_n447), .A2(KEYINPUT17), .ZN(new_n448));
  INV_X1    g262(.A(new_n200), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n449), .A2(KEYINPUT16), .A3(G140), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n200), .A2(G140), .ZN(new_n451));
  OR2_X1    g265(.A1(G125), .A2(G140), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n450), .B1(new_n453), .B2(KEYINPUT16), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(G146), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n453), .A2(KEYINPUT16), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n191), .B1(new_n456), .B2(new_n450), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n445), .A2(new_n317), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT17), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n448), .A2(new_n455), .A3(new_n457), .A4(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT77), .ZN(new_n461));
  NAND2_X1  g275(.A1(G125), .A2(G140), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n452), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT76), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT76), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n452), .A2(new_n465), .A3(new_n462), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n461), .B1(new_n467), .B2(new_n191), .ZN(new_n468));
  AOI211_X1 g282(.A(KEYINPUT77), .B(G146), .C1(new_n464), .C2(new_n466), .ZN(new_n469));
  OAI22_X1  g283(.A1(new_n468), .A2(new_n469), .B1(new_n191), .B2(new_n453), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT18), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n445), .B1(new_n471), .B2(new_n317), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT91), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n473), .B1(new_n458), .B2(KEYINPUT18), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n444), .A2(KEYINPUT91), .A3(new_n471), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n470), .B(new_n472), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  XOR2_X1   g290(.A(G113), .B(G122), .Z(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(KEYINPUT93), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n478), .B(new_n213), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n460), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n451), .A2(KEYINPUT19), .A3(new_n452), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT92), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT19), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT92), .B1(new_n467), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n484), .B1(new_n486), .B2(new_n482), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n455), .B(new_n447), .C1(new_n487), .C2(G146), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n479), .B1(new_n488), .B2(new_n476), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n440), .B(new_n187), .C1(new_n481), .C2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT20), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n489), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n480), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n494), .A2(KEYINPUT20), .A3(new_n440), .A4(new_n187), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n479), .B1(new_n460), .B2(new_n476), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n187), .B1(new_n481), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(G475), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n492), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n275), .A2(G952), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n500), .B1(G234), .B2(G237), .ZN(new_n501));
  XOR2_X1   g315(.A(KEYINPUT21), .B(G898), .Z(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(G234), .A2(G237), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(G902), .A3(G953), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n501), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  NOR4_X1   g321(.A1(new_n438), .A2(new_n439), .A3(new_n499), .A4(new_n507), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n305), .A2(new_n307), .A3(new_n376), .A4(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT100), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n438), .A2(new_n439), .A3(new_n507), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n492), .A2(new_n495), .A3(new_n498), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n512), .A2(new_n376), .A3(new_n513), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n514), .A2(new_n305), .A3(KEYINPUT100), .A4(new_n307), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT78), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT25), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n455), .A2(new_n457), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n236), .A2(G128), .ZN(new_n519));
  OR2_X1    g333(.A1(new_n519), .A2(KEYINPUT72), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(KEYINPUT72), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n520), .A2(new_n521), .B1(G119), .B2(new_n341), .ZN(new_n522));
  XOR2_X1   g336(.A(KEYINPUT24), .B(G110), .Z(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT73), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n524), .B(new_n525), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n236), .A2(KEYINPUT23), .A3(G128), .ZN(new_n527));
  XNOR2_X1  g341(.A(G119), .B(G128), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n527), .B1(new_n528), .B2(KEYINPUT23), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G110), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(KEYINPUT74), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n518), .A2(new_n526), .A3(new_n531), .ZN(new_n532));
  OAI22_X1  g346(.A1(new_n522), .A2(new_n523), .B1(new_n529), .B2(G110), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n455), .B(new_n533), .C1(new_n469), .C2(new_n468), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n275), .A2(G221), .A3(G234), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(KEYINPUT22), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(G137), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n532), .A2(new_n538), .A3(new_n534), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n516), .B(new_n517), .C1(new_n542), .C2(G902), .ZN(new_n543));
  NAND2_X1  g357(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n516), .A2(new_n517), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n540), .A2(new_n187), .A3(new_n541), .A4(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n416), .B1(G234), .B2(new_n187), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n548), .A2(G902), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(KEYINPUT79), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n540), .A2(new_n551), .A3(new_n541), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(G472), .A2(G902), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n335), .A2(new_n339), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n319), .A2(G137), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n328), .A2(KEYINPUT66), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT66), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n331), .A2(new_n558), .A3(new_n327), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n557), .A2(G131), .A3(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n330), .A2(new_n208), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n555), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n262), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT28), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n330), .A2(new_n208), .A3(new_n560), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n199), .B1(new_n330), .B2(new_n334), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n256), .A2(new_n261), .A3(KEYINPUT69), .ZN(new_n568));
  AOI21_X1  g382(.A(KEYINPUT69), .B1(new_n256), .B2(new_n261), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n564), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  NOR4_X1   g386(.A1(new_n565), .A2(new_n566), .A3(new_n570), .A4(KEYINPUT28), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n563), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(G101), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n441), .A2(new_n275), .A3(G210), .ZN(new_n577));
  XOR2_X1   g391(.A(new_n576), .B(new_n577), .Z(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT30), .B1(new_n565), .B2(new_n566), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT30), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n555), .A2(new_n582), .A3(new_n561), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n262), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT31), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n555), .A2(new_n571), .A3(new_n561), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n585), .A2(new_n586), .A3(new_n587), .A4(new_n578), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n580), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n281), .B1(new_n581), .B2(new_n583), .ZN(new_n590));
  INV_X1    g404(.A(new_n587), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n586), .B1(new_n592), .B2(new_n578), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n554), .B1(new_n589), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT32), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g410(.A(KEYINPUT32), .B(new_n554), .C1(new_n589), .C2(new_n593), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(KEYINPUT70), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT70), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n594), .A2(new_n599), .A3(new_n595), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT29), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n587), .A2(KEYINPUT28), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n567), .A2(new_n564), .A3(new_n571), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n579), .B1(new_n605), .B2(new_n563), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n590), .A2(new_n591), .A3(new_n578), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n602), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT71), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT71), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n610), .B(new_n602), .C1(new_n606), .C2(new_n607), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n562), .A2(new_n570), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n605), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(new_n602), .ZN(new_n614));
  AOI21_X1  g428(.A(G902), .B1(new_n614), .B2(new_n578), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n609), .A2(new_n611), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(G472), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n553), .B1(new_n601), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n511), .A2(new_n515), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G101), .ZN(G3));
  AOI21_X1  g434(.A(G478), .B1(new_n434), .B2(new_n187), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  OR3_X1    g436(.A1(new_n424), .A2(KEYINPUT101), .A3(new_n417), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n417), .B1(new_n424), .B2(KEYINPUT101), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(KEYINPUT33), .A3(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT102), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT33), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT102), .B1(new_n434), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n627), .B1(new_n629), .B2(new_n625), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n187), .A2(G478), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n622), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT103), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(new_n633), .A3(new_n499), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n633), .B1(new_n632), .B2(new_n499), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n507), .ZN(new_n638));
  INV_X1    g452(.A(new_n306), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n639), .B1(new_n298), .B2(new_n304), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n637), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n553), .A2(new_n311), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n368), .A2(new_n375), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n187), .B1(new_n589), .B2(new_n593), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(G472), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n646), .A2(new_n594), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n643), .A2(new_n644), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n642), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT104), .B(KEYINPUT34), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G104), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n649), .B(new_n651), .ZN(G6));
  INV_X1    g466(.A(KEYINPUT99), .ZN(new_n653));
  INV_X1    g467(.A(new_n436), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n435), .B1(new_n434), .B2(new_n187), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n499), .B1(new_n656), .B2(new_n437), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n507), .B(KEYINPUT105), .Z(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n648), .A2(new_n640), .A3(new_n657), .A4(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT35), .B(G107), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  NOR2_X1   g476(.A1(new_n539), .A2(KEYINPUT36), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n535), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n551), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n549), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n511), .A2(new_n515), .A3(new_n647), .A4(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n667), .B(KEYINPUT37), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G110), .ZN(G12));
  NAND2_X1  g483(.A1(new_n644), .A2(new_n310), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n617), .B2(new_n601), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n501), .B(KEYINPUT107), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT106), .B(G900), .Z(new_n674));
  OAI21_X1  g488(.A(new_n673), .B1(new_n505), .B2(new_n674), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n657), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n671), .A2(new_n640), .A3(new_n666), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  NOR2_X1   g492(.A1(new_n592), .A2(new_n579), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n612), .A2(new_n587), .A3(new_n579), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n187), .ZN(new_n681));
  OAI21_X1  g495(.A(G472), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n601), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT38), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n298), .A2(new_n686), .A3(new_n304), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n686), .B1(new_n298), .B2(new_n304), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n685), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n689), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(KEYINPUT38), .A3(new_n687), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n684), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  XOR2_X1   g507(.A(new_n675), .B(KEYINPUT39), .Z(new_n694));
  NOR2_X1   g508(.A1(new_n670), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT40), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n666), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n695), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT40), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n306), .B(new_n499), .C1(new_n438), .C2(new_n439), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n693), .A2(new_n697), .A3(new_n699), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G143), .ZN(G45));
  OAI211_X1 g517(.A(new_n626), .B(new_n625), .C1(new_n428), .C2(KEYINPUT33), .ZN(new_n704));
  INV_X1    g518(.A(new_n627), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n631), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n499), .B(new_n675), .C1(new_n706), .C2(new_n621), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n671), .A2(new_n640), .A3(new_n666), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  NAND2_X1  g524(.A1(new_n364), .A2(new_n187), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(G469), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n368), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n311), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n618), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n642), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  NAND3_X1  g533(.A1(new_n640), .A2(new_n657), .A3(new_n659), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(new_n715), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n257), .ZN(G18));
  NAND3_X1  g536(.A1(new_n640), .A2(new_n666), .A3(new_n714), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n601), .A2(new_n617), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n508), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(KEYINPUT109), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  AOI21_X1  g542(.A(new_n700), .B1(new_n298), .B2(new_n304), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n578), .B1(new_n605), .B2(new_n612), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n730), .B1(new_n593), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n613), .A2(new_n579), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n590), .A2(new_n591), .A3(new_n579), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n733), .B(KEYINPUT110), .C1(new_n586), .C2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n732), .A2(new_n735), .A3(new_n588), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n554), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n646), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n738), .A2(new_n553), .A3(new_n658), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n729), .A2(new_n714), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G122), .ZN(G24));
  NOR2_X1   g555(.A1(new_n707), .A2(new_n738), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n640), .A2(new_n666), .A3(new_n742), .A4(new_n714), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G125), .ZN(G27));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n617), .A2(new_n596), .A3(new_n597), .ZN(new_n746));
  INV_X1    g560(.A(new_n553), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n632), .A2(KEYINPUT42), .A3(new_n499), .A4(new_n675), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n298), .A2(new_n304), .A3(new_n306), .A4(new_n376), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n745), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n708), .A2(KEYINPUT42), .A3(new_n747), .A4(new_n746), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n754), .A2(KEYINPUT111), .A3(new_n751), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n724), .A2(new_n747), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n756), .A2(new_n707), .A3(new_n751), .ZN(new_n757));
  OAI22_X1  g571(.A1(new_n753), .A2(new_n755), .B1(new_n757), .B2(KEYINPUT42), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G131), .ZN(G33));
  NOR2_X1   g573(.A1(new_n756), .A2(new_n751), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n676), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G134), .ZN(G36));
  NAND2_X1  g576(.A1(new_n632), .A2(new_n513), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT43), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n632), .A2(KEYINPUT43), .A3(new_n513), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n647), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT44), .B1(new_n767), .B2(new_n666), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n768), .A2(new_n305), .A3(new_n639), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n767), .A2(KEYINPUT44), .A3(new_n666), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n770), .A2(KEYINPUT114), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(KEYINPUT114), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n769), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT115), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n374), .A2(KEYINPUT45), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n374), .A2(KEYINPUT45), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(G469), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(G469), .A2(G902), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT46), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n777), .A2(KEYINPUT46), .A3(new_n778), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(new_n368), .A3(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n694), .ZN(new_n784));
  XNOR2_X1  g598(.A(KEYINPUT112), .B(KEYINPUT113), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n783), .A2(new_n310), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n785), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n783), .A2(new_n310), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n787), .B1(new_n788), .B2(new_n694), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT115), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n769), .A2(new_n771), .A3(new_n790), .A4(new_n772), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n774), .A2(new_n786), .A3(new_n789), .A4(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G137), .ZN(G39));
  XNOR2_X1  g607(.A(new_n788), .B(KEYINPUT47), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n794), .A2(new_n724), .A3(new_n707), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n305), .A2(new_n639), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n553), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G140), .ZN(G42));
  OR2_X1    g612(.A1(new_n713), .A2(KEYINPUT49), .ZN(new_n799));
  AND4_X1   g613(.A1(new_n684), .A2(new_n690), .A3(new_n692), .A4(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n763), .B1(KEYINPUT49), .B2(new_n713), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n800), .A2(new_n307), .A3(new_n643), .A4(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n740), .B1(new_n641), .B2(new_n715), .ZN(new_n803));
  OAI22_X1  g617(.A1(new_n720), .A2(new_n715), .B1(new_n723), .B2(new_n725), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n305), .A2(new_n307), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n632), .A2(new_n499), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n654), .A2(new_n655), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n807), .B1(new_n499), .B2(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n806), .A2(new_n648), .A3(new_n659), .A4(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n667), .A2(new_n619), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n805), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n644), .A2(new_n310), .A3(new_n675), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n305), .A2(new_n701), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n666), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n683), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n813), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n666), .B1(new_n601), .B2(new_n682), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n729), .A2(new_n819), .A3(KEYINPUT116), .A4(new_n814), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n677), .A2(new_n709), .A3(new_n743), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(KEYINPUT52), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n818), .A2(new_n820), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n677), .A2(new_n709), .A3(new_n743), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  AND4_X1   g642(.A1(new_n724), .A2(new_n513), .A3(new_n808), .A4(new_n675), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n666), .B(new_n752), .C1(new_n829), .C2(new_n742), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n758), .A2(new_n761), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n812), .A2(new_n828), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT54), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n713), .A2(new_n306), .A3(new_n311), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n690), .A2(new_n692), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT118), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n765), .A2(new_n766), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n672), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n840), .A2(new_n553), .A3(new_n738), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n690), .A2(new_n692), .A3(new_n842), .A4(new_n836), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n838), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT50), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n796), .A2(new_n714), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n684), .A2(new_n501), .ZN(new_n848));
  NOR4_X1   g662(.A1(new_n847), .A2(new_n848), .A3(new_n553), .A4(new_n632), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n847), .A2(new_n840), .A3(new_n816), .ZN(new_n850));
  INV_X1    g664(.A(new_n738), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n849), .A2(new_n513), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n794), .B1(new_n310), .B2(new_n713), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(new_n796), .A3(new_n841), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n846), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT51), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n500), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n667), .A2(new_n619), .A3(new_n810), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n803), .A2(new_n804), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n750), .A2(new_n752), .A3(new_n745), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT111), .B1(new_n754), .B2(new_n751), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n752), .A2(new_n618), .A3(new_n708), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT42), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n862), .A2(new_n865), .B1(new_n676), .B2(new_n760), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n858), .A2(new_n859), .A3(new_n866), .A4(new_n830), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT52), .B1(new_n821), .B2(new_n822), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n825), .A2(new_n826), .A3(new_n824), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n833), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n859), .A2(KEYINPUT117), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT117), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n874), .B1(new_n803), .B2(new_n804), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n811), .B1(new_n823), .B2(new_n827), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n758), .A2(KEYINPUT53), .A3(new_n761), .A4(new_n830), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n871), .A2(new_n872), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n846), .A2(KEYINPUT51), .A3(new_n852), .A4(new_n854), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n835), .A2(new_n857), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n637), .ZN(new_n885));
  NOR4_X1   g699(.A1(new_n847), .A2(new_n885), .A3(new_n848), .A4(new_n553), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n841), .A2(new_n640), .A3(new_n714), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n847), .A2(new_n840), .A3(new_n748), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT48), .ZN(new_n889));
  NOR4_X1   g703(.A1(new_n884), .A2(new_n886), .A3(new_n887), .A4(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(G952), .A2(G953), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n802), .B1(new_n890), .B2(new_n891), .ZN(G75));
  AOI21_X1  g706(.A(new_n878), .B1(new_n875), .B2(new_n873), .ZN(new_n893));
  AOI22_X1  g707(.A1(new_n833), .A2(new_n832), .B1(new_n893), .B2(new_n877), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n894), .A2(new_n187), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(G210), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT56), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n292), .B(new_n299), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT55), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n896), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n899), .B1(new_n896), .B2(new_n897), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n275), .A2(G952), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT119), .Z(new_n903));
  NOR3_X1   g717(.A1(new_n900), .A2(new_n901), .A3(new_n903), .ZN(G51));
  OR2_X1    g718(.A1(new_n778), .A2(KEYINPUT57), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n778), .A2(KEYINPUT57), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n872), .B1(new_n871), .B2(new_n880), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n905), .B(new_n906), .C1(new_n881), .C2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT120), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n908), .A2(new_n909), .A3(new_n364), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n909), .B1(new_n908), .B2(new_n364), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OR3_X1    g726(.A1(new_n894), .A2(new_n187), .A3(new_n777), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n902), .B1(new_n912), .B2(new_n913), .ZN(G54));
  NAND3_X1  g728(.A1(new_n895), .A2(KEYINPUT58), .A3(G475), .ZN(new_n915));
  INV_X1    g729(.A(new_n494), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n915), .A2(new_n916), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n917), .A2(new_n918), .A3(new_n902), .ZN(G60));
  INV_X1    g733(.A(new_n903), .ZN(new_n920));
  NAND2_X1  g734(.A1(G478), .A2(G902), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT59), .Z(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n835), .B2(new_n882), .ZN(new_n923));
  INV_X1    g737(.A(new_n630), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n924), .B1(new_n881), .B2(new_n907), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n926), .A2(new_n922), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n925), .A2(new_n927), .ZN(G63));
  NAND2_X1  g742(.A1(G217), .A2(G902), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT60), .ZN(new_n930));
  OAI21_X1  g744(.A(KEYINPUT121), .B1(new_n894), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n871), .A2(new_n880), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT121), .ZN(new_n933));
  INV_X1    g747(.A(new_n930), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n931), .A2(new_n542), .A3(new_n935), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n936), .A2(new_n920), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n931), .A2(new_n935), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n664), .A2(KEYINPUT122), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n664), .A2(KEYINPUT122), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n938), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT123), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n937), .B(new_n942), .C1(new_n943), .C2(KEYINPUT61), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n936), .A2(new_n943), .A3(new_n920), .ZN(new_n946));
  INV_X1    g760(.A(new_n941), .ZN(new_n947));
  AOI211_X1 g761(.A(new_n939), .B(new_n947), .C1(new_n931), .C2(new_n935), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n936), .A2(new_n920), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n945), .B(new_n946), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n944), .A2(new_n950), .ZN(G66));
  INV_X1    g765(.A(G224), .ZN(new_n952));
  OAI21_X1  g766(.A(G953), .B1(new_n503), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n812), .B2(G953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n292), .B1(G898), .B2(new_n275), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(G69));
  XOR2_X1   g770(.A(new_n584), .B(KEYINPUT124), .Z(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(new_n487), .Z(new_n958));
  AOI21_X1  g772(.A(new_n698), .B1(new_n809), .B2(KEYINPUT125), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n809), .A2(KEYINPUT125), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n959), .A2(new_n618), .A3(new_n796), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n792), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(KEYINPUT126), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT126), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n792), .A2(new_n964), .A3(new_n961), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n702), .A2(new_n822), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT62), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n969), .A2(new_n797), .ZN(new_n970));
  AOI211_X1 g784(.A(G953), .B(new_n958), .C1(new_n966), .C2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n958), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(new_n314), .B2(G953), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(G900), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n975), .B1(new_n972), .B2(new_n314), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n275), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n748), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n789), .A2(new_n729), .A3(new_n978), .A4(new_n786), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n979), .A2(new_n866), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n792), .A2(new_n797), .A3(new_n822), .A4(new_n980), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n981), .A2(new_n974), .ZN(new_n982));
  OR3_X1    g796(.A1(new_n971), .A2(new_n977), .A3(new_n982), .ZN(G72));
  NAND2_X1  g797(.A1(G472), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT63), .Z(new_n985));
  INV_X1    g799(.A(new_n812), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n985), .B1(new_n981), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n607), .ZN(new_n988));
  INV_X1    g802(.A(new_n607), .ZN(new_n989));
  INV_X1    g803(.A(new_n679), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n834), .A2(new_n989), .A3(new_n990), .A4(new_n985), .ZN(new_n991));
  INV_X1    g805(.A(new_n902), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n988), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT127), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n966), .A2(new_n970), .A3(new_n812), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n995), .A2(new_n985), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n993), .B(new_n994), .C1(new_n996), .C2(new_n990), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n990), .B1(new_n995), .B2(new_n985), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n988), .A2(new_n991), .A3(new_n992), .ZN(new_n999));
  OAI21_X1  g813(.A(KEYINPUT127), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n997), .A2(new_n1000), .ZN(G57));
endmodule


