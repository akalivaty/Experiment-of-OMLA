//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n559, new_n560, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1184,
    new_n1185, new_n1186;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT64), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G236), .A2(G238), .A3(G237), .A4(G235), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT66), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND3_X1  g034(.A1(new_n455), .A2(KEYINPUT67), .A3(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g037(.A(KEYINPUT67), .B1(new_n455), .B2(G2106), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n464), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n467));
  AND3_X1   g042(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(KEYINPUT3), .B1(new_n467), .B2(G2104), .ZN(new_n469));
  OAI211_X1 g044(.A(G137), .B(new_n466), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n475));
  AND2_X1   g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n475), .B1(new_n478), .B2(new_n466), .ZN(new_n479));
  INV_X1    g054(.A(G125), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(new_n471), .ZN(new_n482));
  NAND2_X1  g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI211_X1 g059(.A(KEYINPUT69), .B(G2105), .C1(new_n484), .C2(new_n476), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n474), .B1(new_n479), .B2(new_n485), .ZN(G160));
  OAI21_X1  g061(.A(new_n481), .B1(new_n471), .B2(KEYINPUT70), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n466), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  NOR2_X1   g065(.A1(G100), .A2(G2105), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT72), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(new_n466), .B2(G112), .ZN(new_n493));
  AOI21_X1  g068(.A(G2105), .B1(new_n487), .B2(new_n488), .ZN(new_n494));
  AND3_X1   g069(.A1(new_n494), .A2(KEYINPUT71), .A3(G136), .ZN(new_n495));
  AOI21_X1  g070(.A(KEYINPUT71), .B1(new_n494), .B2(G136), .ZN(new_n496));
  OAI221_X1 g071(.A(new_n490), .B1(new_n492), .B2(new_n493), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  XOR2_X1   g072(.A(new_n497), .B(KEYINPUT73), .Z(G162));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n466), .A2(G138), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n477), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n500), .B1(new_n487), .B2(new_n488), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(new_n499), .ZN(new_n504));
  OAI21_X1  g079(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(G114), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(G2105), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n507), .B1(new_n489), .B2(G126), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  NAND2_X1  g085(.A1(KEYINPUT74), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(KEYINPUT74), .A2(KEYINPUT5), .A3(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G50), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n515), .A2(G62), .ZN(new_n523));
  NAND2_X1  g098(.A1(G75), .A2(G543), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT75), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n522), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n521), .A2(new_n526), .ZN(G166));
  NAND3_X1  g102(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n516), .A2(G51), .A3(G543), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n528), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AND3_X1   g107(.A1(new_n515), .A2(G89), .A3(new_n516), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(G168));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n517), .A2(new_n535), .B1(new_n519), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n515), .A2(G64), .ZN(new_n538));
  NAND2_X1  g113(.A1(G77), .A2(G543), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n522), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n537), .A2(new_n540), .ZN(G171));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(new_n514), .ZN(new_n543));
  AOI21_X1  g118(.A(KEYINPUT5), .B1(KEYINPUT74), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n542), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G651), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(KEYINPUT76), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT76), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n547), .A2(new_n550), .A3(G651), .ZN(new_n551));
  AND2_X1   g126(.A1(new_n515), .A2(new_n516), .ZN(new_n552));
  INV_X1    g127(.A(new_n519), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n552), .A2(G81), .B1(new_n553), .B2(G43), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n549), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n545), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n564), .A2(G651), .B1(new_n552), .B2(G91), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n516), .A2(G53), .A3(G543), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT9), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(G299));
  OR2_X1    g143(.A1(new_n537), .A2(new_n540), .ZN(G301));
  AND2_X1   g144(.A1(new_n530), .A2(new_n531), .ZN(new_n570));
  INV_X1    g145(.A(new_n533), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .A4(new_n528), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT77), .B1(new_n532), .B2(new_n533), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G286));
  INV_X1    g151(.A(G166), .ZN(G303));
  AOI22_X1  g152(.A1(new_n552), .A2(G87), .B1(new_n553), .B2(G49), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(G288));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n581), .B1(new_n513), .B2(new_n514), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n515), .A2(G86), .A3(new_n516), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n516), .A2(G48), .A3(G543), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(G305));
  AOI22_X1  g163(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  OR3_X1    g164(.A1(new_n589), .A2(KEYINPUT78), .A3(new_n522), .ZN(new_n590));
  OAI21_X1  g165(.A(KEYINPUT78), .B1(new_n589), .B2(new_n522), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n552), .A2(G85), .B1(new_n553), .B2(G47), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  INV_X1    g170(.A(G92), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n517), .B2(new_n596), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n515), .A2(KEYINPUT10), .A3(new_n516), .A4(G92), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n545), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(new_n553), .B2(G54), .ZN(new_n603));
  AND2_X1   g178(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n594), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n594), .B1(new_n604), .B2(G868), .ZN(G321));
  AND3_X1   g181(.A1(G286), .A2(KEYINPUT79), .A3(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(G286), .A2(G868), .ZN(new_n608));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  AOI21_X1  g184(.A(KEYINPUT79), .B1(G299), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n607), .B1(new_n608), .B2(new_n610), .ZN(G297));
  AOI21_X1  g186(.A(new_n607), .B1(new_n608), .B2(new_n610), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n604), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n604), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n494), .A2(G135), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT82), .Z(new_n620));
  NAND2_X1  g195(.A1(new_n489), .A2(G123), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT83), .ZN(new_n622));
  OR2_X1    g197(.A1(G99), .A2(G2105), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n623), .B(G2104), .C1(G111), .C2(new_n466), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n620), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n625), .A2(KEYINPUT84), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(KEYINPUT84), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(G2096), .Z(new_n629));
  NAND2_X1  g204(.A1(new_n477), .A2(new_n472), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  INV_X1    g207(.A(G2100), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT80), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n632), .A2(new_n633), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT81), .Z(new_n637));
  NAND3_X1  g212(.A1(new_n629), .A2(new_n635), .A3(new_n637), .ZN(G156));
  INV_X1    g213(.A(KEYINPUT14), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(new_n642), .B2(new_n641), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n644), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  AND3_X1   g227(.A1(new_n651), .A2(new_n652), .A3(G14), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT85), .ZN(G401));
  XNOR2_X1  g229(.A(G2084), .B(G2090), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT86), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(KEYINPUT17), .ZN(new_n661));
  OAI211_X1 g236(.A(new_n656), .B(new_n660), .C1(new_n661), .C2(new_n658), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT87), .ZN(new_n663));
  INV_X1    g238(.A(new_n656), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n664), .A2(new_n661), .A3(new_n658), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT88), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n656), .A2(new_n658), .A3(new_n659), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT18), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n663), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2096), .B(G2100), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  OR2_X1    g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G1971), .B(G1976), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n672), .A2(new_n673), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n674), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n676), .A2(KEYINPUT90), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n672), .A2(new_n673), .A3(KEYINPUT89), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT89), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n676), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT20), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G1981), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT91), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n687), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT92), .B(G1986), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n692), .A2(new_n693), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(G229));
  INV_X1    g271(.A(KEYINPUT102), .ZN(new_n697));
  INV_X1    g272(.A(G25), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n698), .A2(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n494), .A2(G131), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n489), .A2(G119), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n466), .A2(G107), .ZN(new_n702));
  OAI21_X1  g277(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n700), .B(new_n701), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT93), .Z(new_n705));
  AOI21_X1  g280(.A(new_n699), .B1(new_n705), .B2(G29), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT94), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI211_X1 g283(.A(KEYINPUT94), .B(new_n699), .C1(new_n705), .C2(G29), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT35), .B(G1991), .Z(new_n710));
  OR3_X1    g285(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(G16), .A2(G24), .ZN(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(G290), .B2(new_n713), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(KEYINPUT95), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(KEYINPUT95), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G1986), .ZN(new_n718));
  INV_X1    g293(.A(G1986), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n715), .A2(new_n719), .A3(new_n716), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n710), .B1(new_n708), .B2(new_n709), .ZN(new_n722));
  AND3_X1   g297(.A1(new_n711), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT34), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n713), .A2(G23), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G288), .B2(G16), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT33), .B(G1976), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(G166), .A2(new_n713), .ZN(new_n729));
  INV_X1    g304(.A(G1971), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n713), .A2(G22), .ZN(new_n731));
  OR3_X1    g306(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n730), .B1(new_n729), .B2(new_n731), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OR2_X1    g309(.A1(G305), .A2(new_n713), .ZN(new_n735));
  OR2_X1    g310(.A1(G6), .A2(G16), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT32), .B(G1981), .ZN(new_n737));
  AND3_X1   g312(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n737), .B1(new_n735), .B2(new_n736), .ZN(new_n739));
  OAI21_X1  g314(.A(KEYINPUT96), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n735), .A2(new_n736), .ZN(new_n741));
  INV_X1    g316(.A(new_n737), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT96), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n728), .A2(new_n734), .A3(new_n740), .A4(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT97), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n724), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n747), .A2(new_n748), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n747), .A2(new_n748), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n752), .A2(KEYINPUT34), .A3(new_n753), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n723), .A2(new_n751), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(KEYINPUT36), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT36), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n723), .A2(new_n751), .A3(new_n754), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(G29), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(G26), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT28), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n494), .A2(G140), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT98), .ZN(new_n764));
  OAI21_X1  g339(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n765));
  INV_X1    g340(.A(G116), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n765), .B1(new_n766), .B2(G2105), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n489), .B2(G128), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n762), .B1(new_n769), .B2(G29), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2067), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n626), .A2(G29), .A3(new_n627), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n760), .A2(G33), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT25), .Z(new_n775));
  NAND2_X1  g350(.A1(new_n494), .A2(G139), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n775), .B(new_n776), .C1(new_n466), .C2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n773), .B1(new_n778), .B2(G29), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n779), .A2(new_n442), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n713), .A2(G21), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G168), .B2(new_n713), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n782), .A2(G1966), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n779), .A2(new_n442), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n780), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n713), .A2(G20), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT23), .Z(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G299), .B2(G16), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1956), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n771), .A2(new_n772), .A3(new_n785), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n713), .A2(G19), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n556), .B2(new_n713), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G1341), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n713), .A2(G4), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n604), .B2(new_n713), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(G1348), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT24), .ZN(new_n797));
  INV_X1    g372(.A(G34), .ZN(new_n798));
  AOI21_X1  g373(.A(G29), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n797), .B2(new_n798), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G160), .B2(new_n760), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(G2084), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n795), .A2(G1348), .ZN(new_n803));
  NOR2_X1   g378(.A1(G5), .A2(G16), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT99), .Z(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G171), .B2(G16), .ZN(new_n806));
  INV_X1    g381(.A(G1961), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n796), .A2(new_n802), .A3(new_n803), .A4(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(G27), .A2(G29), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G164), .B2(G29), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(new_n443), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n760), .A2(G32), .ZN(new_n813));
  NAND3_X1  g388(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT26), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n814), .A2(new_n815), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n816), .A2(new_n817), .B1(G105), .B2(new_n472), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n494), .A2(G141), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n489), .A2(G129), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n813), .B1(new_n821), .B2(G29), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT27), .B(G1996), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G1966), .B2(new_n782), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n801), .A2(G2084), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT30), .ZN(new_n827));
  AND2_X1   g402(.A1(new_n827), .A2(G28), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n760), .B1(new_n827), .B2(G28), .ZN(new_n829));
  AND2_X1   g404(.A1(KEYINPUT31), .A2(G11), .ZN(new_n830));
  NOR2_X1   g405(.A1(KEYINPUT31), .A2(G11), .ZN(new_n831));
  OAI22_X1  g406(.A1(new_n828), .A2(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(new_n822), .B2(new_n823), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n812), .A2(new_n825), .A3(new_n826), .A4(new_n833), .ZN(new_n834));
  NOR4_X1   g409(.A1(new_n790), .A2(new_n793), .A3(new_n809), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n760), .A2(G35), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT100), .Z(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(G162), .B2(new_n760), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT29), .ZN(new_n839));
  INV_X1    g414(.A(G2090), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT29), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n841), .B(new_n837), .C1(G162), .C2(new_n760), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n839), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT101), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n839), .A2(new_n842), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n844), .B1(new_n845), .B2(G2090), .ZN(new_n846));
  AOI211_X1 g421(.A(KEYINPUT101), .B(new_n840), .C1(new_n839), .C2(new_n842), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n835), .B(new_n843), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n697), .B1(new_n759), .B2(new_n849), .ZN(new_n850));
  AOI211_X1 g425(.A(KEYINPUT102), .B(new_n848), .C1(new_n756), .C2(new_n758), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(G311));
  AOI21_X1  g427(.A(KEYINPUT103), .B1(new_n759), .B2(new_n849), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT103), .ZN(new_n854));
  AOI211_X1 g429(.A(new_n854), .B(new_n848), .C1(new_n756), .C2(new_n758), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n853), .A2(new_n855), .ZN(G150));
  NAND2_X1  g431(.A1(new_n604), .A2(G559), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT38), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n515), .A2(G93), .A3(new_n516), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n516), .A2(G55), .A3(G543), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT104), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT104), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n859), .A2(new_n863), .A3(new_n860), .ZN(new_n864));
  NAND2_X1  g439(.A1(G80), .A2(G543), .ZN(new_n865));
  INV_X1    g440(.A(G67), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n865), .B1(new_n545), .B2(new_n866), .ZN(new_n867));
  AOI22_X1  g442(.A1(new_n862), .A2(new_n864), .B1(G651), .B2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n555), .B(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n858), .B(new_n869), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n870), .A2(KEYINPUT39), .ZN(new_n871));
  INV_X1    g446(.A(G860), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(KEYINPUT39), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n868), .A2(new_n872), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT37), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(G145));
  NAND2_X1  g452(.A1(new_n489), .A2(G130), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT105), .ZN(new_n879));
  NOR3_X1   g454(.A1(new_n879), .A2(new_n466), .A3(G118), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n879), .B1(new_n466), .B2(G118), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n881), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n878), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n883), .B1(G142), .B2(new_n494), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n884), .B(new_n631), .Z(new_n885));
  XNOR2_X1  g460(.A(new_n778), .B(new_n821), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n769), .B(new_n509), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n704), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n887), .B(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(G162), .B(G160), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(new_n628), .ZN(new_n892));
  AOI21_X1  g467(.A(G37), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n893), .B1(new_n892), .B2(new_n890), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g470(.A(G290), .B(G305), .ZN(new_n896));
  XNOR2_X1  g471(.A(G288), .B(G166), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n896), .B(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(KEYINPUT109), .B1(new_n899), .B2(KEYINPUT108), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n898), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT42), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n869), .B(new_n615), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT41), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n565), .A2(new_n567), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n599), .A2(new_n603), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n908), .A2(KEYINPUT106), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n604), .A2(G299), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT106), .B1(new_n908), .B2(new_n909), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n907), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT107), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n908), .A2(new_n909), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n911), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n915), .B1(new_n917), .B2(new_n907), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n916), .A2(new_n911), .A3(KEYINPUT107), .A4(KEYINPUT41), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n914), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n906), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n917), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n921), .B1(new_n906), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n900), .A2(new_n924), .A3(new_n903), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n905), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n923), .B1(new_n905), .B2(new_n925), .ZN(new_n927));
  OAI21_X1  g502(.A(G868), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(G868), .B2(new_n868), .ZN(G295));
  OAI21_X1  g504(.A(new_n928), .B1(G868), .B2(new_n868), .ZN(G331));
  INV_X1    g505(.A(KEYINPUT111), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n573), .A2(new_n574), .A3(G171), .A4(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n575), .A2(G301), .ZN(new_n933));
  INV_X1    g508(.A(G168), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT111), .B1(new_n934), .B2(G171), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n932), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n869), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n931), .B1(G301), .B2(G168), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(G301), .B2(new_n575), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n556), .A2(new_n868), .ZN(new_n940));
  INV_X1    g515(.A(new_n868), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n941), .A2(new_n555), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n939), .B(new_n932), .C1(new_n940), .C2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n937), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n920), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n917), .B1(new_n937), .B2(new_n943), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n899), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G37), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n944), .A2(new_n922), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n949), .B(new_n898), .C1(new_n920), .C2(new_n944), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n947), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT112), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n951), .A2(new_n952), .A3(KEYINPUT43), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n952), .B1(new_n951), .B2(KEYINPUT43), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n922), .B1(new_n944), .B2(new_n907), .ZN(new_n955));
  OR2_X1    g530(.A1(new_n912), .A2(new_n913), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n956), .A2(new_n937), .A3(new_n943), .A4(KEYINPUT41), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n955), .A2(new_n898), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n947), .A2(new_n958), .A3(new_n948), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n953), .A2(new_n954), .A3(new_n960), .ZN(new_n961));
  XOR2_X1   g536(.A(KEYINPUT110), .B(KEYINPUT44), .Z(new_n962));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n963), .B1(new_n959), .B2(KEYINPUT43), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT113), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n947), .A2(new_n950), .A3(new_n966), .A4(new_n948), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n965), .B1(new_n964), .B2(new_n967), .ZN(new_n969));
  OAI22_X1  g544(.A1(new_n961), .A2(new_n962), .B1(new_n968), .B2(new_n969), .ZN(G397));
  INV_X1    g545(.A(G1384), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n499), .A2(new_n466), .A3(G138), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n972), .B1(new_n482), .B2(new_n483), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n501), .B1(new_n468), .B2(new_n469), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n973), .B1(new_n974), .B2(KEYINPUT4), .ZN(new_n975));
  OAI211_X1 g550(.A(G126), .B(G2105), .C1(new_n468), .C2(new_n469), .ZN(new_n976));
  INV_X1    g551(.A(new_n507), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n971), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n479), .A2(new_n485), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n470), .A2(new_n473), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n982), .A2(G40), .A3(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n769), .A2(G2067), .ZN(new_n986));
  INV_X1    g561(.A(G2067), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n764), .A2(new_n987), .A3(new_n768), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n821), .A2(G1996), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n985), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n985), .A2(G1996), .A3(new_n821), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n992), .A2(new_n993), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n991), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  XOR2_X1   g571(.A(new_n996), .B(KEYINPUT115), .Z(new_n997));
  INV_X1    g572(.A(new_n985), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n704), .B(new_n710), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(G290), .B(G1986), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1000), .B1(new_n985), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT127), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n1004));
  INV_X1    g579(.A(G40), .ZN(new_n1005));
  AOI211_X1 g580(.A(new_n1005), .B(new_n474), .C1(new_n479), .C2(new_n485), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n980), .A2(G1384), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(new_n975), .B2(new_n978), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT116), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT116), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n509), .A2(new_n1010), .A3(new_n1007), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1006), .A2(new_n981), .A3(new_n1009), .A4(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1004), .B1(new_n1012), .B2(G2078), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT124), .ZN(new_n1014));
  XNOR2_X1  g589(.A(KEYINPUT118), .B(KEYINPUT50), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n971), .B(new_n1015), .C1(new_n975), .C2(new_n978), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1016), .A2(G160), .A3(G40), .ZN(new_n1017));
  AOI21_X1  g592(.A(G1384), .B1(new_n504), .B2(new_n508), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1014), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n979), .A2(KEYINPUT50), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1006), .A2(new_n1022), .A3(KEYINPUT124), .A4(new_n1016), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1021), .A2(new_n807), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1013), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n981), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1026));
  OAI21_X1  g601(.A(G2105), .B1(new_n484), .B2(new_n476), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n983), .A2(KEYINPUT125), .A3(G40), .A4(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT125), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(G40), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1029), .B1(new_n1030), .B2(new_n474), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1004), .A2(G2078), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1028), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT126), .B1(new_n1026), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1033), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT126), .ZN(new_n1036));
  AOI22_X1  g611(.A1(KEYINPUT116), .A2(new_n1008), .B1(new_n979), .B2(new_n980), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1011), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(G171), .B1(new_n1025), .B2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1006), .A2(new_n981), .A3(new_n1008), .A4(new_n1032), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1013), .A2(new_n1024), .A3(G301), .A4(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1040), .A2(KEYINPUT54), .A3(new_n1042), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1017), .A2(G2090), .A3(new_n1020), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1012), .A2(new_n730), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1044), .B1(new_n1045), .B2(KEYINPUT117), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1012), .A2(new_n1047), .A3(new_n730), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n1051));
  INV_X1    g626(.A(G8), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1051), .B1(G166), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1050), .A2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1054), .B(KEYINPUT119), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1049), .A2(G8), .A3(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(G8), .B1(new_n984), .B2(new_n979), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n578), .A2(G1976), .A3(new_n579), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(KEYINPUT52), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1006), .A2(new_n1018), .ZN(new_n1061));
  INV_X1    g636(.A(G1976), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT52), .B1(G288), .B2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1061), .A2(new_n1063), .A3(G8), .A4(new_n1058), .ZN(new_n1064));
  NAND2_X1  g639(.A1(G305), .A2(G1981), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n1066));
  INV_X1    g641(.A(G1981), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n585), .A2(new_n1067), .A3(new_n586), .A4(new_n587), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1065), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT49), .ZN(new_n1070));
  NAND3_X1  g645(.A1(G305), .A2(KEYINPUT120), .A3(G1981), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1072), .A2(G8), .A3(new_n1061), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1070), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1060), .B(new_n1064), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n1012), .A2(new_n730), .ZN(new_n1076));
  OR2_X1    g651(.A1(new_n1018), .A2(new_n1015), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n1006), .A3(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1079), .A2(G2090), .ZN(new_n1080));
  OAI21_X1  g655(.A(G8), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1054), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1075), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G1966), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1008), .B1(new_n1018), .B2(KEYINPUT45), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1084), .B1(new_n1085), .B2(new_n984), .ZN(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT121), .B(G2084), .Z(new_n1087));
  NAND4_X1  g662(.A1(new_n1006), .A2(new_n1022), .A3(new_n1016), .A4(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1086), .A2(new_n1088), .A3(G168), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(G8), .ZN(new_n1090));
  AOI21_X1  g665(.A(G168), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT51), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT51), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1089), .A2(new_n1093), .A3(G8), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1043), .A2(new_n1056), .A3(new_n1083), .A4(new_n1095), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n1025), .A2(new_n1039), .A3(G171), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1013), .A2(new_n1024), .A3(new_n1041), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(G171), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT54), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1003), .B1(new_n1096), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1056), .A2(new_n1083), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1042), .A2(KEYINPUT54), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1105), .A2(new_n1040), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1100), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1107), .B1(new_n1108), .B2(new_n1097), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1104), .A2(new_n1106), .A3(KEYINPUT127), .A4(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G1956), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1079), .A2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT56), .B(G2072), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1037), .A2(new_n1006), .A3(new_n1011), .A4(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n565), .B(new_n567), .C1(KEYINPUT123), .C2(KEYINPUT57), .ZN(new_n1116));
  NAND2_X1  g691(.A1(KEYINPUT123), .A2(KEYINPUT57), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1116), .B(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(G1348), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1021), .A2(new_n1121), .A3(new_n1023), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1006), .A2(new_n987), .A3(new_n1018), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n909), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1118), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1120), .A2(new_n1125), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  XOR2_X1   g704(.A(KEYINPUT58), .B(G1341), .Z(new_n1130));
  NAND2_X1  g705(.A1(new_n1061), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1131), .B1(new_n1012), .B2(G1996), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1132), .A2(KEYINPUT59), .A3(new_n556), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT59), .B1(new_n1132), .B2(new_n556), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT60), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1122), .A2(new_n1136), .A3(new_n604), .A4(new_n1123), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1120), .A2(KEYINPUT61), .A3(new_n1125), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1129), .A2(new_n1135), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1124), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1122), .A2(new_n909), .A3(new_n1123), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1136), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1120), .B(new_n1126), .C1(new_n1139), .C2(new_n1142), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1102), .A2(new_n1110), .A3(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n578), .A2(new_n1062), .A3(new_n579), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1068), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1147), .A2(G8), .A3(new_n1061), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1148), .B1(new_n1056), .B2(new_n1075), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1095), .A2(KEYINPUT62), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1150), .A2(new_n1103), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1100), .B1(new_n1095), .B2(KEYINPUT62), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1149), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT63), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1155), .A2(G8), .A3(new_n575), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1154), .B1(new_n1103), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1075), .A2(new_n1156), .A3(new_n1154), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1056), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1054), .B1(new_n1049), .B2(G8), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1158), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1161), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1163), .A2(KEYINPUT122), .A3(new_n1056), .A4(new_n1159), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1157), .A2(new_n1162), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1153), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1002), .B1(new_n1144), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n985), .B1(new_n989), .B2(new_n821), .ZN(new_n1168));
  NOR3_X1   g743(.A1(new_n998), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT46), .ZN(new_n1170));
  INV_X1    g745(.A(G1996), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1170), .B1(new_n985), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1168), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT47), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n998), .A2(G1986), .A3(G290), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1175), .B(KEYINPUT48), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1174), .B1(new_n1000), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(new_n705), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n997), .A2(new_n710), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n998), .B1(new_n1179), .B2(new_n988), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1167), .A2(new_n1181), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g757(.A1(new_n653), .A2(G227), .A3(new_n463), .A4(new_n462), .ZN(new_n1184));
  AND3_X1   g758(.A1(new_n694), .A2(new_n695), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g759(.A1(new_n1185), .A2(new_n894), .ZN(new_n1186));
  NOR2_X1   g760(.A1(new_n961), .A2(new_n1186), .ZN(G308));
  OR2_X1    g761(.A1(new_n961), .A2(new_n1186), .ZN(G225));
endmodule


