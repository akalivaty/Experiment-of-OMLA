//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 0 1 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1357, new_n1358, new_n1359;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT64), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n206), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n209), .B(new_n215), .C1(new_n222), .C2(KEYINPUT1), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XOR2_X1   g0024(.A(G250), .B(G257), .Z(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT65), .ZN(new_n226));
  XNOR2_X1  g0026(.A(G264), .B(G270), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n228), .B(new_n233), .Z(G358));
  XNOR2_X1  g0034(.A(G68), .B(G77), .ZN(new_n235));
  INV_X1    g0035(.A(G58), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT66), .B(G50), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(G1), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n244), .A2(G13), .A3(G20), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n212), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n244), .A2(G20), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n249), .A2(G50), .A3(new_n250), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(G50), .B2(new_n245), .ZN(new_n252));
  INV_X1    g0052(.A(new_n248), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT8), .B(G58), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n213), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT67), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n213), .A2(KEYINPUT67), .A3(G33), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n255), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n253), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n252), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(KEYINPUT9), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n265), .B(KEYINPUT74), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT3), .B(G33), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n267), .A2(G223), .A3(G1698), .ZN(new_n268));
  INV_X1    g0068(.A(G77), .ZN(new_n269));
  INV_X1    g0069(.A(G1698), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G222), .ZN(new_n272));
  OAI221_X1 g0072(.A(new_n268), .B1(new_n269), .B2(new_n267), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G41), .ZN(new_n276));
  INV_X1    g0076(.A(G45), .ZN(new_n277));
  AOI21_X1  g0077(.A(G1), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G1), .A3(G13), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n278), .A2(new_n280), .A3(G274), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n244), .B1(G41), .B2(G45), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n282), .B1(G226), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n275), .A2(new_n286), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n287), .A2(G200), .B1(new_n264), .B2(KEYINPUT9), .ZN(new_n288));
  INV_X1    g0088(.A(G190), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n266), .B(new_n288), .C1(new_n289), .C2(new_n287), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n290), .B(KEYINPUT10), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n287), .A2(G179), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT68), .ZN(new_n293));
  INV_X1    g0093(.A(G169), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n264), .B1(new_n287), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n249), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n255), .A2(new_n250), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n298), .A2(new_n299), .B1(new_n245), .B2(new_n255), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT76), .ZN(new_n301));
  AND2_X1   g0101(.A1(KEYINPUT3), .A2(G33), .ZN(new_n302));
  NOR2_X1   g0102(.A1(KEYINPUT3), .A2(G33), .ZN(new_n303));
  NOR3_X1   g0103(.A1(new_n302), .A2(new_n303), .A3(G20), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n301), .B1(new_n304), .B2(KEYINPUT7), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT3), .ZN(new_n306));
  INV_X1    g0106(.A(G33), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(KEYINPUT3), .A2(G33), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n308), .A2(KEYINPUT7), .A3(new_n213), .A4(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT77), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n302), .A2(new_n303), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT77), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n312), .A2(new_n313), .A3(KEYINPUT7), .A4(new_n213), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n308), .A2(new_n213), .A3(new_n309), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT7), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(KEYINPUT76), .A3(new_n316), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n305), .A2(new_n311), .A3(new_n314), .A4(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G68), .ZN(new_n319));
  INV_X1    g0119(.A(G68), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n236), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(G20), .B1(new_n321), .B2(new_n201), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n261), .A2(G159), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT16), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n253), .B1(new_n319), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n315), .A2(new_n316), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT78), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(new_n329), .A3(new_n310), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n304), .A2(KEYINPUT78), .A3(KEYINPUT7), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n330), .A2(G68), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n324), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT16), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n300), .B1(new_n327), .B2(new_n335), .ZN(new_n336));
  OAI211_X1 g0136(.A(G226), .B(G1698), .C1(new_n302), .C2(new_n303), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT79), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT79), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n267), .A2(new_n339), .A3(G226), .A4(G1698), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(G223), .B(new_n270), .C1(new_n302), .C2(new_n303), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G33), .A2(G87), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n280), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n280), .A2(G232), .A3(new_n283), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n281), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT80), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT80), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n281), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(G169), .B1(new_n346), .B2(new_n352), .ZN(new_n353));
  AND3_X1   g0153(.A1(new_n281), .A2(new_n347), .A3(new_n350), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n350), .B1(new_n281), .B2(new_n347), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n344), .B1(new_n340), .B2(new_n338), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n356), .B(G179), .C1(new_n357), .C2(new_n280), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT18), .B1(new_n336), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT18), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n353), .A2(new_n358), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT16), .B1(new_n332), .B2(new_n324), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n325), .B1(new_n318), .B2(G68), .ZN(new_n364));
  NOR3_X1   g0164(.A1(new_n363), .A2(new_n364), .A3(new_n253), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n361), .B(new_n362), .C1(new_n365), .C2(new_n300), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n360), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n319), .A2(new_n326), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n335), .A2(new_n368), .A3(new_n248), .ZN(new_n369));
  INV_X1    g0169(.A(new_n300), .ZN(new_n370));
  INV_X1    g0170(.A(G200), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n346), .B2(new_n352), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n356), .B(new_n289), .C1(new_n357), .C2(new_n280), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AND4_X1   g0174(.A1(KEYINPUT17), .A2(new_n369), .A3(new_n370), .A4(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT17), .B1(new_n336), .B2(new_n374), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n367), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n230), .A2(G1698), .ZN(new_n380));
  OAI221_X1 g0180(.A(new_n380), .B1(G226), .B2(G1698), .C1(new_n302), .C2(new_n303), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G33), .A2(G97), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n274), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT13), .ZN(new_n385));
  INV_X1    g0185(.A(G274), .ZN(new_n386));
  AND2_X1   g0186(.A1(G1), .A2(G13), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n386), .B1(new_n387), .B2(new_n279), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n285), .A2(G238), .B1(new_n278), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n384), .A2(new_n385), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n280), .B1(new_n381), .B2(new_n382), .ZN(new_n391));
  INV_X1    g0191(.A(G238), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n281), .B1(new_n392), .B2(new_n284), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT13), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G200), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n390), .A2(G190), .A3(new_n394), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n258), .A2(G77), .A3(new_n259), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n261), .A2(G50), .B1(G20), .B2(new_n320), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT11), .B1(new_n401), .B2(new_n248), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n401), .A2(KEYINPUT11), .A3(new_n248), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(KEYINPUT75), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT75), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT11), .ZN(new_n407));
  AOI211_X1 g0207(.A(new_n407), .B(new_n253), .C1(new_n399), .C2(new_n400), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n406), .B1(new_n402), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n246), .A2(new_n320), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n410), .B(KEYINPUT12), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n249), .A2(G68), .A3(new_n250), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n405), .A2(new_n409), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n398), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n395), .A2(G169), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT14), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n390), .A2(G179), .A3(new_n394), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT14), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n385), .B1(new_n384), .B2(new_n389), .ZN(new_n419));
  NOR3_X1   g0219(.A1(new_n391), .A2(new_n393), .A3(KEYINPUT13), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n418), .B(G169), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n416), .A2(new_n417), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n414), .B1(new_n413), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(G244), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n281), .B1(new_n424), .B2(new_n284), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n267), .A2(G238), .A3(G1698), .ZN(new_n426));
  OR2_X1    g0226(.A1(KEYINPUT69), .A2(G107), .ZN(new_n427));
  NAND2_X1  g0227(.A1(KEYINPUT69), .A2(G107), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n312), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n426), .B(new_n430), .C1(new_n271), .C2(new_n230), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n425), .B1(new_n431), .B2(new_n274), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n432), .A2(new_n371), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(G190), .B2(new_n432), .ZN(new_n434));
  INV_X1    g0234(.A(new_n261), .ZN(new_n435));
  OAI22_X1  g0235(.A1(new_n254), .A2(new_n435), .B1(new_n213), .B2(new_n269), .ZN(new_n436));
  XNOR2_X1  g0236(.A(KEYINPUT15), .B(G87), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n437), .A2(new_n256), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n248), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT70), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT70), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n441), .B(new_n248), .C1(new_n436), .C2(new_n438), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT72), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n245), .A2(G77), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n445), .B(KEYINPUT71), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n269), .B1(new_n244), .B2(G20), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n446), .B1(new_n249), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n443), .A2(new_n444), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n443), .A2(new_n448), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT72), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n434), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT73), .ZN(new_n454));
  INV_X1    g0254(.A(new_n432), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n454), .B1(new_n455), .B2(G179), .ZN(new_n456));
  INV_X1    g0256(.A(G179), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n432), .A2(KEYINPUT73), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n455), .A2(new_n294), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n444), .B1(new_n443), .B2(new_n448), .ZN(new_n461));
  INV_X1    g0261(.A(new_n449), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n459), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n423), .A2(new_n453), .A3(new_n463), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n297), .A2(new_n379), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n267), .A2(new_n213), .A3(G87), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT22), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT22), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n267), .A2(new_n469), .A3(new_n213), .A4(G87), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n213), .A2(KEYINPUT23), .A3(G107), .ZN(new_n472));
  NAND2_X1  g0272(.A1(G33), .A2(G116), .ZN(new_n473));
  OAI21_X1  g0273(.A(KEYINPUT91), .B1(new_n473), .B2(G20), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT91), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n475), .A2(new_n213), .A3(G33), .A4(G116), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n472), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n427), .A2(G20), .A3(new_n428), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT23), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n477), .A2(new_n479), .A3(KEYINPUT92), .ZN(new_n480));
  AOI21_X1  g0280(.A(KEYINPUT92), .B1(new_n477), .B2(new_n479), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n471), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT24), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT24), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n484), .B(new_n471), .C1(new_n480), .C2(new_n481), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n248), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n267), .A2(G257), .A3(G1698), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n267), .A2(G250), .A3(new_n270), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G294), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n276), .A2(KEYINPUT5), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n244), .B(G45), .C1(new_n276), .C2(KEYINPUT5), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(new_n274), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n491), .A2(new_n274), .B1(new_n496), .B2(G264), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT83), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n494), .A2(KEYINPUT82), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n277), .A2(G1), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT82), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G41), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n500), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n280), .A2(G274), .A3(new_n492), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n498), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n506), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n508), .A2(KEYINPUT83), .A3(new_n504), .A4(new_n499), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n497), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n371), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(G190), .B2(new_n511), .ZN(new_n513));
  INV_X1    g0313(.A(G107), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n246), .A2(KEYINPUT25), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(KEYINPUT25), .B1(new_n246), .B2(new_n514), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n244), .A2(G33), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n245), .A2(new_n518), .A3(new_n212), .A4(new_n247), .ZN(new_n519));
  OAI22_X1  g0319(.A1(new_n516), .A2(new_n517), .B1(new_n514), .B2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n487), .A2(new_n513), .A3(new_n521), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n497), .A2(new_n510), .A3(new_n457), .ZN(new_n523));
  AOI21_X1  g0323(.A(G169), .B1(new_n497), .B2(new_n510), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n253), .B1(new_n483), .B2(new_n485), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n525), .B1(new_n526), .B2(new_n520), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n280), .A2(G274), .A3(new_n500), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT86), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n388), .A2(KEYINPUT86), .A3(new_n500), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n424), .A2(G1698), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(G238), .B2(G1698), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n473), .B1(new_n534), .B2(new_n312), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n274), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n280), .B(G250), .C1(G1), .C2(new_n277), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n532), .A2(new_n536), .A3(G190), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT87), .ZN(new_n539));
  INV_X1    g0339(.A(G250), .ZN(new_n540));
  NOR3_X1   g0340(.A1(new_n274), .A2(new_n540), .A3(new_n500), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n541), .B1(new_n535), .B2(new_n274), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT87), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n542), .A2(new_n543), .A3(G190), .A4(new_n532), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT88), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT88), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n539), .A2(new_n547), .A3(new_n544), .ZN(new_n548));
  INV_X1    g0348(.A(new_n437), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n549), .A2(new_n245), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT19), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n213), .B1(new_n382), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(G87), .ZN(new_n553));
  INV_X1    g0353(.A(G97), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n552), .B1(new_n429), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n267), .A2(new_n213), .A3(G68), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n551), .B1(new_n256), .B2(new_n554), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n550), .B1(new_n559), .B2(new_n248), .ZN(new_n560));
  OR2_X1    g0360(.A1(new_n519), .A2(new_n553), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n371), .B1(new_n542), .B2(new_n532), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n546), .A2(new_n548), .A3(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(G238), .A2(G1698), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n566), .B1(new_n424), .B2(G1698), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n567), .A2(new_n267), .B1(G33), .B2(G116), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n537), .B1(new_n568), .B2(new_n280), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n530), .A2(new_n531), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n457), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n560), .B1(new_n437), .B2(new_n519), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n542), .A2(new_n532), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n294), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n572), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n522), .A2(new_n527), .A3(new_n565), .A4(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(G244), .B(new_n270), .C1(new_n302), .C2(new_n303), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT4), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(G33), .A2(G283), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n579), .A2(new_n424), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n267), .A2(new_n270), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(G250), .B(G1698), .C1(new_n302), .C2(new_n303), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT81), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n267), .A2(KEYINPUT81), .A3(G250), .A4(G1698), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n274), .B1(new_n584), .B2(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(G257), .B(new_n280), .C1(new_n493), .C2(new_n494), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n590), .A2(new_n510), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT85), .ZN(new_n593));
  INV_X1    g0393(.A(new_n591), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n594), .B1(new_n507), .B2(new_n509), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT85), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n596), .A3(new_n590), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n593), .A2(G190), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n246), .A2(new_n554), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n519), .B2(new_n554), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n330), .A2(new_n331), .A3(new_n429), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n514), .A2(KEYINPUT6), .A3(G97), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n554), .A2(new_n514), .ZN(new_n603));
  NOR2_X1   g0403(.A1(G97), .A2(G107), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n602), .B1(new_n605), .B2(KEYINPUT6), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n606), .A2(G20), .B1(G77), .B2(new_n261), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n601), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n600), .B1(new_n608), .B2(new_n248), .ZN(new_n609));
  AOI21_X1  g0409(.A(KEYINPUT84), .B1(new_n592), .B2(G200), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n592), .A2(KEYINPUT84), .A3(G200), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n598), .B(new_n609), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n595), .A2(new_n596), .A3(new_n590), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n596), .B1(new_n595), .B2(new_n590), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n294), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n595), .A2(new_n457), .A3(new_n590), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n616), .A2(new_n609), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  OAI211_X1 g0418(.A(G270), .B(new_n280), .C1(new_n493), .C2(new_n494), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n267), .A2(G257), .A3(new_n270), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n267), .A2(G264), .A3(G1698), .ZN(new_n621));
  INV_X1    g0421(.A(G303), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n620), .B(new_n621), .C1(new_n622), .C2(new_n267), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n274), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n510), .A2(new_n619), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(G200), .ZN(new_n626));
  INV_X1    g0426(.A(G116), .ZN(new_n627));
  OR3_X1    g0427(.A1(new_n519), .A2(KEYINPUT89), .A3(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT89), .B1(new_n519), .B2(new_n627), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n627), .A2(G20), .ZN(new_n631));
  INV_X1    g0431(.A(G13), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n631), .A2(G1), .A3(new_n632), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n581), .B(new_n213), .C1(G33), .C2(new_n554), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(new_n248), .A3(new_n631), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT20), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n634), .A2(KEYINPUT20), .A3(new_n248), .A4(new_n631), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n633), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n626), .A2(KEYINPUT90), .A3(new_n630), .A4(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT90), .ZN(new_n641));
  INV_X1    g0441(.A(new_n619), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n507), .B2(new_n509), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n371), .B1(new_n643), .B2(new_n624), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n630), .A2(new_n639), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n641), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n643), .A2(G190), .A3(new_n624), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n640), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n625), .A2(KEYINPUT21), .A3(new_n645), .A4(G169), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n457), .B1(new_n623), .B2(new_n274), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n645), .A2(new_n643), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n294), .B1(new_n643), .B2(new_n624), .ZN(new_n653));
  AOI21_X1  g0453(.A(KEYINPUT21), .B1(new_n653), .B2(new_n645), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n612), .A2(new_n618), .A3(new_n648), .A4(new_n655), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n466), .A2(new_n577), .A3(new_n656), .ZN(G372));
  AOI21_X1  g0457(.A(new_n253), .B1(new_n601), .B2(new_n607), .ZN(new_n658));
  OAI22_X1  g0458(.A1(new_n592), .A2(G179), .B1(new_n658), .B2(new_n600), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n593), .A2(new_n597), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n294), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n661), .A2(KEYINPUT26), .A3(new_n565), .A4(new_n576), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n564), .A2(new_n545), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n615), .A2(new_n617), .A3(new_n576), .A4(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n654), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n649), .A2(new_n651), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n527), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n520), .B1(new_n486), .B2(new_n248), .ZN(new_n671));
  AOI22_X1  g0471(.A1(new_n671), .A2(new_n513), .B1(new_n545), .B2(new_n564), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n670), .A2(new_n672), .A3(new_n618), .A4(new_n612), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n667), .A2(new_n673), .A3(new_n576), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n465), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT93), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n421), .A2(new_n417), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n418), .B1(new_n395), .B2(G169), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n413), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n463), .B2(new_n414), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n377), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n367), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n291), .A2(new_n682), .B1(new_n293), .B2(new_n295), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n676), .A2(new_n683), .ZN(G369));
  AND2_X1   g0484(.A1(new_n648), .A2(new_n655), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n632), .A2(G1), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n213), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT27), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n686), .A2(new_n689), .A3(new_n213), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n688), .A2(G213), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G343), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT94), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n645), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n694), .B(KEYINPUT95), .Z(new_n695));
  NAND2_X1  g0495(.A1(new_n685), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n655), .B2(new_n695), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n522), .A2(new_n527), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n692), .B(KEYINPUT94), .Z(new_n700));
  NOR2_X1   g0500(.A1(new_n671), .A2(new_n700), .ZN(new_n701));
  OAI22_X1  g0501(.A1(new_n699), .A2(new_n701), .B1(new_n527), .B2(new_n700), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n669), .A2(new_n668), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n700), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n699), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n527), .A2(new_n693), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n703), .A2(new_n709), .ZN(G399));
  INV_X1    g0510(.A(new_n207), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(G41), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n211), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n244), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  OR3_X1    g0515(.A1(new_n429), .A2(G116), .A3(new_n555), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n713), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT28), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT31), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n613), .A2(new_n614), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n571), .A2(new_n643), .A3(new_n497), .A4(new_n650), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n511), .A2(new_n457), .A3(new_n574), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n592), .A2(new_n625), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n720), .A2(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n722), .B1(new_n660), .B2(new_n721), .ZN(new_n727));
  AOI211_X1 g0527(.A(new_n719), .B(new_n700), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  AND4_X1   g0528(.A1(new_n497), .A2(new_n571), .A3(new_n643), .A4(new_n650), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n729), .A2(new_n593), .A3(KEYINPUT30), .A4(new_n597), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n571), .A2(G179), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n731), .A2(new_n511), .A3(new_n592), .A4(new_n625), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n613), .A2(new_n721), .A3(new_n614), .ZN(new_n733));
  OAI211_X1 g0533(.A(new_n730), .B(new_n732), .C1(new_n733), .C2(KEYINPUT30), .ZN(new_n734));
  AOI21_X1  g0534(.A(KEYINPUT31), .B1(new_n734), .B2(new_n693), .ZN(new_n735));
  OAI21_X1  g0535(.A(KEYINPUT96), .B1(new_n728), .B2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(KEYINPUT30), .B1(new_n720), .B2(new_n729), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n496), .A2(G264), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n491), .A2(new_n274), .ZN(new_n739));
  AND4_X1   g0539(.A1(new_n738), .A2(new_n739), .A3(new_n542), .A4(new_n532), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n740), .A2(KEYINPUT30), .A3(new_n643), .A4(new_n650), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n732), .B1(new_n660), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n693), .B1(new_n737), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n719), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT96), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n693), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n577), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n612), .A2(new_n618), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n748), .A2(new_n749), .A3(new_n685), .A4(new_n700), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n736), .A2(new_n747), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G330), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT97), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n751), .A2(KEYINPUT97), .A3(G330), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(KEYINPUT29), .B1(new_n674), .B2(new_n700), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n673), .A2(new_n576), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n664), .A2(new_n665), .ZN(new_n759));
  INV_X1    g0559(.A(new_n576), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n560), .B(new_n561), .C1(new_n571), .C2(new_n371), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n761), .B1(new_n545), .B2(KEYINPUT88), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n760), .B1(new_n762), .B2(new_n548), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n661), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n759), .B1(new_n665), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n758), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n693), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n757), .B1(new_n767), .B2(KEYINPUT29), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n756), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n718), .B1(new_n769), .B2(G1), .ZN(G364));
  NOR3_X1   g0570(.A1(new_n632), .A2(new_n277), .A3(G20), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT98), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n715), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n698), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(G330), .B2(new_n697), .ZN(new_n775));
  INV_X1    g0575(.A(new_n773), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n213), .A2(new_n457), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n289), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT102), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(KEYINPUT103), .B(G326), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G190), .A2(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n777), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G311), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n213), .A2(G179), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n784), .ZN(new_n788));
  INV_X1    g0588(.A(G329), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n785), .A2(new_n786), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n777), .A2(G190), .A3(new_n371), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n267), .B(new_n790), .C1(G322), .C2(new_n792), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n289), .A2(G179), .A3(G200), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n213), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n778), .A2(G190), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT33), .B(G317), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G294), .A2(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n787), .A2(G190), .A3(G200), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n787), .A2(new_n289), .A3(G200), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n801), .A2(G303), .B1(new_n803), .B2(G283), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n783), .A2(new_n793), .A3(new_n799), .A4(new_n804), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n791), .A2(new_n236), .B1(new_n785), .B2(new_n269), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(G68), .B2(new_n797), .ZN(new_n807));
  INV_X1    g0607(.A(G159), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n788), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT32), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n779), .A2(G50), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n796), .A2(G97), .B1(new_n803), .B2(G107), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n807), .A2(new_n810), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n267), .B1(new_n800), .B2(new_n553), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT101), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n805), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n212), .B1(G20), .B2(new_n294), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n776), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n711), .A2(new_n267), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(new_n277), .B2(new_n211), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n239), .B2(new_n277), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n711), .A2(new_n312), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT99), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n824), .A2(G355), .B1(new_n627), .B2(new_n711), .ZN(new_n825));
  AOI21_X1  g0625(.A(KEYINPUT100), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n822), .A2(KEYINPUT100), .A3(new_n825), .ZN(new_n827));
  NOR2_X1   g0627(.A1(G13), .A2(G33), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(G20), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(new_n817), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n830), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n818), .B1(new_n826), .B2(new_n832), .C1(new_n697), .C2(new_n833), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n775), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(G396));
  INV_X1    g0636(.A(new_n756), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n674), .A2(new_n700), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n700), .B1(new_n451), .B2(new_n449), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n463), .B1(new_n452), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n462), .A2(new_n461), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n842), .A2(new_n459), .A3(new_n460), .A4(new_n700), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n838), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n844), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n674), .A2(new_n846), .A3(new_n700), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n773), .B1(new_n837), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n837), .B2(new_n848), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n817), .A2(new_n828), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n773), .B1(G77), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n779), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n854), .A2(new_n622), .B1(new_n800), .B2(new_n514), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(G87), .B2(new_n803), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n267), .B1(new_n792), .B2(G294), .ZN(new_n857));
  INV_X1    g0657(.A(new_n785), .ZN(new_n858));
  INV_X1    g0658(.A(new_n788), .ZN(new_n859));
  AOI22_X1  g0659(.A1(G116), .A2(new_n858), .B1(new_n859), .B2(G311), .ZN(new_n860));
  AOI22_X1  g0660(.A1(G97), .A2(new_n796), .B1(new_n797), .B2(G283), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n856), .A2(new_n857), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n792), .A2(G143), .B1(new_n858), .B2(G159), .ZN(new_n863));
  INV_X1    g0663(.A(G137), .ZN(new_n864));
  INV_X1    g0664(.A(G150), .ZN(new_n865));
  INV_X1    g0665(.A(new_n797), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n863), .B1(new_n854), .B2(new_n864), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT34), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(G132), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n267), .B1(new_n788), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(G68), .B2(new_n803), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n796), .A2(G58), .B1(new_n801), .B2(G50), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n869), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n867), .A2(new_n868), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n862), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n853), .B1(new_n876), .B2(new_n817), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(new_n846), .B2(new_n829), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n850), .A2(new_n878), .ZN(G384));
  OAI21_X1  g0679(.A(G1), .B1(new_n632), .B2(G20), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n413), .A2(new_n693), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n679), .B(new_n881), .C1(new_n413), .C2(new_n398), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n413), .B(new_n693), .C1(new_n677), .C2(new_n678), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n884), .A2(new_n843), .A3(new_n840), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n728), .A2(new_n735), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n885), .B1(new_n886), .B2(new_n750), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT40), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT105), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n375), .B2(new_n376), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n369), .A2(new_n370), .A3(new_n374), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT17), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n336), .A2(KEYINPUT17), .A3(new_n374), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n893), .A2(KEYINPUT105), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n890), .A2(new_n367), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n691), .B1(new_n365), .B2(new_n300), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n362), .B1(new_n365), .B2(new_n300), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(new_n897), .A3(new_n891), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT37), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT37), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n900), .A2(new_n897), .A3(new_n903), .A4(new_n891), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n899), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT38), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n906), .A2(KEYINPUT106), .A3(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT106), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n896), .A2(new_n898), .B1(new_n904), .B2(new_n902), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n909), .B1(new_n910), .B2(KEYINPUT38), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT104), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n315), .A2(KEYINPUT76), .A3(new_n316), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT76), .B1(new_n315), .B2(new_n316), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n311), .A2(new_n314), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n320), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n324), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n334), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n300), .B1(new_n920), .B2(new_n327), .ZN(new_n921));
  INV_X1    g0721(.A(new_n691), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n913), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n248), .B1(new_n918), .B2(new_n325), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT16), .B1(new_n319), .B2(new_n324), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n370), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(KEYINPUT104), .A3(new_n691), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n362), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n923), .A2(new_n927), .A3(new_n891), .A4(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT37), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n904), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n923), .A2(new_n927), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n378), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n931), .A2(new_n933), .A3(KEYINPUT38), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n888), .B1(new_n912), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT40), .ZN(new_n936));
  INV_X1    g0736(.A(new_n904), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(KEYINPUT37), .B2(new_n929), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n367), .A2(new_n377), .B1(new_n923), .B2(new_n927), .ZN(new_n939));
  NOR3_X1   g0739(.A1(new_n938), .A2(new_n907), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT38), .B1(new_n931), .B2(new_n933), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n887), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n935), .B1(new_n936), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n744), .A2(new_n746), .ZN(new_n944));
  NOR3_X1   g0744(.A1(new_n656), .A2(new_n577), .A3(new_n693), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n466), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(G330), .B1(new_n943), .B2(new_n947), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n948), .B1(new_n949), .B2(KEYINPUT107), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(KEYINPUT107), .B2(new_n949), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT39), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n907), .B1(new_n938), .B2(new_n939), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n952), .B1(new_n953), .B2(new_n934), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n934), .A2(new_n952), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n954), .B1(new_n912), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n422), .A2(new_n413), .A3(new_n700), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n847), .A2(new_n843), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n884), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n953), .A2(new_n934), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n960), .A2(new_n962), .B1(new_n367), .B2(new_n691), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n958), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n768), .A2(new_n465), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n683), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n964), .B(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n880), .B1(new_n951), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(new_n967), .B2(new_n951), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n606), .A2(KEYINPUT35), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n606), .A2(KEYINPUT35), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n970), .A2(G116), .A3(new_n214), .A4(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT36), .Z(new_n973));
  OAI211_X1 g0773(.A(new_n211), .B(G77), .C1(new_n236), .C2(new_n320), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n202), .A2(G68), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n244), .B(G13), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  OR3_X1    g0776(.A1(new_n969), .A2(new_n973), .A3(new_n976), .ZN(G367));
  AOI22_X1  g0777(.A1(new_n796), .A2(new_n429), .B1(new_n803), .B2(G97), .ZN(new_n978));
  INV_X1    g0778(.A(G294), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n978), .B1(new_n979), .B2(new_n866), .C1(new_n780), .C2(new_n786), .ZN(new_n980));
  AND3_X1   g0780(.A1(new_n801), .A2(KEYINPUT46), .A3(G116), .ZN(new_n981));
  AOI21_X1  g0781(.A(KEYINPUT46), .B1(new_n801), .B2(G116), .ZN(new_n982));
  AOI22_X1  g0782(.A1(G283), .A2(new_n858), .B1(new_n859), .B2(G317), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n983), .B(new_n312), .C1(new_n622), .C2(new_n791), .ZN(new_n984));
  NOR4_X1   g0784(.A1(new_n980), .A2(new_n981), .A3(new_n982), .A4(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT111), .Z(new_n986));
  NAND2_X1  g0786(.A1(new_n781), .A2(G143), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n791), .A2(new_n865), .B1(new_n788), .B2(new_n864), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n312), .B(new_n988), .C1(G50), .C2(new_n858), .ZN(new_n989));
  AOI22_X1  g0789(.A1(G68), .A2(new_n796), .B1(new_n797), .B2(G159), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n801), .A2(G58), .B1(new_n803), .B2(G77), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n987), .A2(new_n989), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n986), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT47), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n817), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n228), .A2(new_n819), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n817), .B(new_n830), .C1(new_n711), .C2(new_n549), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n776), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n760), .A2(new_n562), .A3(new_n693), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n693), .A2(new_n562), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n663), .A2(new_n1000), .A3(new_n576), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n995), .B(new_n998), .C1(new_n833), .C2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n772), .A2(new_n244), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n703), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n749), .B1(new_n609), .B2(new_n700), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n661), .A2(new_n693), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g0810(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  AND3_X1   g0812(.A1(new_n1010), .A2(new_n709), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1012), .B1(new_n1010), .B2(new_n709), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT44), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n1010), .B2(new_n709), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n1013), .A2(new_n1014), .B1(new_n1016), .B2(KEYINPUT110), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n705), .A2(new_n699), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n707), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1019), .A2(KEYINPUT44), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1020));
  AND3_X1   g0820(.A1(new_n1016), .A2(new_n1020), .A3(KEYINPUT110), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1007), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1016), .A2(KEYINPUT110), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1016), .A2(new_n1020), .A3(KEYINPUT110), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1023), .A2(new_n703), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1022), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n705), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1018), .B1(new_n702), .B2(new_n1028), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n698), .B(new_n1029), .Z(new_n1030));
  OAI21_X1  g0830(.A(new_n769), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n712), .B(new_n1032), .Z(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1006), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1010), .A2(new_n706), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1036), .A2(KEYINPUT42), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n618), .B1(new_n1008), .B2(new_n527), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1036), .A2(KEYINPUT42), .B1(new_n1038), .B2(new_n700), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n1037), .A2(new_n1039), .B1(KEYINPUT43), .B2(new_n1003), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(KEYINPUT43), .B2(new_n1003), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT43), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1037), .A2(new_n1039), .A3(new_n1042), .A4(new_n1002), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1010), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1044), .B1(new_n703), .B2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1041), .A2(new_n1007), .A3(new_n1010), .A4(new_n1043), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1004), .B1(new_n1035), .B2(new_n1048), .ZN(G387));
  NOR2_X1   g0849(.A1(new_n1030), .A2(new_n1005), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT112), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n702), .A2(new_n833), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n824), .A2(new_n716), .B1(new_n514), .B2(new_n711), .ZN(new_n1053));
  AOI211_X1 g0853(.A(G45), .B(new_n716), .C1(G68), .C2(G77), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n254), .A2(G50), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT50), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n819), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n233), .A2(new_n277), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1053), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT113), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1062), .A2(new_n831), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n773), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT114), .Z(new_n1066));
  OAI22_X1  g0866(.A1(new_n785), .A2(new_n320), .B1(new_n788), .B2(new_n865), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n312), .B(new_n1067), .C1(G50), .C2(new_n792), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n801), .A2(G77), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n549), .A2(new_n796), .B1(new_n797), .B2(new_n255), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n779), .A2(G159), .B1(new_n803), .B2(G97), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n781), .A2(G322), .B1(G311), .B2(new_n797), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1074), .A2(KEYINPUT115), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(KEYINPUT115), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n792), .A2(G317), .B1(new_n858), .B2(G303), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT48), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(G283), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n795), .A2(new_n1081), .B1(new_n800), .B2(new_n979), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1080), .A2(KEYINPUT49), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n267), .B1(new_n859), .B2(new_n782), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1084), .B(new_n1085), .C1(new_n627), .C2(new_n802), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT49), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1072), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1052), .B(new_n1066), .C1(new_n1088), .C2(new_n817), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1051), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1030), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n769), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n769), .A2(new_n1091), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n712), .B(KEYINPUT116), .Z(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1090), .B1(new_n1092), .B2(new_n1095), .ZN(G393));
  NAND3_X1  g0896(.A1(new_n1022), .A2(new_n1026), .A3(new_n1006), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n831), .B1(new_n554), .B2(new_n207), .C1(new_n242), .C2(new_n820), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n773), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n796), .A2(G77), .B1(new_n801), .B2(G68), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n797), .A2(G50), .B1(new_n803), .B2(G87), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n858), .A2(new_n255), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n312), .B1(new_n859), .B2(G143), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(G150), .A2(new_n779), .B1(new_n792), .B2(G159), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(KEYINPUT117), .B(KEYINPUT51), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1105), .B(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G317), .A2(new_n779), .B1(new_n792), .B2(G311), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT52), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(G116), .A2(new_n796), .B1(new_n797), .B2(G303), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n312), .B1(new_n785), .B2(new_n979), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(G322), .B2(new_n859), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n801), .A2(G283), .B1(new_n803), .B2(G107), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1110), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n1104), .A2(new_n1107), .B1(new_n1109), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1099), .B1(new_n1115), .B2(new_n817), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n1010), .B2(new_n833), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1094), .B1(new_n1093), .B2(new_n1027), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n769), .A2(new_n1091), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1097), .B(new_n1117), .C1(new_n1118), .C2(new_n1119), .ZN(G390));
  INV_X1    g0920(.A(new_n1094), .ZN(new_n1121));
  OAI21_X1  g0921(.A(G330), .B1(new_n944), .B2(new_n945), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n466), .A2(new_n1122), .ZN(new_n1123));
  OR2_X1    g0923(.A1(new_n966), .A2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1122), .A2(new_n885), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n844), .B1(new_n754), .B2(new_n755), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1126), .B1(new_n1127), .B2(new_n884), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n959), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n700), .B(new_n840), .C1(new_n758), .C2(new_n765), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n843), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n883), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n423), .B2(new_n881), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n1122), .B2(new_n844), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT118), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g0936(.A(KEYINPUT118), .B(new_n1133), .C1(new_n1122), .C2(new_n844), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1131), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n751), .A2(KEYINPUT97), .A3(G330), .ZN(new_n1139));
  AOI21_X1  g0939(.A(KEYINPUT97), .B1(new_n751), .B2(G330), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n846), .B(new_n884), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1124), .B1(new_n1129), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n960), .A2(new_n957), .ZN(new_n1144));
  AOI21_X1  g0944(.A(KEYINPUT106), .B1(new_n906), .B2(new_n907), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n910), .A2(new_n909), .A3(KEYINPUT38), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n955), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n954), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1144), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n912), .A2(new_n934), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1133), .B1(new_n1130), .B2(new_n843), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n957), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1149), .A2(new_n1154), .A3(new_n1141), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n956), .A2(new_n1144), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1155), .B1(new_n1156), .B2(new_n1126), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1121), .B1(new_n1143), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT119), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n934), .A2(new_n952), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n908), .B2(new_n911), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1152), .B1(new_n959), .B2(new_n884), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n1162), .A2(new_n1163), .A3(new_n954), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n940), .B1(new_n908), .B2(new_n911), .ZN(new_n1165));
  NOR3_X1   g0965(.A1(new_n1165), .A2(new_n1152), .A3(new_n1151), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1125), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n846), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1125), .B1(new_n1168), .B2(new_n1133), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n959), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1142), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n966), .A2(new_n1123), .ZN(new_n1172));
  AOI221_X4 g0972(.A(new_n1160), .B1(new_n1167), .B2(new_n1155), .C1(new_n1171), .C2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT119), .B1(new_n1174), .B2(new_n1157), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1159), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n956), .A2(new_n828), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n854), .A2(new_n1081), .B1(new_n269), .B2(new_n795), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n801), .A2(G87), .B1(new_n803), .B2(G68), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n792), .A2(G116), .B1(new_n859), .B2(G294), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n267), .B1(new_n858), .B2(G97), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1178), .B(new_n1182), .C1(new_n429), .C2(new_n797), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT120), .ZN(new_n1184));
  INV_X1    g0984(.A(G125), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n791), .A2(new_n870), .B1(new_n788), .B2(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(KEYINPUT54), .B(G143), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n312), .B(new_n1186), .C1(new_n858), .C2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(KEYINPUT53), .B1(new_n800), .B2(new_n865), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(G128), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n854), .A2(new_n1192), .B1(new_n802), .B2(new_n202), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n866), .A2(new_n864), .B1(new_n808), .B2(new_n795), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n800), .A2(KEYINPUT53), .A3(new_n865), .ZN(new_n1195));
  NOR4_X1   g0995(.A1(new_n1191), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n817), .B1(new_n1184), .B2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n776), .B1(new_n254), .B2(new_n851), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1177), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT121), .Z(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n1006), .B2(new_n1158), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1176), .A2(new_n1201), .ZN(G378));
  AOI22_X1  g1002(.A1(new_n1128), .A2(new_n959), .B1(new_n1141), .B2(new_n1138), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1172), .B1(new_n1203), .B2(new_n1157), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT122), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1133), .A2(new_n844), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n944), .B2(new_n945), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(new_n953), .B2(new_n934), .ZN(new_n1208));
  OAI21_X1  g1008(.A(G330), .B1(new_n1208), .B2(KEYINPUT40), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1205), .B1(new_n935), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(G330), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n942), .B2(new_n936), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1212), .B(KEYINPUT122), .C1(new_n1165), .C2(new_n888), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n291), .A2(new_n296), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n264), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1214), .A2(new_n1215), .A3(new_n691), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n291), .B(new_n296), .C1(new_n264), .C2(new_n922), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1218));
  AND3_X1   g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1218), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1210), .A2(new_n1213), .A3(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n935), .A2(new_n1209), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1224), .A2(KEYINPUT122), .A3(new_n1221), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n964), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1223), .A2(new_n964), .A3(new_n1225), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1204), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT57), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1204), .A2(new_n1228), .A3(KEYINPUT57), .A4(new_n1229), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1232), .A2(new_n1094), .A3(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1228), .A2(new_n1006), .A3(new_n1229), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n773), .B1(G50), .B2(new_n852), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n854), .A2(new_n627), .B1(new_n802), .B2(new_n236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G97), .B2(new_n797), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n312), .A2(new_n276), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(G283), .B2(new_n859), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n792), .A2(G107), .B1(new_n858), .B2(new_n549), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n796), .A2(G68), .B1(new_n801), .B2(G77), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1238), .A2(new_n1240), .A3(new_n1241), .A4(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT58), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1239), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n1185), .A2(new_n854), .B1(new_n866), .B2(new_n870), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n792), .A2(G128), .B1(new_n858), .B2(G137), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1249), .B1(new_n800), .B2(new_n1187), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n1248), .B(new_n1250), .C1(G150), .C2(new_n796), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(KEYINPUT59), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n803), .A2(G159), .ZN(new_n1254));
  AOI211_X1 g1054(.A(G33), .B(G41), .C1(new_n859), .C2(G124), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1252), .A2(KEYINPUT59), .ZN(new_n1257));
  OAI221_X1 g1057(.A(new_n1247), .B1(new_n1244), .B2(new_n1243), .C1(new_n1256), .C2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1236), .B1(new_n1258), .B2(new_n817), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1259), .B1(new_n1222), .B2(new_n829), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1235), .A2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1234), .A2(new_n1261), .ZN(G375));
  NAND3_X1  g1062(.A1(new_n1129), .A2(new_n1142), .A3(new_n1124), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1174), .A2(new_n1263), .A3(new_n1034), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1133), .A2(new_n828), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n773), .B1(G68), .B2(new_n852), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1266), .B(KEYINPUT123), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n627), .A2(new_n866), .B1(new_n854), .B2(new_n979), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(G97), .B2(new_n801), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n267), .B1(new_n792), .B2(G283), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n429), .A2(new_n858), .B1(new_n859), .B2(G303), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n796), .A2(new_n549), .B1(new_n803), .B2(G77), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1269), .A2(new_n1270), .A3(new_n1271), .A4(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n779), .A2(G132), .ZN(new_n1274));
  XOR2_X1   g1074(.A(new_n1274), .B(KEYINPUT124), .Z(new_n1275));
  AOI22_X1  g1075(.A1(new_n796), .A2(G50), .B1(new_n801), .B2(G159), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n797), .A2(new_n1188), .B1(new_n803), .B2(G58), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n312), .B1(new_n792), .B2(G137), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(G150), .A2(new_n858), .B1(new_n859), .B2(G128), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1276), .A2(new_n1277), .A3(new_n1278), .A4(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1273), .B1(new_n1275), .B2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1267), .B1(new_n1281), .B2(new_n817), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n1171), .A2(new_n1006), .B1(new_n1265), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1264), .A2(new_n1283), .ZN(G381));
  INV_X1    g1084(.A(G390), .ZN(new_n1285));
  INV_X1    g1085(.A(G384), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  OR4_X1    g1087(.A1(G396), .A2(new_n1287), .A3(G387), .A4(G393), .ZN(new_n1288));
  OR4_X1    g1088(.A1(G378), .A2(new_n1288), .A3(G375), .A4(G381), .ZN(G407));
  INV_X1    g1089(.A(G378), .ZN(new_n1290));
  INV_X1    g1090(.A(G343), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(G213), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1290), .A2(new_n1293), .ZN(new_n1294));
  OAI211_X1 g1094(.A(G407), .B(G213), .C1(G375), .C2(new_n1294), .ZN(G409));
  NAND2_X1  g1095(.A1(G387), .A2(new_n1285), .ZN(new_n1296));
  OAI211_X1 g1096(.A(G390), .B(new_n1004), .C1(new_n1035), .C2(new_n1048), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT126), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(KEYINPUT125), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(G393), .B(new_n835), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT125), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1298), .A2(new_n1303), .A3(new_n1299), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1301), .A2(new_n1302), .A3(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1302), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1303), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1307));
  AOI211_X1 g1107(.A(KEYINPUT125), .B(KEYINPUT126), .C1(new_n1296), .C2(new_n1297), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1306), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1305), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT61), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1234), .A2(G378), .A3(new_n1261), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1235), .B(new_n1260), .C1(new_n1230), .C2(new_n1033), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1313), .A2(new_n1176), .A3(new_n1201), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1293), .B1(new_n1312), .B2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT60), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1263), .A2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1203), .A2(KEYINPUT60), .A3(new_n1124), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1317), .A2(new_n1094), .A3(new_n1174), .A4(new_n1318), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1319), .A2(G384), .A3(new_n1283), .ZN(new_n1320));
  AOI21_X1  g1120(.A(G384), .B1(new_n1319), .B2(new_n1283), .ZN(new_n1321));
  OAI211_X1 g1121(.A(G2897), .B(new_n1293), .C1(new_n1320), .C2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1319), .A2(new_n1283), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(new_n1286), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1319), .A2(G384), .A3(new_n1283), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1293), .A2(G2897), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1324), .A2(new_n1325), .A3(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1322), .A2(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1311), .B1(new_n1315), .B2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT62), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1330), .B1(new_n1315), .B2(new_n1332), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1329), .A2(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1315), .A2(new_n1330), .A3(new_n1332), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1310), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1315), .A2(KEYINPUT63), .A3(new_n1332), .ZN(new_n1337));
  OAI211_X1 g1137(.A(new_n1337), .B(new_n1311), .C1(new_n1315), .C2(new_n1328), .ZN(new_n1338));
  AOI211_X1 g1138(.A(new_n1293), .B(new_n1331), .C1(new_n1312), .C2(new_n1314), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1310), .B1(new_n1339), .B2(KEYINPUT63), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1338), .A2(new_n1340), .ZN(new_n1341));
  OAI21_X1  g1141(.A(KEYINPUT127), .B1(new_n1336), .B2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1315), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1328), .ZN(new_n1344));
  AOI21_X1  g1144(.A(KEYINPUT61), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1315), .A2(new_n1332), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1346), .A2(KEYINPUT62), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1345), .A2(new_n1347), .A3(new_n1335), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1310), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT127), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT63), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1346), .A2(new_n1352), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1345), .A2(new_n1353), .A3(new_n1310), .A4(new_n1337), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1350), .A2(new_n1351), .A3(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1342), .A2(new_n1355), .ZN(G405));
  NAND2_X1  g1156(.A1(G375), .A2(new_n1290), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1357), .A2(new_n1312), .ZN(new_n1358));
  XNOR2_X1  g1158(.A(new_n1358), .B(new_n1331), .ZN(new_n1359));
  XNOR2_X1  g1159(.A(new_n1359), .B(new_n1310), .ZN(G402));
endmodule


