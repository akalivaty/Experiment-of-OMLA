//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n832, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(KEYINPUT16), .A3(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G8gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT101), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n204), .B(new_n206), .C1(new_n203), .C2(new_n202), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n205), .A2(KEYINPUT101), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT21), .ZN(new_n210));
  XNOR2_X1  g009(.A(G57gat), .B(G64gat), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G71gat), .B(G78gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n213), .B(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n209), .B1(new_n210), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n217), .B(G183gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(G231gat), .A2(G233gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n218), .B(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(KEYINPUT107), .B(KEYINPUT20), .Z(new_n221));
  XNOR2_X1  g020(.A(new_n220), .B(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n215), .A2(KEYINPUT21), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT108), .B(KEYINPUT19), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n224), .B(G211gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n223), .B(new_n225), .ZN(new_n226));
  XOR2_X1   g025(.A(G127gat), .B(G155gat), .Z(new_n227));
  XNOR2_X1  g026(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g027(.A(new_n222), .B(new_n228), .Z(new_n229));
  NAND2_X1  g028(.A1(G85gat), .A2(G92gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n230), .B(KEYINPUT7), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT8), .ZN(new_n232));
  AND2_X1   g031(.A1(G99gat), .A2(G106gat), .ZN(new_n233));
  OAI221_X1 g032(.A(new_n231), .B1(new_n232), .B2(new_n233), .C1(G85gat), .C2(G92gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(G99gat), .A2(G106gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n234), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n237), .B(KEYINPUT109), .ZN(new_n238));
  XNOR2_X1  g037(.A(G43gat), .B(G50gat), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n239), .A2(KEYINPUT15), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(KEYINPUT98), .ZN(new_n242));
  OR3_X1    g041(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(KEYINPUT99), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G29gat), .ZN(new_n245));
  INV_X1    g044(.A(G36gat), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT99), .B1(new_n242), .B2(new_n243), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n240), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n239), .A2(KEYINPUT15), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n240), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n243), .B(KEYINPUT100), .ZN(new_n252));
  INV_X1    g051(.A(new_n242), .ZN(new_n253));
  OAI221_X1 g052(.A(new_n251), .B1(new_n245), .B2(new_n246), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT41), .ZN(new_n257));
  NAND2_X1  g056(.A1(G232gat), .A2(G233gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n255), .A2(KEYINPUT102), .A3(KEYINPUT17), .ZN(new_n259));
  OR2_X1    g058(.A1(KEYINPUT102), .A2(KEYINPUT17), .ZN(new_n260));
  NAND2_X1  g059(.A1(KEYINPUT102), .A2(KEYINPUT17), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n249), .A2(new_n254), .A3(new_n260), .A4(new_n261), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  OAI221_X1 g062(.A(new_n256), .B1(new_n257), .B2(new_n258), .C1(new_n263), .C2(new_n238), .ZN(new_n264));
  XNOR2_X1  g063(.A(G134gat), .B(G162gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  XOR2_X1   g065(.A(G190gat), .B(G218gat), .Z(new_n267));
  NAND2_X1  g066(.A1(new_n258), .A2(new_n257), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  OR2_X1    g069(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n266), .A2(new_n270), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n229), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT35), .ZN(new_n276));
  XNOR2_X1  g075(.A(G78gat), .B(G106gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(KEYINPUT31), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(G50gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT91), .ZN(new_n280));
  XNOR2_X1  g079(.A(G141gat), .B(G148gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(G155gat), .A2(G162gat), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n281), .B1(KEYINPUT2), .B2(new_n282), .ZN(new_n283));
  OR2_X1    g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n284), .A2(KEYINPUT81), .A3(new_n282), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT81), .ZN(new_n286));
  AND2_X1   g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(G155gat), .A2(G162gat), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n283), .A2(new_n290), .ZN(new_n291));
  OR2_X1    g090(.A1(KEYINPUT83), .A2(G155gat), .ZN(new_n292));
  INV_X1    g091(.A(G162gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT84), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT84), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(G162gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(KEYINPUT83), .A2(G155gat), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n292), .A2(new_n294), .A3(new_n296), .A4(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n281), .B1(new_n298), .B2(KEYINPUT2), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT82), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n284), .A2(new_n300), .A3(new_n282), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT82), .B1(new_n287), .B2(new_n288), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT85), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n299), .A2(new_n303), .A3(KEYINPUT85), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n291), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  XOR2_X1   g107(.A(KEYINPUT87), .B(KEYINPUT3), .Z(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT29), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G197gat), .B(G204gat), .ZN(new_n314));
  INV_X1    g113(.A(G211gat), .ZN(new_n315));
  INV_X1    g114(.A(G218gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n314), .B1(KEYINPUT22), .B2(new_n317), .ZN(new_n318));
  XOR2_X1   g117(.A(G211gat), .B(G218gat), .Z(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT74), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n320), .B(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n308), .A2(KEYINPUT29), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n313), .A2(new_n323), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n291), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n299), .A2(KEYINPUT85), .A3(new_n303), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT85), .B1(new_n299), .B2(new_n303), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n309), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(G228gat), .ZN(new_n332));
  INV_X1    g131(.A(G233gat), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G22gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n329), .A2(KEYINPUT3), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n325), .A2(G228gat), .A3(G233gat), .A4(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n334), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n335), .B1(new_n334), .B2(new_n337), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n280), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT91), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n340), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT92), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n344), .A2(new_n345), .A3(new_n338), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n338), .A2(new_n345), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n340), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n341), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n343), .B1(new_n349), .B2(new_n279), .ZN(new_n350));
  NAND2_X1  g149(.A1(G183gat), .A2(G190gat), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT66), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT24), .ZN(new_n354));
  NAND3_X1  g153(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n357));
  OR2_X1    g156(.A1(new_n357), .A2(KEYINPUT67), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT68), .B(G183gat), .ZN(new_n359));
  INV_X1    g158(.A(G190gat), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT67), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n357), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n356), .B(new_n358), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(G169gat), .ZN(new_n364));
  INV_X1    g163(.A(G176gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT23), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT23), .B1(new_n364), .B2(new_n365), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n368), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n363), .A2(KEYINPUT25), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT69), .ZN(new_n372));
  OR2_X1    g171(.A1(new_n368), .A2(KEYINPUT65), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n369), .A2(new_n366), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n351), .A2(new_n354), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n375), .B(new_n357), .C1(G183gat), .C2(G190gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n368), .A2(KEYINPUT65), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n373), .A2(new_n374), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT25), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT69), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n363), .A2(new_n381), .A3(KEYINPUT25), .A4(new_n370), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n372), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n364), .A2(new_n365), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n366), .B(KEYINPUT26), .ZN(new_n385));
  XOR2_X1   g184(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n386));
  INV_X1    g185(.A(G183gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n387), .A2(KEYINPUT27), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n388), .B(KEYINPUT70), .ZN(new_n389));
  AOI21_X1  g188(.A(G190gat), .B1(new_n359), .B2(KEYINPUT27), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n386), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  XOR2_X1   g190(.A(KEYINPUT27), .B(G183gat), .Z(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  AND3_X1   g192(.A1(new_n393), .A2(KEYINPUT28), .A3(new_n360), .ZN(new_n394));
  OAI221_X1 g193(.A(new_n351), .B1(new_n384), .B2(new_n385), .C1(new_n391), .C2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n383), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(G127gat), .B(G134gat), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(KEYINPUT72), .B2(KEYINPUT1), .ZN(new_n398));
  XNOR2_X1  g197(.A(G113gat), .B(G120gat), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n399), .A2(KEYINPUT1), .ZN(new_n400));
  XOR2_X1   g199(.A(new_n398), .B(new_n400), .Z(new_n401));
  XNOR2_X1  g200(.A(new_n396), .B(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(G227gat), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n403), .A2(new_n333), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(KEYINPUT64), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  OR3_X1    g205(.A1(new_n402), .A2(KEYINPUT34), .A3(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT34), .B1(new_n402), .B2(new_n404), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n402), .A2(new_n406), .ZN(new_n411));
  XNOR2_X1  g210(.A(G15gat), .B(G43gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(G71gat), .ZN(new_n413));
  INV_X1    g212(.A(G99gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT33), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n411), .A2(KEYINPUT32), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT73), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n411), .A2(KEYINPUT73), .A3(KEYINPUT32), .A4(new_n416), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT33), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n411), .B1(KEYINPUT32), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n415), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n410), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n421), .A2(new_n424), .A3(new_n410), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n350), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n396), .A2(new_n312), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT77), .ZN(new_n431));
  NAND2_X1  g230(.A1(G226gat), .A2(G233gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(KEYINPUT75), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n430), .A2(new_n431), .A3(new_n434), .ZN(new_n435));
  XOR2_X1   g234(.A(new_n433), .B(KEYINPUT76), .Z(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n396), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT29), .B1(new_n383), .B2(new_n395), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT77), .B1(new_n439), .B2(new_n433), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n435), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n322), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n434), .B1(new_n383), .B2(new_n395), .ZN(new_n443));
  AOI211_X1 g242(.A(new_n322), .B(new_n443), .C1(new_n430), .C2(new_n436), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(G64gat), .B(G92gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n446), .B(G36gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(KEYINPUT78), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n448), .B(new_n205), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n442), .A2(new_n445), .A3(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(KEYINPUT80), .B(KEYINPUT30), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n449), .B1(new_n442), .B2(new_n445), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n442), .A2(new_n445), .ZN(new_n456));
  INV_X1    g255(.A(new_n449), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(KEYINPUT30), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT79), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT79), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n453), .A2(new_n460), .A3(KEYINPUT30), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n455), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT5), .ZN(new_n463));
  INV_X1    g262(.A(new_n401), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n308), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n329), .A2(new_n401), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(G225gat), .A2(G233gat), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n463), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT4), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n308), .A2(KEYINPUT4), .A3(new_n464), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT86), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT3), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n475), .B1(new_n308), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n329), .A2(KEYINPUT86), .A3(KEYINPUT3), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n477), .A2(new_n401), .A3(new_n478), .A4(new_n311), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT88), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n306), .A2(new_n307), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n476), .B1(new_n481), .B2(new_n326), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n464), .B1(new_n482), .B2(KEYINPUT86), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n336), .A2(new_n475), .B1(new_n308), .B2(new_n310), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT88), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  AOI211_X1 g285(.A(new_n469), .B(new_n474), .C1(new_n480), .C2(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n463), .A2(KEYINPUT89), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n470), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n474), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n479), .A2(KEYINPUT88), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n485), .B1(new_n483), .B2(new_n484), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n468), .B(new_n490), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n470), .ZN(new_n494));
  INV_X1    g293(.A(new_n488), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n489), .A2(new_n496), .ZN(new_n497));
  XOR2_X1   g296(.A(G1gat), .B(G29gat), .Z(new_n498));
  XNOR2_X1  g297(.A(KEYINPUT90), .B(KEYINPUT0), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n498), .B(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G57gat), .B(G85gat), .ZN(new_n501));
  XOR2_X1   g300(.A(new_n500), .B(new_n501), .Z(new_n502));
  AOI21_X1  g301(.A(KEYINPUT6), .B1(new_n497), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n503), .B1(new_n497), .B2(new_n502), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n474), .B1(new_n480), .B2(new_n486), .ZN(new_n505));
  AOI211_X1 g304(.A(new_n470), .B(new_n488), .C1(new_n505), .C2(new_n468), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n494), .B1(new_n493), .B2(new_n495), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n502), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n508), .A2(KEYINPUT6), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n462), .B1(new_n504), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n276), .B1(new_n429), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT94), .B1(new_n506), .B2(new_n507), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT94), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n489), .A2(new_n515), .A3(new_n496), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n509), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n503), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT93), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n462), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n460), .B1(new_n453), .B2(KEYINPUT30), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n444), .B1(new_n322), .B2(new_n441), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT30), .ZN(new_n524));
  NOR4_X1   g323(.A1(new_n523), .A2(KEYINPUT79), .A3(new_n524), .A4(new_n449), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n526), .A2(KEYINPUT93), .A3(new_n455), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n510), .A2(new_n519), .B1(new_n521), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n429), .B1(new_n528), .B2(KEYINPUT97), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n502), .B1(new_n514), .B2(new_n516), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT6), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n531), .B1(new_n508), .B2(new_n509), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n510), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT93), .B1(new_n526), .B2(new_n455), .ZN(new_n534));
  AND4_X1   g333(.A1(KEYINPUT93), .A2(new_n455), .A3(new_n459), .A4(new_n461), .ZN(new_n535));
  OAI211_X1 g334(.A(KEYINPUT97), .B(new_n533), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(new_n276), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n513), .B1(new_n529), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n465), .A2(new_n466), .A3(new_n468), .ZN(new_n539));
  OAI211_X1 g338(.A(KEYINPUT39), .B(new_n539), .C1(new_n505), .C2(new_n468), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(new_n469), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n540), .B(new_n502), .C1(KEYINPUT39), .C2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT40), .ZN(new_n544));
  OR3_X1    g343(.A1(new_n505), .A2(KEYINPUT39), .A3(new_n468), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT40), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n545), .A2(new_n546), .A3(new_n502), .A4(new_n540), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n517), .A2(new_n509), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n521), .A2(new_n527), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT95), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n349), .A2(new_n279), .ZN(new_n552));
  INV_X1    g351(.A(new_n343), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OR2_X1    g353(.A1(new_n523), .A2(KEYINPUT37), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n457), .B1(new_n523), .B2(KEYINPUT37), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n453), .B1(new_n557), .B2(KEYINPUT38), .ZN(new_n558));
  AOI211_X1 g357(.A(new_n323), .B(new_n443), .C1(new_n430), .C2(new_n436), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT96), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n441), .A2(new_n323), .ZN(new_n561));
  OAI21_X1  g360(.A(KEYINPUT37), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT38), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n562), .A2(new_n563), .A3(new_n449), .A4(new_n555), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n519), .A2(new_n558), .A3(new_n510), .A4(new_n564), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n521), .A2(new_n527), .A3(new_n548), .A4(KEYINPUT95), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n551), .A2(new_n554), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT36), .ZN(new_n568));
  INV_X1    g367(.A(new_n427), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n568), .B1(new_n569), .B2(new_n425), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n426), .A2(KEYINPUT36), .A3(new_n427), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n511), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n572), .B1(new_n573), .B2(new_n350), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n567), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n275), .B1(new_n538), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT10), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n216), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n238), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n234), .A2(new_n236), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT111), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n236), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n234), .B(new_n583), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n582), .B(new_n215), .C1(new_n584), .C2(new_n581), .ZN(new_n585));
  AND3_X1   g384(.A1(new_n237), .A2(KEYINPUT110), .A3(new_n216), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT110), .B1(new_n237), .B2(new_n216), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n577), .B(new_n585), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n579), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(G230gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n590), .A2(new_n333), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(new_n591), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G120gat), .B(G148gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(new_n365), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n598), .B(G204gat), .Z(new_n599));
  NAND2_X1  g398(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n599), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n593), .A2(new_n595), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n209), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n605), .B1(new_n259), .B2(new_n262), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT103), .ZN(new_n607));
  NAND2_X1  g406(.A1(G229gat), .A2(G233gat), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT103), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n609), .B1(new_n255), .B2(new_n605), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n607), .B(new_n608), .C1(new_n606), .C2(new_n610), .ZN(new_n611));
  OR2_X1    g410(.A1(KEYINPUT104), .A2(KEYINPUT18), .ZN(new_n612));
  NAND2_X1  g411(.A1(KEYINPUT104), .A2(KEYINPUT18), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(KEYINPUT105), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n606), .A2(new_n610), .ZN(new_n616));
  AOI211_X1 g415(.A(new_n609), .B(new_n605), .C1(new_n259), .C2(new_n262), .ZN(new_n617));
  INV_X1    g416(.A(new_n608), .ZN(new_n618));
  NOR3_X1   g417(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n255), .B(new_n605), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n608), .B(KEYINPUT13), .Z(new_n621));
  AOI22_X1  g420(.A1(new_n619), .A2(KEYINPUT18), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT11), .B(G169gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(G197gat), .ZN(new_n624));
  XOR2_X1   g423(.A(G113gat), .B(G141gat), .Z(new_n625));
  XOR2_X1   g424(.A(new_n624), .B(new_n625), .Z(new_n626));
  XOR2_X1   g425(.A(new_n626), .B(KEYINPUT12), .Z(new_n627));
  INV_X1    g426(.A(KEYINPUT105), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n611), .A2(new_n628), .A3(new_n612), .A4(new_n613), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n615), .A2(new_n622), .A3(new_n627), .A4(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n627), .ZN(new_n631));
  INV_X1    g430(.A(new_n614), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n620), .A2(new_n621), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT18), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n633), .B1(new_n611), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n631), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(KEYINPUT106), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT106), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n630), .A2(new_n639), .A3(new_n636), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n576), .A2(new_n604), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n504), .A2(new_n510), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT112), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(new_n203), .ZN(G1324gat));
  NOR2_X1   g447(.A1(new_n534), .A2(new_n535), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n643), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT16), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n652), .A2(new_n205), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n205), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n651), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n651), .A2(KEYINPUT42), .A3(new_n654), .A4(new_n655), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n658), .B(new_n659), .C1(new_n205), .C2(new_n651), .ZN(G1325gat));
  INV_X1    g459(.A(new_n643), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n569), .A2(new_n425), .ZN(new_n662));
  AOI21_X1  g461(.A(G15gat), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(G15gat), .ZN(new_n664));
  INV_X1    g463(.A(new_n572), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n643), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  OR3_X1    g465(.A1(new_n663), .A2(KEYINPUT113), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT113), .B1(new_n663), .B2(new_n666), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(G1326gat));
  NOR2_X1   g468(.A1(new_n643), .A2(new_n554), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT43), .B(G22gat), .Z(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1327gat));
  OAI21_X1  g471(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT97), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n675), .A2(new_n276), .A3(new_n429), .A4(new_n536), .ZN(new_n676));
  AOI22_X1  g475(.A1(new_n676), .A2(new_n513), .B1(new_n567), .B2(new_n574), .ZN(new_n677));
  INV_X1    g476(.A(new_n273), .ZN(new_n678));
  INV_X1    g477(.A(new_n229), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n679), .A2(new_n603), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n642), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n677), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n682), .A2(new_n245), .A3(new_n645), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT45), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n685), .B1(new_n677), .B2(new_n678), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n567), .A2(new_n574), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n536), .A2(new_n276), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n554), .A2(new_n662), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n689), .B1(new_n673), .B2(new_n674), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n512), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  OAI211_X1 g490(.A(KEYINPUT44), .B(new_n273), .C1(new_n687), .C2(new_n691), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n686), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n637), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n679), .A2(new_n694), .A3(new_n603), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n693), .A2(new_n645), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n684), .B1(new_n245), .B2(new_n696), .ZN(G1328gat));
  NAND3_X1  g496(.A1(new_n682), .A2(new_n246), .A3(new_n649), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(KEYINPUT46), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n698), .A2(KEYINPUT46), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n693), .A2(new_n649), .A3(new_n695), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n699), .B(new_n700), .C1(new_n701), .C2(new_n246), .ZN(G1329gat));
  AOI21_X1  g501(.A(new_n678), .B1(new_n538), .B2(new_n575), .ZN(new_n703));
  INV_X1    g502(.A(G43gat), .ZN(new_n704));
  INV_X1    g503(.A(new_n681), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n703), .A2(new_n704), .A3(new_n662), .A4(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT114), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n682), .A2(KEYINPUT114), .A3(new_n704), .A4(new_n662), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n686), .A2(new_n692), .A3(new_n572), .A4(new_n695), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G43gat), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT47), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n710), .A2(KEYINPUT47), .A3(new_n712), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(G1330gat));
  NOR2_X1   g516(.A1(new_n554), .A2(G50gat), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n718), .B(KEYINPUT115), .Z(new_n719));
  AND3_X1   g518(.A1(new_n703), .A2(new_n705), .A3(new_n719), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n686), .A2(new_n692), .A3(new_n350), .A4(new_n695), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n720), .B1(new_n721), .B2(G50gat), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT48), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n722), .A2(KEYINPUT116), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n723), .A2(KEYINPUT116), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n723), .A2(KEYINPUT116), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n722), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n724), .A2(new_n727), .ZN(G1331gat));
  NOR2_X1   g527(.A1(new_n637), .A2(new_n604), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n576), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(new_n646), .ZN(new_n731));
  XOR2_X1   g530(.A(KEYINPUT117), .B(G57gat), .Z(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(G1332gat));
  NOR2_X1   g532(.A1(new_n730), .A2(new_n650), .ZN(new_n734));
  NOR2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  AND2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(new_n734), .B2(new_n735), .ZN(G1333gat));
  INV_X1    g537(.A(KEYINPUT50), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n538), .A2(new_n575), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n740), .A2(new_n662), .A3(new_n274), .A4(new_n729), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT118), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT118), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n576), .A2(new_n743), .A3(new_n662), .A4(new_n729), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(G71gat), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(G71gat), .B1(new_n730), .B2(new_n665), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n739), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(G71gat), .B1(new_n742), .B2(new_n744), .ZN(new_n750));
  INV_X1    g549(.A(new_n748), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n750), .A2(new_n751), .A3(KEYINPUT50), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n749), .A2(new_n752), .ZN(G1334gat));
  NOR2_X1   g552(.A1(new_n730), .A2(new_n554), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n754), .B(G78gat), .Z(G1335gat));
  NAND4_X1  g554(.A1(new_n686), .A2(new_n692), .A3(new_n229), .A4(new_n729), .ZN(new_n756));
  OAI21_X1  g555(.A(G85gat), .B1(new_n756), .B2(new_n646), .ZN(new_n757));
  INV_X1    g556(.A(G85gat), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n679), .A2(new_n637), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT51), .B1(new_n703), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT51), .ZN(new_n761));
  INV_X1    g560(.A(new_n759), .ZN(new_n762));
  NOR4_X1   g561(.A1(new_n677), .A2(new_n761), .A3(new_n678), .A4(new_n762), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n760), .A2(new_n763), .A3(KEYINPUT119), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT119), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n740), .A2(new_n273), .A3(new_n759), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n761), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n703), .A2(KEYINPUT51), .A3(new_n759), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n765), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n758), .B(new_n603), .C1(new_n764), .C2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n757), .B1(new_n770), .B2(new_n646), .ZN(G1336gat));
  OAI21_X1  g570(.A(G92gat), .B1(new_n756), .B2(new_n650), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n650), .A2(G92gat), .A3(new_n604), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT120), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(new_n760), .B2(new_n763), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT52), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n772), .A2(new_n778), .A3(new_n775), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(G1337gat));
  OAI21_X1  g579(.A(G99gat), .B1(new_n756), .B2(new_n665), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n414), .B(new_n603), .C1(new_n764), .C2(new_n769), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n781), .B1(new_n782), .B2(new_n428), .ZN(G1338gat));
  OAI21_X1  g582(.A(G106gat), .B1(new_n756), .B2(new_n554), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n554), .A2(G106gat), .A3(new_n604), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(new_n760), .B2(new_n763), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT121), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n788), .B1(new_n786), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n784), .B(new_n786), .C1(new_n789), .C2(new_n788), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(G1339gat));
  INV_X1    g592(.A(new_n626), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n616), .A2(new_n617), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n795), .A2(new_n608), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n620), .A2(new_n621), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n794), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n630), .A2(new_n603), .A3(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n579), .A2(new_n588), .A3(new_n591), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n593), .A2(KEYINPUT54), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n591), .B1(new_n579), .B2(new_n588), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n601), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n801), .A2(KEYINPUT55), .A3(new_n804), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(new_n602), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT122), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n807), .A2(new_n602), .A3(new_n808), .A4(KEYINPUT122), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n799), .B1(new_n813), .B2(new_n694), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT123), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT123), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n816), .B(new_n799), .C1(new_n813), .C2(new_n694), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(new_n678), .A3(new_n817), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n273), .A2(new_n630), .A3(new_n798), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n819), .A2(new_n811), .A3(new_n812), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n679), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n274), .A2(new_n604), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n822), .A2(new_n637), .ZN(new_n823));
  OR2_X1    g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n646), .A2(new_n649), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n824), .A2(new_n429), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(G113gat), .B1(new_n826), .B2(new_n641), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n826), .A2(G113gat), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n827), .B1(new_n828), .B2(new_n694), .ZN(G1340gat));
  NOR2_X1   g628(.A1(new_n826), .A2(new_n604), .ZN(new_n830));
  XOR2_X1   g629(.A(new_n830), .B(G120gat), .Z(G1341gat));
  NOR2_X1   g630(.A1(new_n826), .A2(new_n229), .ZN(new_n832));
  XOR2_X1   g631(.A(new_n832), .B(G127gat), .Z(G1342gat));
  NOR2_X1   g632(.A1(new_n826), .A2(new_n678), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT56), .ZN(new_n835));
  INV_X1    g634(.A(G134gat), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n837), .B(new_n838), .ZN(G1343gat));
  OAI21_X1  g638(.A(new_n350), .B1(new_n821), .B2(new_n823), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n665), .ZN(new_n841));
  NOR4_X1   g640(.A1(new_n840), .A2(new_n841), .A3(G141gat), .A4(new_n641), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n842), .A2(KEYINPUT58), .ZN(new_n843));
  XOR2_X1   g642(.A(KEYINPUT124), .B(KEYINPUT57), .Z(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n809), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n638), .A2(new_n847), .A3(new_n640), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n799), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n678), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n679), .B1(new_n850), .B2(new_n820), .ZN(new_n851));
  OAI211_X1 g650(.A(KEYINPUT57), .B(new_n350), .C1(new_n851), .C2(new_n823), .ZN(new_n852));
  AOI211_X1 g651(.A(new_n641), .B(new_n841), .C1(new_n846), .C2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(G141gat), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n843), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n841), .B1(new_n846), .B2(new_n852), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n637), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n842), .B1(new_n857), .B2(G141gat), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT58), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n855), .B1(new_n858), .B2(new_n859), .ZN(G1344gat));
  NOR2_X1   g659(.A1(new_n840), .A2(new_n841), .ZN(new_n861));
  INV_X1    g660(.A(G148gat), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n861), .A2(new_n862), .A3(new_n603), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT59), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n822), .A2(new_n642), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n819), .A2(new_n847), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n866), .B1(new_n868), .B2(new_n229), .ZN(new_n869));
  OAI211_X1 g668(.A(KEYINPUT125), .B(new_n865), .C1(new_n869), .C2(new_n554), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT125), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n273), .B1(new_n848), .B2(new_n799), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n819), .A2(new_n847), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n229), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n866), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n554), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n871), .B1(new_n876), .B2(KEYINPUT57), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n350), .B(new_n844), .C1(new_n821), .C2(new_n823), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n870), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n879), .A2(new_n603), .A3(new_n665), .A4(new_n825), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n864), .B1(new_n880), .B2(G148gat), .ZN(new_n881));
  AOI211_X1 g680(.A(KEYINPUT59), .B(new_n862), .C1(new_n856), .C2(new_n603), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n863), .B1(new_n881), .B2(new_n882), .ZN(G1345gat));
  NAND2_X1  g682(.A1(new_n292), .A2(new_n297), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n229), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n861), .A2(new_n679), .ZN(new_n886));
  AOI22_X1  g685(.A1(new_n856), .A2(new_n885), .B1(new_n886), .B2(new_n884), .ZN(G1346gat));
  NAND2_X1  g686(.A1(new_n294), .A2(new_n296), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n678), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n861), .A2(new_n273), .ZN(new_n890));
  AOI22_X1  g689(.A1(new_n856), .A2(new_n889), .B1(new_n890), .B2(new_n888), .ZN(G1347gat));
  NOR2_X1   g690(.A1(new_n645), .A2(new_n650), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n824), .A2(new_n429), .A3(new_n892), .ZN(new_n893));
  OR3_X1    g692(.A1(new_n893), .A2(G169gat), .A3(new_n694), .ZN(new_n894));
  OAI21_X1  g693(.A(G169gat), .B1(new_n893), .B2(new_n641), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1348gat));
  NOR2_X1   g695(.A1(new_n893), .A2(new_n604), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(new_n365), .ZN(G1349gat));
  INV_X1    g697(.A(KEYINPUT60), .ZN(new_n899));
  OAI22_X1  g698(.A1(new_n893), .A2(new_n229), .B1(KEYINPUT126), .B2(new_n359), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT126), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n359), .A2(new_n902), .ZN(new_n903));
  NOR4_X1   g702(.A1(new_n893), .A2(new_n393), .A3(new_n229), .A4(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n899), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n893), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(new_n392), .A3(new_n679), .ZN(new_n907));
  OAI211_X1 g706(.A(KEYINPUT60), .B(new_n900), .C1(new_n907), .C2(new_n903), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n905), .A2(new_n908), .ZN(G1350gat));
  OAI22_X1  g708(.A1(new_n893), .A2(new_n678), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n910));
  NAND2_X1  g709(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n910), .B(new_n911), .ZN(G1351gat));
  NAND2_X1  g711(.A1(new_n892), .A2(new_n665), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n879), .A2(new_n642), .A3(new_n914), .ZN(new_n915));
  XNOR2_X1  g714(.A(KEYINPUT127), .B(G197gat), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n840), .A2(new_n913), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n694), .A2(new_n916), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(G1352gat));
  NOR2_X1   g720(.A1(new_n919), .A2(G204gat), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(new_n603), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(KEYINPUT62), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n879), .A2(new_n603), .A3(new_n914), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(G204gat), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT62), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n922), .A2(new_n927), .A3(new_n603), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n924), .A2(new_n926), .A3(new_n928), .ZN(G1353gat));
  NAND3_X1  g728(.A1(new_n918), .A2(new_n315), .A3(new_n679), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n879), .A2(new_n679), .A3(new_n914), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n931), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n932));
  AOI21_X1  g731(.A(KEYINPUT63), .B1(new_n931), .B2(G211gat), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(G1354gat));
  NAND3_X1  g733(.A1(new_n918), .A2(new_n316), .A3(new_n273), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n879), .A2(new_n273), .A3(new_n914), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n935), .B1(new_n936), .B2(new_n316), .ZN(G1355gat));
endmodule


