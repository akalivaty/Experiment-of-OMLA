//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1 1 0 1 1 0 1 0 1 1 1 1 0 1 0 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n820, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957;
  INV_X1    g000(.A(KEYINPUT30), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT73), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT71), .B(KEYINPUT22), .Z(new_n204));
  INV_X1    g003(.A(G218gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT72), .B(G211gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G197gat), .B(G204gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n209), .B1(new_n207), .B2(new_n208), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n203), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n212), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(KEYINPUT73), .A3(new_n210), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(G226gat), .A2(G233gat), .ZN(new_n217));
  XOR2_X1   g016(.A(new_n217), .B(KEYINPUT74), .Z(new_n218));
  XNOR2_X1  g017(.A(KEYINPUT27), .B(G183gat), .ZN(new_n219));
  INV_X1    g018(.A(G190gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(KEYINPUT28), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n222));
  AOI21_X1  g021(.A(G190gat), .B1(new_n222), .B2(KEYINPUT27), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT27), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n224), .A2(KEYINPUT65), .A3(G183gat), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n221), .B1(new_n226), .B2(KEYINPUT28), .ZN(new_n227));
  INV_X1    g026(.A(G183gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n228), .A2(new_n220), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT66), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT26), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n235), .B1(new_n232), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n234), .B1(new_n233), .B2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n227), .A2(new_n230), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n228), .A2(new_n220), .ZN(new_n240));
  NAND3_X1  g039(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT64), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n240), .B(new_n241), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n244), .B1(new_n243), .B2(new_n242), .ZN(new_n245));
  OR2_X1    g044(.A1(new_n232), .A2(KEYINPUT23), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n232), .A2(KEYINPUT23), .ZN(new_n247));
  NAND2_X1  g046(.A1(G169gat), .A2(G176gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT25), .B1(new_n245), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT25), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n246), .A2(new_n251), .A3(new_n247), .A4(new_n248), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n240), .A2(new_n241), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(new_n242), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n239), .A2(new_n250), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT29), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n218), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  OR2_X1    g058(.A1(new_n233), .A2(new_n237), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n229), .B1(new_n260), .B2(new_n234), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n255), .B1(new_n261), .B2(new_n227), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n217), .B1(new_n262), .B2(new_n250), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n216), .B1(new_n259), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n213), .A2(new_n215), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n257), .A2(new_n218), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT29), .B1(new_n262), .B2(new_n250), .ZN(new_n267));
  INV_X1    g066(.A(new_n217), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n265), .B(new_n266), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n264), .A2(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(G8gat), .B(G36gat), .Z(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT75), .ZN(new_n272));
  XNOR2_X1  g071(.A(G64gat), .B(G92gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n202), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n270), .A2(new_n274), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT40), .ZN(new_n278));
  INV_X1    g077(.A(G148gat), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n279), .A2(G141gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT76), .B(G141gat), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n280), .B1(new_n281), .B2(G148gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G155gat), .ZN(new_n284));
  INV_X1    g083(.A(G162gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT2), .ZN(new_n287));
  NOR2_X1   g086(.A1(G155gat), .A2(G162gat), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n279), .A2(G141gat), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n287), .B1(new_n280), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n286), .A2(new_n288), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n283), .A2(new_n290), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G113gat), .B(G120gat), .ZN(new_n295));
  OAI211_X1 g094(.A(KEYINPUT67), .B(G127gat), .C1(new_n295), .C2(KEYINPUT1), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT1), .ZN(new_n297));
  INV_X1    g096(.A(G127gat), .ZN(new_n298));
  INV_X1    g097(.A(G113gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n299), .A2(G120gat), .ZN(new_n300));
  INV_X1    g099(.A(G120gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(G113gat), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n297), .B(new_n298), .C1(new_n300), .C2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G134gat), .ZN(new_n304));
  AND3_X1   g103(.A1(new_n296), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n304), .B1(new_n296), .B2(new_n303), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n294), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT78), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n296), .A2(new_n303), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G134gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n296), .A2(new_n303), .A3(new_n304), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n313), .A2(KEYINPUT78), .A3(new_n294), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT4), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n292), .A2(new_n293), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n317), .B1(new_n282), .B2(new_n289), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT3), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT3), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n317), .B(new_n320), .C1(new_n282), .C2(new_n289), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n319), .A2(new_n321), .A3(new_n311), .A4(new_n312), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT77), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n305), .A2(new_n306), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT77), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n324), .A2(new_n325), .A3(new_n321), .A4(new_n319), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT4), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n307), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n316), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT39), .ZN(new_n331));
  NAND2_X1  g130(.A1(G225gat), .A2(G233gat), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n330), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  XOR2_X1   g133(.A(KEYINPUT79), .B(KEYINPUT0), .Z(new_n335));
  XNOR2_X1  g134(.A(new_n335), .B(KEYINPUT80), .ZN(new_n336));
  XNOR2_X1  g135(.A(G1gat), .B(G29gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G57gat), .B(G85gat), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n338), .B(new_n339), .Z(new_n340));
  NAND2_X1  g139(.A1(new_n334), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n318), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n309), .A2(new_n314), .A3(new_n332), .A4(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT39), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n344), .B1(new_n330), .B2(new_n333), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n278), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n345), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n347), .A2(KEYINPUT40), .A3(new_n340), .A4(new_n334), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n309), .A2(new_n314), .A3(new_n328), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n313), .A2(KEYINPUT4), .A3(new_n294), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n327), .A2(new_n349), .A3(new_n332), .A4(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT5), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n309), .A2(new_n314), .A3(new_n342), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n352), .B1(new_n353), .B2(new_n333), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n333), .B1(new_n323), .B2(new_n326), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n356), .A2(new_n316), .A3(new_n352), .A4(new_n329), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n340), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n277), .A2(new_n346), .A3(new_n348), .A4(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT6), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n355), .A2(new_n340), .A3(new_n357), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n360), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n358), .A2(KEYINPUT6), .A3(new_n359), .ZN(new_n365));
  INV_X1    g164(.A(new_n276), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n216), .B(new_n266), .C1(new_n267), .C2(new_n268), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n265), .B1(new_n259), .B2(new_n263), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(new_n369), .A3(KEYINPUT37), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT81), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n368), .A2(new_n369), .A3(KEYINPUT81), .A4(KEYINPUT37), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT37), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n264), .A2(new_n269), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT82), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT82), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n264), .A2(new_n269), .A3(new_n378), .A4(new_n375), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n274), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n381), .A2(KEYINPUT38), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n374), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n375), .B1(new_n264), .B2(new_n269), .ZN(new_n384));
  AOI211_X1 g183(.A(new_n381), .B(new_n384), .C1(new_n377), .C2(new_n379), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT38), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n383), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n361), .B1(new_n367), .B2(new_n387), .ZN(new_n388));
  XOR2_X1   g187(.A(G71gat), .B(G99gat), .Z(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(KEYINPUT69), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(G15gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(G43gat), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT68), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n257), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n262), .A2(KEYINPUT68), .A3(new_n250), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n394), .A2(new_n395), .A3(new_n313), .ZN(new_n396));
  INV_X1    g195(.A(G227gat), .ZN(new_n397));
  INV_X1    g196(.A(G233gat), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n262), .A2(new_n324), .A3(KEYINPUT68), .A4(new_n250), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n396), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT33), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n392), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(KEYINPUT32), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n401), .B(KEYINPUT32), .C1(new_n402), .C2(new_n392), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT70), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n396), .A2(new_n400), .ZN(new_n409));
  INV_X1    g208(.A(new_n399), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT34), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT34), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n409), .A2(new_n413), .A3(new_n410), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n407), .A2(new_n408), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n415), .B1(new_n407), .B2(new_n408), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT36), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n415), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n407), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n415), .A2(new_n405), .A3(new_n406), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT36), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT29), .B1(new_n214), .B2(new_n210), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n318), .B1(new_n425), .B2(KEYINPUT3), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n321), .A2(new_n258), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n426), .B1(new_n265), .B2(new_n427), .ZN(new_n428));
  XOR2_X1   g227(.A(G78gat), .B(G106gat), .Z(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(G228gat), .A2(G233gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n431), .B(G22gat), .ZN(new_n432));
  XOR2_X1   g231(.A(KEYINPUT31), .B(G50gat), .Z(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n430), .B(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n388), .A2(new_n418), .A3(new_n424), .A4(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT35), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n364), .A2(new_n365), .ZN(new_n439));
  INV_X1    g238(.A(new_n277), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(new_n440), .A3(new_n436), .ZN(new_n441));
  INV_X1    g240(.A(new_n422), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n438), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n418), .A2(new_n424), .A3(new_n435), .ZN(new_n444));
  NOR3_X1   g243(.A1(new_n416), .A2(new_n417), .A3(new_n435), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT35), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n439), .A2(new_n440), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n437), .B(new_n443), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(G113gat), .B(G141gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n450), .B(G197gat), .ZN(new_n451));
  XOR2_X1   g250(.A(KEYINPUT11), .B(G169gat), .Z(new_n452));
  XNOR2_X1  g251(.A(new_n451), .B(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n453), .B(KEYINPUT12), .ZN(new_n454));
  XNOR2_X1  g253(.A(G15gat), .B(G22gat), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT16), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n455), .B1(new_n456), .B2(G1gat), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n457), .B1(G1gat), .B2(new_n455), .ZN(new_n458));
  XOR2_X1   g257(.A(new_n458), .B(G8gat), .Z(new_n459));
  INV_X1    g258(.A(G29gat), .ZN(new_n460));
  INV_X1    g259(.A(G36gat), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT14), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT14), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n463), .B1(G29gat), .B2(G36gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(G29gat), .A2(G36gat), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(G50gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(G43gat), .ZN(new_n468));
  INV_X1    g267(.A(G43gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(G50gat), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n470), .A3(KEYINPUT15), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT83), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n468), .A2(new_n470), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT15), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n468), .A2(new_n470), .A3(KEYINPUT83), .A4(KEYINPUT15), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n474), .A2(new_n466), .A3(new_n477), .A4(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT84), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT15), .B1(new_n468), .B2(new_n470), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n484), .A2(KEYINPUT84), .A3(new_n474), .A4(new_n478), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n472), .B1(new_n481), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n459), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n472), .ZN(new_n488));
  XNOR2_X1  g287(.A(G43gat), .B(G50gat), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT83), .B1(new_n489), .B2(KEYINPUT15), .ZN(new_n490));
  INV_X1    g289(.A(new_n478), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT84), .B1(new_n492), .B2(new_n484), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n479), .A2(new_n480), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n488), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT17), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT17), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n486), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n487), .B1(new_n499), .B2(new_n459), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT85), .ZN(new_n501));
  NAND2_X1  g300(.A1(G229gat), .A2(G233gat), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT18), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n481), .A2(new_n485), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n497), .B1(new_n504), .B2(new_n488), .ZN(new_n505));
  AOI211_X1 g304(.A(KEYINPUT17), .B(new_n472), .C1(new_n481), .C2(new_n485), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n459), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n459), .A2(new_n486), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n507), .A2(KEYINPUT18), .A3(new_n502), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT85), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n503), .A2(new_n510), .ZN(new_n511));
  XOR2_X1   g310(.A(new_n502), .B(KEYINPUT13), .Z(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n459), .A2(new_n486), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n513), .B1(new_n508), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n507), .A2(new_n502), .A3(new_n508), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT18), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n454), .B1(new_n511), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n509), .A2(KEYINPUT85), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n509), .A2(KEYINPUT85), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n454), .B(new_n518), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n449), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT21), .ZN(new_n526));
  AND2_X1   g325(.A1(G71gat), .A2(G78gat), .ZN(new_n527));
  NOR2_X1   g326(.A1(G71gat), .A2(G78gat), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n527), .B1(KEYINPUT9), .B2(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(KEYINPUT86), .B(G57gat), .Z(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(G64gat), .ZN(new_n531));
  INV_X1    g330(.A(G64gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(G57gat), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n529), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  XOR2_X1   g333(.A(G57gat), .B(G64gat), .Z(new_n535));
  AOI211_X1 g334(.A(new_n527), .B(new_n528), .C1(new_n535), .C2(KEYINPUT9), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n459), .B1(new_n526), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(KEYINPUT90), .ZN(new_n540));
  XNOR2_X1  g339(.A(G127gat), .B(G155gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(G231gat), .A2(G233gat), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(KEYINPUT87), .B(KEYINPUT21), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n537), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n543), .B1(new_n537), .B2(new_n544), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n548), .B1(new_n546), .B2(new_n547), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n541), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n551), .ZN(new_n553));
  INV_X1    g352(.A(new_n541), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(new_n554), .A3(new_n549), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n540), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G183gat), .B(G211gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT89), .B(KEYINPUT20), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n552), .A2(new_n555), .A3(new_n540), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n557), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n560), .ZN(new_n563));
  INV_X1    g362(.A(new_n561), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n563), .B1(new_n564), .B2(new_n556), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G134gat), .B(G162gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(G232gat), .A2(G233gat), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT41), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n567), .B(new_n570), .Z(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT91), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT7), .ZN(new_n574));
  NAND2_X1  g373(.A1(G85gat), .A2(G92gat), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n574), .B(new_n575), .Z(new_n576));
  NOR2_X1   g375(.A1(G85gat), .A2(G92gat), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT8), .ZN(new_n578));
  NAND2_X1  g377(.A1(G99gat), .A2(G106gat), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT92), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(KEYINPUT92), .A2(G99gat), .A3(G106gat), .ZN(new_n582));
  AOI211_X1 g381(.A(KEYINPUT93), .B(new_n577), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT93), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n579), .A2(new_n580), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n585), .A2(KEYINPUT8), .A3(new_n582), .ZN(new_n586));
  INV_X1    g385(.A(new_n577), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n584), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n576), .B1(new_n583), .B2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G99gat), .B(G106gat), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n590), .B(new_n576), .C1(new_n583), .C2(new_n588), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI22_X1  g393(.A1(new_n594), .A2(new_n486), .B1(new_n569), .B2(new_n568), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT95), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n594), .B1(new_n505), .B2(new_n506), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT94), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT94), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n600), .B(new_n594), .C1(new_n505), .C2(new_n506), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(G190gat), .B(G218gat), .Z(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n597), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n604), .B1(new_n597), .B2(new_n602), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n572), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n597), .A2(new_n602), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(new_n603), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n597), .A2(new_n602), .A3(new_n604), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n609), .A2(new_n571), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G230gat), .A2(G233gat), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n586), .A2(new_n587), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT93), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n586), .A2(new_n584), .A3(new_n587), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n590), .B1(new_n618), .B2(new_n576), .ZN(new_n619));
  INV_X1    g418(.A(new_n593), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n538), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT10), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n592), .A2(new_n537), .A3(new_n593), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n592), .A2(KEYINPUT10), .A3(new_n537), .A4(new_n593), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n614), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n613), .B1(new_n621), .B2(new_n623), .ZN(new_n627));
  XNOR2_X1  g426(.A(G120gat), .B(G148gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(G176gat), .B(G204gat), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n628), .B(new_n629), .Z(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n626), .A2(new_n627), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n631), .B1(new_n626), .B2(new_n627), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n566), .A2(new_n612), .A3(new_n636), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n525), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n439), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g441(.A(KEYINPUT16), .B(G8gat), .Z(new_n643));
  NAND3_X1  g442(.A1(new_n639), .A2(new_n277), .A3(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(G8gat), .B1(new_n638), .B2(new_n440), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  MUX2_X1   g445(.A(new_n644), .B(new_n646), .S(KEYINPUT42), .Z(G1325gat));
  OR3_X1    g446(.A1(new_n638), .A2(G15gat), .A3(new_n442), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n418), .A2(new_n424), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(G15gat), .B1(new_n638), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT96), .ZN(G1326gat));
  NOR2_X1   g452(.A1(new_n638), .A2(new_n436), .ZN(new_n654));
  XOR2_X1   g453(.A(KEYINPUT43), .B(G22gat), .Z(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(G1327gat));
  AND2_X1   g455(.A1(new_n607), .A2(new_n611), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n437), .A2(new_n443), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n448), .B1(new_n444), .B2(new_n446), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT44), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI211_X1 g461(.A(KEYINPUT44), .B(new_n657), .C1(new_n658), .C2(new_n659), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n635), .B(KEYINPUT98), .Z(new_n664));
  INV_X1    g463(.A(new_n524), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n664), .A2(new_n665), .A3(new_n566), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n662), .A2(new_n663), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(KEYINPUT99), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT99), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n662), .A2(new_n669), .A3(new_n663), .A4(new_n666), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n668), .A2(new_n640), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(G29gat), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n566), .A2(new_n612), .A3(new_n635), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n524), .B(new_n673), .C1(new_n658), .C2(new_n659), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT97), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n439), .A2(G29gat), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n677), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT97), .B1(new_n674), .B2(new_n679), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n678), .A2(KEYINPUT45), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(KEYINPUT45), .B1(new_n678), .B2(new_n680), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n672), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT100), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n672), .A2(new_n683), .A3(KEYINPUT100), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(G1328gat));
  NAND3_X1  g487(.A1(new_n668), .A2(new_n277), .A3(new_n670), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n461), .B1(new_n689), .B2(KEYINPUT101), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(KEYINPUT101), .B2(new_n689), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n674), .A2(G36gat), .A3(new_n440), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT46), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(G1329gat));
  OAI21_X1  g493(.A(G43gat), .B1(new_n667), .B2(new_n650), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n674), .A2(G43gat), .A3(new_n442), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n695), .A2(KEYINPUT47), .A3(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n668), .A2(new_n649), .A3(new_n670), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n696), .B1(new_n699), .B2(G43gat), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n700), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g500(.A1(new_n674), .A2(G50gat), .A3(new_n436), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT48), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n705), .B1(new_n667), .B2(new_n436), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(G50gat), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n667), .A2(new_n705), .A3(new_n436), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n704), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n668), .A2(new_n435), .A3(new_n670), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n702), .B1(new_n710), .B2(G50gat), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n709), .B1(new_n711), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g511(.A(new_n664), .ZN(new_n713));
  INV_X1    g512(.A(new_n566), .ZN(new_n714));
  NOR4_X1   g513(.A1(new_n713), .A2(new_n714), .A3(new_n524), .A4(new_n657), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n449), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n640), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(new_n530), .Z(G1332gat));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n277), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n720));
  XOR2_X1   g519(.A(KEYINPUT49), .B(G64gat), .Z(new_n721));
  OAI21_X1  g520(.A(new_n720), .B1(new_n719), .B2(new_n721), .ZN(G1333gat));
  NAND3_X1  g521(.A1(new_n716), .A2(G71gat), .A3(new_n649), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT103), .ZN(new_n724));
  INV_X1    g523(.A(G71gat), .ZN(new_n725));
  INV_X1    g524(.A(new_n716), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n422), .B(KEYINPUT104), .Z(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT50), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT50), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n724), .A2(new_n731), .A3(new_n728), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(G1334gat));
  NAND2_X1  g532(.A1(new_n716), .A2(new_n435), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g534(.A1(new_n524), .A2(new_n566), .A3(new_n636), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n662), .A2(new_n663), .A3(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n662), .A2(KEYINPUT105), .A3(new_n663), .A4(new_n736), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n739), .A2(new_n640), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G85gat), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n449), .A2(new_n665), .A3(new_n714), .A4(new_n657), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n439), .A2(G85gat), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n745), .A2(new_n635), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n742), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT106), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n742), .A2(new_n747), .A3(KEYINPUT106), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(G1336gat));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753));
  OAI21_X1  g552(.A(G92gat), .B1(new_n737), .B2(new_n440), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n743), .B(KEYINPUT51), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n713), .A2(G92gat), .A3(new_n440), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n753), .B(new_n754), .C1(new_n755), .C2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n744), .A2(KEYINPUT107), .ZN(new_n759));
  XOR2_X1   g558(.A(new_n743), .B(new_n759), .Z(new_n760));
  NAND3_X1  g559(.A1(new_n739), .A2(new_n277), .A3(new_n740), .ZN(new_n761));
  AOI22_X1  g560(.A1(new_n760), .A2(new_n756), .B1(new_n761), .B2(G92gat), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n758), .B1(new_n762), .B2(new_n753), .ZN(G1337gat));
  OR4_X1    g562(.A1(G99gat), .A2(new_n755), .A3(new_n442), .A4(new_n636), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n739), .A2(new_n649), .A3(new_n740), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G99gat), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(G1338gat));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n768));
  OAI21_X1  g567(.A(G106gat), .B1(new_n737), .B2(new_n436), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n713), .A2(G106gat), .A3(new_n436), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n768), .B(new_n769), .C1(new_n755), .C2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n739), .A2(new_n435), .A3(new_n740), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n760), .A2(new_n770), .B1(new_n773), .B2(G106gat), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n772), .B1(new_n774), .B2(new_n768), .ZN(G1339gat));
  INV_X1    g574(.A(KEYINPUT54), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n777));
  INV_X1    g576(.A(new_n625), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n776), .B(new_n613), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n625), .A2(new_n614), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT54), .B1(new_n777), .B2(new_n780), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n779), .B(new_n631), .C1(new_n781), .C2(new_n626), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n613), .B1(new_n777), .B2(new_n778), .ZN(new_n785));
  INV_X1    g584(.A(new_n780), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n776), .B1(new_n786), .B2(new_n624), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n783), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n630), .B1(new_n626), .B2(new_n776), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n632), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n523), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n784), .B(new_n790), .C1(new_n791), .C2(new_n519), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n508), .A2(new_n514), .A3(new_n513), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT108), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n500), .A2(new_n502), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n453), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n796), .A2(new_n523), .A3(new_n635), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n657), .B1(new_n792), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n790), .A2(new_n784), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n796), .A2(new_n523), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n612), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n714), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  OR2_X1    g601(.A1(new_n637), .A2(new_n524), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n439), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n804), .A2(new_n440), .A3(new_n445), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(KEYINPUT109), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n524), .A2(new_n299), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT110), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n435), .B1(new_n802), .B2(new_n803), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n439), .A2(new_n277), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n810), .A2(new_n422), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(G113gat), .B1(new_n812), .B2(new_n665), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n809), .A2(new_n813), .ZN(G1340gat));
  NAND2_X1  g613(.A1(new_n635), .A2(new_n301), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT111), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n806), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(G120gat), .B1(new_n812), .B2(new_n713), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(G1341gat));
  NAND3_X1  g618(.A1(new_n805), .A2(new_n298), .A3(new_n566), .ZN(new_n820));
  OAI21_X1  g619(.A(G127gat), .B1(new_n812), .B2(new_n714), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(G1342gat));
  XOR2_X1   g621(.A(KEYINPUT67), .B(G134gat), .Z(new_n823));
  NAND3_X1  g622(.A1(new_n805), .A2(new_n657), .A3(new_n823), .ZN(new_n824));
  XOR2_X1   g623(.A(new_n824), .B(KEYINPUT56), .Z(new_n825));
  OAI21_X1  g624(.A(G134gat), .B1(new_n812), .B2(new_n612), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(G1343gat));
  INV_X1    g626(.A(new_n281), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n650), .A2(new_n811), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n802), .A2(new_n803), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n831), .A2(KEYINPUT113), .A3(KEYINPUT57), .A4(new_n435), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n436), .B1(new_n802), .B2(new_n803), .ZN(new_n833));
  XNOR2_X1  g632(.A(KEYINPUT112), .B(KEYINPUT57), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n832), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n837));
  AOI211_X1 g636(.A(new_n837), .B(new_n436), .C1(new_n802), .C2(new_n803), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(KEYINPUT113), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n830), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n828), .B1(new_n840), .B2(new_n665), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n444), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n804), .A2(new_n843), .ZN(new_n844));
  NOR4_X1   g643(.A1(new_n844), .A2(G141gat), .A3(new_n665), .A4(new_n277), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT58), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT114), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT114), .B1(new_n804), .B2(new_n843), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n848), .A2(new_n277), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n665), .A2(G141gat), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT58), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n852), .A2(new_n841), .A3(KEYINPUT115), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT115), .B1(new_n852), .B2(new_n841), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n846), .B1(new_n853), .B2(new_n854), .ZN(G1344gat));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n799), .B1(new_n520), .B2(new_n523), .ZN(new_n858));
  INV_X1    g657(.A(new_n797), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n612), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n801), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n566), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n637), .A2(new_n524), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n435), .B(new_n835), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n864), .B1(KEYINPUT57), .B2(new_n833), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT116), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n811), .A2(new_n418), .A3(new_n866), .A4(new_n424), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n635), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n868), .B1(KEYINPUT116), .B2(new_n829), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n279), .B1(new_n865), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT59), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n857), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n869), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n831), .A2(new_n435), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n837), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n873), .B1(new_n875), .B2(new_n864), .ZN(new_n876));
  OAI211_X1 g675(.A(KEYINPUT117), .B(KEYINPUT59), .C1(new_n876), .C2(new_n279), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n635), .B(new_n830), .C1(new_n836), .C2(new_n839), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n279), .A2(KEYINPUT59), .ZN(new_n879));
  AOI22_X1  g678(.A1(new_n872), .A2(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n850), .A2(new_n279), .A3(new_n635), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n856), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n878), .A2(new_n879), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT57), .B1(new_n831), .B2(new_n435), .ZN(new_n885));
  AOI211_X1 g684(.A(new_n436), .B(new_n834), .C1(new_n802), .C2(new_n803), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n869), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(G148gat), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT117), .B1(new_n888), .B2(KEYINPUT59), .ZN(new_n889));
  AOI211_X1 g688(.A(new_n857), .B(new_n871), .C1(new_n887), .C2(G148gat), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n884), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(KEYINPUT118), .A3(new_n881), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n883), .A2(new_n892), .ZN(G1345gat));
  OAI21_X1  g692(.A(G155gat), .B1(new_n840), .B2(new_n714), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n850), .A2(new_n284), .A3(new_n566), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1346gat));
  NOR3_X1   g695(.A1(new_n840), .A2(new_n285), .A3(new_n612), .ZN(new_n897));
  AOI21_X1  g696(.A(G162gat), .B1(new_n850), .B2(new_n657), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n897), .A2(new_n898), .ZN(G1347gat));
  NOR2_X1   g698(.A1(new_n640), .A2(new_n440), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n831), .A2(new_n900), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n901), .A2(new_n445), .ZN(new_n902));
  AOI21_X1  g701(.A(G169gat), .B1(new_n902), .B2(new_n524), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n900), .B(KEYINPUT119), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n904), .A2(new_n727), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n905), .A2(new_n810), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n524), .A2(G169gat), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(G1348gat));
  NAND3_X1  g707(.A1(new_n906), .A2(G176gat), .A3(new_n664), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT120), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n909), .A2(new_n910), .ZN(new_n912));
  AOI21_X1  g711(.A(G176gat), .B1(new_n902), .B2(new_n635), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(G1349gat));
  AOI21_X1  g713(.A(new_n228), .B1(new_n906), .B2(new_n566), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n566), .A2(new_n219), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n902), .B2(new_n916), .ZN(new_n917));
  XOR2_X1   g716(.A(new_n917), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g717(.A(new_n220), .B1(new_n906), .B2(new_n657), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT61), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OR2_X1    g720(.A1(new_n921), .A2(KEYINPUT122), .ZN(new_n922));
  OR3_X1    g721(.A1(new_n919), .A2(KEYINPUT121), .A3(new_n920), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT121), .B1(new_n919), .B2(new_n920), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n921), .A2(KEYINPUT122), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n922), .A2(new_n923), .A3(new_n924), .A4(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n902), .A2(new_n220), .A3(new_n657), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1351gat));
  AND2_X1   g727(.A1(new_n901), .A2(new_n843), .ZN(new_n929));
  XOR2_X1   g728(.A(KEYINPUT123), .B(G197gat), .Z(new_n930));
  NAND3_X1  g729(.A1(new_n929), .A2(new_n524), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n904), .A2(new_n649), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT124), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(new_n865), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n934), .A2(new_n665), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n931), .B1(new_n935), .B2(new_n930), .ZN(G1352gat));
  INV_X1    g735(.A(G204gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n929), .A2(new_n937), .A3(new_n635), .ZN(new_n938));
  XOR2_X1   g737(.A(new_n938), .B(KEYINPUT62), .Z(new_n939));
  NOR3_X1   g738(.A1(new_n934), .A2(KEYINPUT125), .A3(new_n713), .ZN(new_n940));
  OAI21_X1  g739(.A(KEYINPUT125), .B1(new_n934), .B2(new_n713), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G204gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n939), .B1(new_n940), .B2(new_n942), .ZN(G1353gat));
  NAND3_X1  g742(.A1(new_n933), .A2(new_n566), .A3(new_n865), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(G211gat), .B1(new_n944), .B2(new_n945), .ZN(new_n948));
  OAI21_X1  g747(.A(KEYINPUT63), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n944), .A2(new_n945), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT63), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n950), .A2(new_n951), .A3(G211gat), .A4(new_n946), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n929), .A2(new_n206), .A3(new_n566), .ZN(new_n953));
  XOR2_X1   g752(.A(new_n953), .B(KEYINPUT126), .Z(new_n954));
  NAND3_X1  g753(.A1(new_n949), .A2(new_n952), .A3(new_n954), .ZN(G1354gat));
  OAI21_X1  g754(.A(G218gat), .B1(new_n934), .B2(new_n612), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n929), .A2(new_n205), .A3(new_n657), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(G1355gat));
endmodule


