//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 0 0 1 1 1 1 0 1 1 0 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  INV_X1    g001(.A(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  INV_X1    g007(.A(G218gat), .ZN(new_n209));
  INV_X1    g008(.A(G211gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT72), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT72), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G211gat), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n209), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n207), .B(new_n208), .C1(new_n214), .C2(KEYINPUT22), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT22), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT72), .B(G211gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n217), .B1(new_n218), .B2(new_n209), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n208), .B1(new_n219), .B2(new_n207), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n216), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(G141gat), .B(G148gat), .Z(new_n222));
  NAND2_X1  g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT2), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(new_n223), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT76), .ZN(new_n228));
  NAND3_X1  g027(.A1(KEYINPUT75), .A2(G155gat), .A3(G162gat), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n228), .B1(new_n227), .B2(new_n229), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n225), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT2), .ZN(new_n233));
  INV_X1    g032(.A(G155gat), .ZN(new_n234));
  INV_X1    g033(.A(G162gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n222), .A2(new_n233), .A3(new_n223), .A4(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT3), .B1(new_n232), .B2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n221), .B1(new_n238), .B2(KEYINPUT29), .ZN(new_n239));
  INV_X1    g038(.A(new_n237), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n227), .A2(new_n229), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT76), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n240), .B1(new_n244), .B2(new_n225), .ZN(new_n245));
  INV_X1    g044(.A(new_n208), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n211), .A2(new_n213), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT22), .B1(new_n247), .B2(G218gat), .ZN(new_n248));
  INV_X1    g047(.A(new_n207), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n246), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT29), .B1(new_n250), .B2(new_n215), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n245), .B1(new_n251), .B2(KEYINPUT3), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n239), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G228gat), .ZN(new_n254));
  INV_X1    g053(.A(G233gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT29), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n259), .B1(new_n216), .B2(new_n220), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT3), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT81), .B1(new_n262), .B2(new_n245), .ZN(new_n263));
  OAI211_X1 g062(.A(KEYINPUT81), .B(new_n245), .C1(new_n251), .C2(KEYINPUT3), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n256), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n239), .A2(KEYINPUT82), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT82), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n221), .B(new_n268), .C1(new_n238), .C2(KEYINPUT29), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n258), .B1(new_n266), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(G22gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n271), .A2(G22gat), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n206), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT83), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n271), .A2(new_n277), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n258), .B(KEYINPUT83), .C1(new_n266), .C2(new_n270), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n278), .A2(KEYINPUT84), .A3(G22gat), .A4(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n206), .B1(new_n272), .B2(new_n273), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n273), .B1(new_n271), .B2(new_n277), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT84), .B1(new_n283), .B2(new_n279), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n276), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n245), .A2(KEYINPUT3), .ZN(new_n286));
  XOR2_X1   g085(.A(G127gat), .B(G134gat), .Z(new_n287));
  XNOR2_X1  g086(.A(G113gat), .B(G120gat), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n287), .B1(KEYINPUT1), .B2(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(G113gat), .B(G120gat), .Z(new_n290));
  INV_X1    g089(.A(KEYINPUT1), .ZN(new_n291));
  XNOR2_X1  g090(.A(G127gat), .B(G134gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT77), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n289), .A2(new_n293), .A3(KEYINPUT77), .ZN(new_n297));
  AND2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n232), .A2(new_n237), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(new_n261), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n286), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT5), .ZN(new_n302));
  NAND2_X1  g101(.A1(G225gat), .A2(G233gat), .ZN(new_n303));
  AND3_X1   g102(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n294), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n299), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT4), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT79), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n306), .A2(KEYINPUT79), .A3(KEYINPUT4), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT67), .B1(new_n289), .B2(new_n293), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n289), .A2(new_n293), .A3(KEYINPUT67), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT4), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n314), .A2(new_n315), .A3(new_n299), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n309), .A2(new_n310), .A3(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n314), .A2(KEYINPUT4), .A3(new_n299), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n306), .A2(new_n315), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n301), .A2(new_n303), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n296), .A2(new_n297), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n306), .B1(new_n321), .B2(new_n299), .ZN(new_n322));
  INV_X1    g121(.A(new_n303), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n302), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n304), .A2(new_n317), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT6), .ZN(new_n326));
  XOR2_X1   g125(.A(G1gat), .B(G29gat), .Z(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G57gat), .B(G85gat), .ZN(new_n330));
  XOR2_X1   g129(.A(new_n329), .B(new_n330), .Z(new_n331));
  NOR3_X1   g130(.A1(new_n325), .A2(new_n326), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n304), .A2(new_n317), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n320), .A2(new_n324), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n331), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT6), .B1(new_n325), .B2(new_n331), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n332), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  XOR2_X1   g138(.A(G8gat), .B(G36gat), .Z(new_n340));
  XNOR2_X1  g139(.A(G64gat), .B(G92gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(G226gat), .A2(G233gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n343), .B(KEYINPUT73), .ZN(new_n344));
  NAND3_X1  g143(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G183gat), .ZN(new_n348));
  INV_X1    g147(.A(G190gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n345), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT64), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT25), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G169gat), .ZN(new_n354));
  INV_X1    g153(.A(G176gat), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT23), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(G169gat), .A2(G176gat), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n357), .A2(KEYINPUT23), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n351), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n353), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n360), .B1(new_n358), .B2(new_n356), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n364), .B(new_n351), .C1(new_n352), .C2(KEYINPUT25), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n354), .A2(new_n355), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT26), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n367), .B1(new_n368), .B2(new_n357), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n358), .A2(KEYINPUT26), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n350), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n348), .A2(KEYINPUT27), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT27), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(G183gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT66), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT66), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n372), .A2(new_n374), .A3(new_n377), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n349), .A2(KEYINPUT28), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT65), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(G190gat), .B1(new_n372), .B2(KEYINPUT65), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT28), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n371), .B1(new_n380), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n366), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n344), .B1(new_n386), .B2(new_n259), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n343), .B1(new_n366), .B2(new_n385), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n221), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n386), .A2(new_n344), .ZN(new_n390));
  INV_X1    g189(.A(new_n221), .ZN(new_n391));
  INV_X1    g190(.A(new_n343), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT29), .B1(new_n366), .B2(new_n385), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n390), .B(new_n391), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n342), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT30), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n389), .A2(new_n394), .A3(new_n342), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n389), .A2(KEYINPUT30), .A3(new_n394), .A4(new_n342), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n399), .A2(KEYINPUT74), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n399), .A2(KEYINPUT74), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n398), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n339), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n314), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n289), .A2(new_n293), .A3(KEYINPUT67), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n405), .A2(new_n311), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n406), .A2(new_n366), .A3(new_n385), .ZN(new_n407));
  INV_X1    g206(.A(G227gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n408), .A2(new_n255), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n404), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  XOR2_X1   g209(.A(G71gat), .B(G99gat), .Z(new_n411));
  XNOR2_X1  g210(.A(G15gat), .B(G43gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT33), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT68), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n410), .A2(KEYINPUT32), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n404), .A2(new_n407), .A3(new_n409), .A4(new_n413), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n414), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT68), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n410), .A2(KEYINPUT32), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n418), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT70), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n404), .A2(new_n407), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n409), .A2(KEYINPUT34), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n426), .ZN(new_n428));
  AOI211_X1 g227(.A(KEYINPUT70), .B(new_n428), .C1(new_n404), .C2(new_n407), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n406), .A2(new_n366), .A3(new_n385), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n366), .A2(new_n385), .B1(new_n312), .B2(new_n313), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT69), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT69), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n404), .A2(new_n434), .A3(new_n407), .ZN(new_n435));
  INV_X1    g234(.A(new_n409), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n433), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT34), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n430), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n415), .B1(new_n419), .B2(new_n414), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n410), .A2(KEYINPUT32), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n417), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n443), .A2(new_n438), .A3(new_n430), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT71), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n440), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n423), .A2(new_n439), .A3(KEYINPUT71), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n285), .A2(new_n403), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT35), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT88), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT88), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n449), .A2(new_n452), .A3(KEYINPUT35), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n335), .A2(KEYINPUT6), .A3(new_n336), .ZN(new_n455));
  OR2_X1    g254(.A1(new_n455), .A2(KEYINPUT87), .ZN(new_n456));
  XOR2_X1   g255(.A(new_n331), .B(KEYINPUT85), .Z(new_n457));
  OAI21_X1  g256(.A(new_n338), .B1(new_n325), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n455), .A2(KEYINPUT87), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n456), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n440), .A2(new_n444), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  OR2_X1    g261(.A1(new_n402), .A2(KEYINPUT35), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n285), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n454), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n395), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT37), .ZN(new_n468));
  OR2_X1    g267(.A1(new_n342), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n468), .B1(new_n389), .B2(new_n394), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT38), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n393), .A2(new_n392), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n474), .B1(new_n344), .B2(new_n386), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n468), .B1(new_n475), .B2(new_n221), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n391), .B1(new_n387), .B2(new_n388), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT38), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n470), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n460), .A2(new_n397), .A3(new_n473), .A4(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n303), .B1(new_n317), .B2(new_n301), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT39), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT39), .B1(new_n322), .B2(new_n323), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n483), .B(new_n457), .C1(new_n481), .C2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT40), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  XOR2_X1   g286(.A(new_n487), .B(KEYINPUT86), .Z(new_n488));
  OAI221_X1 g287(.A(new_n402), .B1(new_n325), .B2(new_n457), .C1(new_n486), .C2(new_n485), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n480), .B(new_n285), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n448), .A2(KEYINPUT36), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n461), .A2(KEYINPUT36), .ZN(new_n492));
  OR2_X1    g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OR2_X1    g292(.A1(new_n285), .A2(new_n403), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n490), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n466), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G43gat), .B(G50gat), .ZN(new_n497));
  OR2_X1    g296(.A1(new_n497), .A2(KEYINPUT15), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(KEYINPUT15), .ZN(new_n499));
  NAND2_X1  g298(.A1(G29gat), .A2(G36gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NOR3_X1   g301(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n503), .B(KEYINPUT91), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT92), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n505), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n503), .A2(KEYINPUT91), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n503), .A2(KEYINPUT91), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n512), .A2(KEYINPUT92), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n502), .B1(new_n508), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n503), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n505), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT90), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n516), .A2(new_n517), .B1(G29gat), .B2(G36gat), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n515), .A2(KEYINPUT90), .A3(new_n505), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n499), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n514), .A2(KEYINPUT17), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT17), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n507), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n512), .A2(KEYINPUT92), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n501), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n523), .B1(new_n526), .B2(new_n520), .ZN(new_n527));
  XNOR2_X1  g326(.A(G15gat), .B(G22gat), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT93), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(G8gat), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT16), .ZN(new_n532));
  AOI21_X1  g331(.A(G1gat), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n531), .B(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n522), .A2(new_n527), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n514), .A2(new_n521), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n531), .B(new_n533), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G229gat), .A2(G233gat), .ZN(new_n541));
  XOR2_X1   g340(.A(new_n541), .B(KEYINPUT94), .Z(new_n542));
  NOR2_X1   g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n543), .A2(KEYINPUT18), .ZN(new_n544));
  XOR2_X1   g343(.A(KEYINPUT95), .B(KEYINPUT13), .Z(new_n545));
  XNOR2_X1  g344(.A(new_n542), .B(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n537), .A2(KEYINPUT96), .A3(new_n538), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n535), .A2(new_n521), .A3(new_n514), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT96), .B1(new_n537), .B2(new_n538), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n547), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n542), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n536), .A2(KEYINPUT18), .A3(new_n553), .A4(new_n539), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G113gat), .B(G141gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(G197gat), .ZN(new_n557));
  XOR2_X1   g356(.A(KEYINPUT11), .B(G169gat), .Z(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT12), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NOR3_X1   g360(.A1(new_n544), .A2(new_n555), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT97), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n555), .A2(new_n563), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n543), .A2(KEYINPUT18), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n552), .A2(KEYINPUT97), .A3(new_n554), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n560), .B(KEYINPUT89), .Z(new_n568));
  AOI21_X1  g367(.A(new_n562), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(G85gat), .A2(G92gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT7), .ZN(new_n572));
  NAND2_X1  g371(.A1(G99gat), .A2(G106gat), .ZN(new_n573));
  INV_X1    g372(.A(G85gat), .ZN(new_n574));
  INV_X1    g373(.A(G92gat), .ZN(new_n575));
  AOI22_X1  g374(.A1(KEYINPUT8), .A2(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT100), .ZN(new_n577));
  XNOR2_X1  g376(.A(G99gat), .B(G106gat), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n572), .B(new_n576), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n577), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n522), .A2(new_n527), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n581), .ZN(new_n583));
  AND2_X1   g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584));
  AOI22_X1  g383(.A1(new_n537), .A2(new_n583), .B1(KEYINPUT41), .B2(new_n584), .ZN(new_n585));
  AND3_X1   g384(.A1(new_n582), .A2(new_n585), .A3(new_n349), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n349), .B1(new_n582), .B2(new_n585), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n209), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n582), .A2(new_n585), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(G190gat), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n582), .A2(new_n585), .A3(new_n349), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n590), .A2(G218gat), .A3(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT99), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n588), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n584), .A2(KEYINPUT41), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n595), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n588), .A2(new_n592), .A3(new_n593), .A4(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(G134gat), .B(G162gat), .Z(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(G57gat), .B(G64gat), .Z(new_n603));
  NAND2_X1  g402(.A1(G71gat), .A2(G78gat), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT9), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(G71gat), .A2(G78gat), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  AOI22_X1  g408(.A1(new_n604), .A2(new_n609), .B1(new_n606), .B2(KEYINPUT98), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n607), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n613), .A2(KEYINPUT21), .ZN(new_n614));
  NAND2_X1  g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(G127gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n538), .B1(KEYINPUT21), .B2(new_n613), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(G155gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(G183gat), .B(G211gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n620), .B(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n596), .A2(new_n600), .A3(new_n598), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n602), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT101), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n602), .A2(new_n625), .A3(KEYINPUT101), .A4(new_n626), .ZN(new_n630));
  XOR2_X1   g429(.A(G120gat), .B(G148gat), .Z(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT102), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n632), .B(KEYINPUT103), .Z(new_n633));
  XNOR2_X1  g432(.A(G176gat), .B(G204gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n613), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n581), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT10), .ZN(new_n639));
  AND2_X1   g438(.A1(new_n578), .A2(new_n577), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n579), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n579), .A2(new_n640), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n613), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n638), .A2(new_n639), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n583), .A2(KEYINPUT10), .A3(new_n613), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(G230gat), .A2(G233gat), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n647), .B1(new_n638), .B2(new_n643), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n636), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(KEYINPUT104), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT104), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n646), .A2(new_n653), .A3(new_n647), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n649), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n651), .B1(new_n655), .B2(new_n636), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AND3_X1   g456(.A1(new_n629), .A2(new_n630), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n496), .A2(new_n570), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n339), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n661), .B(G1gat), .Z(G1324gat));
  INV_X1    g461(.A(KEYINPUT42), .ZN(new_n663));
  INV_X1    g462(.A(new_n402), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n659), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT16), .B(G8gat), .Z(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n663), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n665), .A2(KEYINPUT42), .A3(new_n667), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n666), .A2(G8gat), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(G1325gat));
  OAI21_X1  g471(.A(G15gat), .B1(new_n659), .B2(new_n493), .ZN(new_n673));
  OR2_X1    g472(.A1(new_n462), .A2(G15gat), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n673), .B1(new_n659), .B2(new_n674), .ZN(G1326gat));
  NOR2_X1   g474(.A1(new_n659), .A2(new_n285), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT43), .B(G22gat), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n676), .B(new_n677), .Z(G1327gat));
  INV_X1    g477(.A(KEYINPUT105), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n679), .B1(new_n454), .B2(new_n465), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n449), .A2(new_n452), .A3(KEYINPUT35), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n452), .B1(new_n449), .B2(KEYINPUT35), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n679), .B(new_n465), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n495), .B1(new_n680), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT106), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n495), .B(KEYINPUT106), .C1(new_n680), .C2(new_n684), .ZN(new_n688));
  INV_X1    g487(.A(new_n626), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n600), .B1(new_n596), .B2(new_n598), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n691), .A2(KEYINPUT44), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n687), .A2(new_n688), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n691), .B1(new_n466), .B2(new_n495), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n625), .A2(new_n569), .A3(new_n656), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(G29gat), .B1(new_n699), .B2(new_n660), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n694), .A2(new_n698), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n701), .A2(G29gat), .A3(new_n660), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n702), .A2(KEYINPUT45), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(KEYINPUT45), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n700), .A2(new_n703), .A3(new_n704), .ZN(G1328gat));
  OAI21_X1  g504(.A(G36gat), .B1(new_n699), .B2(new_n664), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n701), .A2(G36gat), .A3(new_n664), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT46), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(G1329gat));
  NOR3_X1   g508(.A1(new_n701), .A2(G43gat), .A3(new_n462), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT47), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n493), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n697), .A2(new_n713), .A3(new_n698), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n715));
  OAI21_X1  g514(.A(G43gat), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n699), .A2(KEYINPUT108), .A3(new_n493), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n712), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(G43gat), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n710), .B(KEYINPUT107), .Z(new_n721));
  OAI21_X1  g520(.A(new_n711), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n718), .A2(new_n722), .ZN(G1330gat));
  OAI21_X1  g522(.A(G50gat), .B1(new_n699), .B2(new_n285), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT110), .ZN(new_n725));
  INV_X1    g524(.A(new_n285), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n203), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT109), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n694), .A2(new_n698), .A3(new_n728), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n697), .A2(new_n726), .A3(new_n698), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(new_n730), .B2(new_n203), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT48), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n725), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n724), .B(new_n729), .C1(KEYINPUT110), .C2(KEYINPUT48), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(G1331gat));
  AND2_X1   g534(.A1(new_n687), .A2(new_n688), .ZN(new_n736));
  AND4_X1   g535(.A1(new_n569), .A2(new_n629), .A3(new_n630), .A4(new_n656), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n339), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n402), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n742));
  XOR2_X1   g541(.A(KEYINPUT49), .B(G64gat), .Z(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n741), .B2(new_n743), .ZN(G1333gat));
  INV_X1    g543(.A(G71gat), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n738), .A2(new_n745), .A3(new_n461), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n736), .A2(new_n713), .A3(new_n737), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G71gat), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT50), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(G1334gat));
  NAND2_X1  g550(.A1(new_n738), .A2(new_n726), .ZN(new_n752));
  XNOR2_X1  g551(.A(KEYINPUT111), .B(G78gat), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1335gat));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755));
  INV_X1    g554(.A(new_n685), .ZN(new_n756));
  INV_X1    g555(.A(new_n691), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n570), .A2(new_n625), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n755), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n756), .A2(new_n755), .A3(new_n759), .ZN(new_n762));
  OR2_X1    g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n763), .A2(new_n574), .A3(new_n339), .A4(new_n656), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n697), .A2(new_n656), .A3(new_n758), .ZN(new_n765));
  OAI21_X1  g564(.A(G85gat), .B1(new_n765), .B2(new_n660), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(G1336gat));
  NAND4_X1  g566(.A1(new_n697), .A2(new_n402), .A3(new_n656), .A4(new_n758), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G92gat), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n657), .A2(new_n664), .A3(G92gat), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n763), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n769), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n770), .B(KEYINPUT112), .ZN(new_n774));
  AOI22_X1  g573(.A1(new_n763), .A2(new_n774), .B1(new_n768), .B2(G92gat), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n773), .B1(new_n775), .B2(new_n776), .ZN(G1337gat));
  OAI21_X1  g576(.A(G99gat), .B1(new_n765), .B2(new_n493), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n462), .A2(G99gat), .A3(new_n657), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(G1338gat));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n758), .A2(new_n656), .ZN(new_n783));
  AOI211_X1 g582(.A(new_n285), .B(new_n783), .C1(new_n693), .C2(new_n696), .ZN(new_n784));
  INV_X1    g583(.A(G106gat), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n782), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n285), .A2(G106gat), .A3(new_n657), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(new_n761), .B2(new_n762), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n788), .B1(new_n784), .B2(new_n785), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n786), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  OAI221_X1 g590(.A(new_n788), .B1(new_n782), .B2(KEYINPUT53), .C1(new_n784), .C2(new_n785), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(G1339gat));
  INV_X1    g592(.A(KEYINPUT117), .ZN(new_n794));
  AND4_X1   g593(.A1(new_n569), .A2(new_n629), .A3(new_n630), .A4(new_n657), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n797));
  INV_X1    g596(.A(new_n551), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n798), .A2(new_n549), .A3(new_n548), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n797), .B1(new_n799), .B2(new_n547), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n550), .A2(new_n551), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n801), .A2(KEYINPUT115), .A3(new_n546), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n540), .A2(new_n542), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n800), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n559), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n565), .A2(new_n552), .A3(new_n554), .A4(new_n560), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n805), .A2(new_n806), .A3(new_n656), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n809));
  AND3_X1   g608(.A1(new_n652), .A2(new_n809), .A3(new_n654), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n648), .A2(KEYINPUT54), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n646), .A2(new_n647), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n635), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n808), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n652), .A2(new_n809), .A3(new_n654), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n809), .B1(new_n646), .B2(new_n647), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n816), .B1(new_n647), .B2(new_n646), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n815), .A2(KEYINPUT55), .A3(new_n635), .A4(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n814), .A2(new_n651), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n807), .B1(new_n569), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n820), .A2(new_n626), .A3(new_n602), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n689), .B2(new_n690), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n796), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(new_n625), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n821), .A2(new_n824), .A3(new_n796), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n795), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n794), .B1(new_n828), .B2(new_n726), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n660), .A2(new_n402), .ZN(new_n830));
  INV_X1    g629(.A(new_n827), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n831), .A2(new_n825), .A3(new_n625), .ZN(new_n832));
  OAI211_X1 g631(.A(KEYINPUT117), .B(new_n285), .C1(new_n832), .C2(new_n795), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n829), .A2(new_n461), .A3(new_n830), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT118), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n285), .B1(new_n832), .B2(new_n795), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n462), .B1(new_n836), .B2(new_n794), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n837), .A2(new_n838), .A3(new_n830), .A4(new_n833), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n835), .A2(new_n839), .A3(new_n570), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(G113gat), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n569), .A2(G113gat), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n339), .B1(new_n832), .B2(new_n795), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n285), .A2(new_n448), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n402), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n847), .A2(KEYINPUT119), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n847), .A2(KEYINPUT119), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n842), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n841), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT120), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n841), .A2(new_n853), .A3(new_n850), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(G1340gat));
  NAND3_X1  g654(.A1(new_n835), .A2(new_n839), .A3(new_n656), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(G120gat), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n657), .A2(G120gat), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n858), .B1(new_n848), .B2(new_n849), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(G1341gat));
  AND3_X1   g659(.A1(new_n835), .A2(new_n839), .A3(new_n625), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n625), .A2(new_n617), .ZN(new_n862));
  OAI22_X1  g661(.A1(new_n861), .A2(new_n617), .B1(new_n847), .B2(new_n862), .ZN(G1342gat));
  NOR3_X1   g662(.A1(new_n847), .A2(G134gat), .A3(new_n691), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT56), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n835), .A2(new_n839), .A3(new_n757), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(G134gat), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(G1343gat));
  AND2_X1   g667(.A1(new_n493), .A2(new_n830), .ZN(new_n869));
  INV_X1    g668(.A(new_n795), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n821), .A2(new_n824), .ZN(new_n871));
  INV_X1    g670(.A(new_n625), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n285), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n869), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n828), .A2(KEYINPUT57), .A3(new_n285), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(G141gat), .A3(new_n570), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n844), .A2(KEYINPUT121), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n713), .A2(new_n402), .A3(new_n285), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT121), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n843), .B2(new_n882), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n880), .A2(new_n883), .A3(new_n569), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n879), .B1(new_n884), .B2(G141gat), .ZN(new_n885));
  XNOR2_X1  g684(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n886));
  XOR2_X1   g685(.A(new_n885), .B(new_n886), .Z(G1344gat));
  INV_X1    g686(.A(new_n878), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(new_n657), .ZN(new_n889));
  OAI21_X1  g688(.A(KEYINPUT57), .B1(new_n828), .B2(new_n285), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XOR2_X1   g691(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n893));
  NOR2_X1   g692(.A1(new_n657), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n869), .A2(new_n894), .ZN(new_n895));
  OAI22_X1  g694(.A1(new_n889), .A2(KEYINPUT59), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n883), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n656), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n893), .A2(G148gat), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n896), .A2(G148gat), .B1(new_n898), .B2(new_n899), .ZN(G1345gat));
  OAI21_X1  g699(.A(G155gat), .B1(new_n888), .B2(new_n872), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n897), .A2(new_n234), .A3(new_n625), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1346gat));
  NOR3_X1   g702(.A1(new_n888), .A2(new_n235), .A3(new_n691), .ZN(new_n904));
  AOI21_X1  g703(.A(G162gat), .B1(new_n897), .B2(new_n757), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n904), .A2(new_n905), .ZN(G1347gat));
  NOR2_X1   g705(.A1(new_n664), .A2(new_n339), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n837), .A2(new_n833), .A3(new_n907), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n908), .A2(new_n354), .A3(new_n569), .ZN(new_n909));
  NOR4_X1   g708(.A1(new_n828), .A2(new_n339), .A3(new_n664), .A4(new_n845), .ZN(new_n910));
  AOI21_X1  g709(.A(G169gat), .B1(new_n910), .B2(new_n570), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n909), .A2(new_n911), .ZN(G1348gat));
  OAI21_X1  g711(.A(G176gat), .B1(new_n908), .B2(new_n657), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n910), .A2(new_n355), .A3(new_n656), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1349gat));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n916), .A2(KEYINPUT60), .ZN(new_n917));
  OAI21_X1  g716(.A(G183gat), .B1(new_n908), .B2(new_n872), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n910), .A2(new_n376), .A3(new_n378), .A4(new_n625), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n916), .A2(KEYINPUT60), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n920), .B(new_n921), .ZN(G1350gat));
  NAND3_X1  g721(.A1(new_n910), .A2(new_n349), .A3(new_n757), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n908), .A2(new_n691), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT61), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n924), .A2(new_n925), .A3(G190gat), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n925), .B1(new_n924), .B2(G190gat), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(G1351gat));
  NAND2_X1  g727(.A1(new_n493), .A2(new_n907), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(G197gat), .A3(new_n570), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n892), .A2(KEYINPUT125), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n892), .A2(KEYINPUT125), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n828), .A2(new_n339), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n713), .A2(new_n664), .A3(new_n285), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(G197gat), .B1(new_n938), .B2(new_n570), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n934), .A2(new_n939), .ZN(G1352gat));
  NOR3_X1   g739(.A1(new_n937), .A2(G204gat), .A3(new_n657), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT62), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n930), .A2(new_n656), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n943), .B1(new_n932), .B2(new_n933), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n944), .A2(KEYINPUT126), .ZN(new_n945));
  OAI21_X1  g744(.A(G204gat), .B1(new_n944), .B2(KEYINPUT126), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n942), .B1(new_n945), .B2(new_n946), .ZN(G1353gat));
  NAND3_X1  g746(.A1(new_n938), .A2(new_n218), .A3(new_n625), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n890), .A2(new_n891), .A3(new_n625), .A4(new_n930), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n949), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n950));
  AOI21_X1  g749(.A(KEYINPUT63), .B1(new_n949), .B2(G211gat), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(G1354gat));
  NAND3_X1  g751(.A1(new_n930), .A2(G218gat), .A3(new_n757), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n953), .B1(new_n932), .B2(new_n933), .ZN(new_n954));
  AOI21_X1  g753(.A(G218gat), .B1(new_n938), .B2(new_n757), .ZN(new_n955));
  OR3_X1    g754(.A1(new_n954), .A2(KEYINPUT127), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(KEYINPUT127), .B1(new_n954), .B2(new_n955), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(G1355gat));
endmodule


