//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072;
  XNOR2_X1  g000(.A(G125), .B(G140), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  AND3_X1   g002(.A1(new_n187), .A2(KEYINPUT80), .A3(new_n188), .ZN(new_n189));
  AOI21_X1  g003(.A(KEYINPUT80), .B1(new_n187), .B2(new_n188), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G125), .ZN(new_n193));
  INV_X1    g007(.A(G125), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G140), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n193), .A2(new_n195), .A3(KEYINPUT78), .ZN(new_n196));
  OR3_X1    g010(.A1(new_n194), .A2(KEYINPUT78), .A3(G140), .ZN(new_n197));
  AND3_X1   g011(.A1(new_n196), .A2(KEYINPUT94), .A3(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(KEYINPUT94), .B1(new_n196), .B2(new_n197), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n191), .B1(new_n200), .B2(G146), .ZN(new_n201));
  INV_X1    g015(.A(G953), .ZN(new_n202));
  AND2_X1   g016(.A1(KEYINPUT67), .A2(G237), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT67), .A2(G237), .ZN(new_n204));
  OAI211_X1 g018(.A(G214), .B(new_n202), .C1(new_n203), .C2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(G237), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n208), .A2(G143), .A3(G214), .A4(new_n202), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT18), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  NOR3_X1   g026(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT93), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(new_n213), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n207), .A2(new_n209), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  OR2_X1    g031(.A1(new_n201), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n210), .A2(G131), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT96), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n210), .A2(KEYINPUT96), .A3(G131), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT95), .B1(new_n210), .B2(G131), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT95), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n207), .A2(new_n209), .A3(new_n224), .A4(new_n212), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(KEYINPUT17), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n196), .A2(new_n197), .A3(KEYINPUT16), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT16), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n193), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n231), .A2(G146), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n188), .B1(new_n228), .B2(new_n230), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n212), .B1(new_n207), .B2(new_n209), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n235), .B(new_n220), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT17), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n234), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n218), .B1(new_n227), .B2(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(G113), .B(G122), .ZN(new_n240));
  INV_X1    g054(.A(G104), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n242), .B(new_n218), .C1(new_n227), .C2(new_n238), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G902), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G475), .ZN(new_n249));
  INV_X1    g063(.A(G116), .ZN(new_n250));
  OAI21_X1  g064(.A(KEYINPUT100), .B1(new_n250), .B2(G122), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT100), .ZN(new_n252));
  INV_X1    g066(.A(G122), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(G116), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G107), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n250), .A2(G122), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n206), .A2(G128), .ZN(new_n259));
  INV_X1    g073(.A(G128), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G143), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G134), .ZN(new_n263));
  INV_X1    g077(.A(G134), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n259), .A2(new_n261), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n257), .A2(KEYINPUT14), .ZN(new_n267));
  OR3_X1    g081(.A1(new_n253), .A2(KEYINPUT14), .A3(G116), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n255), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n258), .B(new_n266), .C1(new_n269), .C2(new_n256), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT13), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n261), .B1(new_n259), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n259), .A2(new_n271), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT101), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n259), .A2(KEYINPUT101), .A3(new_n271), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n272), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n265), .B1(new_n277), .B2(new_n264), .ZN(new_n278));
  INV_X1    g092(.A(new_n258), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n256), .B1(new_n255), .B2(new_n257), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n270), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(KEYINPUT9), .B(G234), .ZN(new_n283));
  INV_X1    g097(.A(G217), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n283), .A2(new_n284), .A3(G953), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n270), .B(new_n285), .C1(new_n278), .C2(new_n281), .ZN(new_n288));
  AOI21_X1  g102(.A(G902), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G478), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(KEYINPUT15), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  AOI211_X1 g107(.A(G902), .B(new_n291), .C1(new_n287), .C2(new_n288), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n202), .A2(G952), .ZN(new_n296));
  NAND2_X1  g110(.A1(G234), .A2(G237), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n297), .A2(G902), .A3(G953), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT21), .B(G898), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n295), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  AND4_X1   g119(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n225), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n196), .A2(new_n197), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT94), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n196), .A2(new_n197), .A3(KEYINPUT94), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(KEYINPUT19), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n193), .A2(new_n195), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n311), .B(new_n188), .C1(KEYINPUT19), .C2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n233), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n218), .B(KEYINPUT97), .C1(new_n306), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n243), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n201), .A2(new_n217), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n312), .A2(KEYINPUT19), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n319), .B1(new_n200), .B2(KEYINPUT19), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n233), .B1(new_n320), .B2(new_n188), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n318), .B1(new_n321), .B2(new_n226), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n322), .A2(KEYINPUT97), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n245), .B1(new_n317), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT99), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT20), .ZN(new_n327));
  NOR2_X1   g141(.A1(G475), .A2(G902), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(KEYINPUT98), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  AOI22_X1  g144(.A1(new_n326), .A2(new_n327), .B1(new_n324), .B2(new_n330), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n324), .A2(KEYINPUT99), .A3(new_n327), .A4(new_n330), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n249), .B(new_n305), .C1(new_n331), .C2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(G210), .B1(G237), .B2(G902), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n241), .A2(KEYINPUT85), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT85), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G104), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(new_n338), .A3(G107), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT3), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(new_n256), .A3(G104), .ZN(new_n341));
  AOI21_X1  g155(.A(G107), .B1(new_n336), .B2(new_n338), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n339), .B(new_n341), .C1(new_n342), .C2(new_n340), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G101), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT85), .B(G104), .ZN(new_n345));
  OAI21_X1  g159(.A(KEYINPUT3), .B1(new_n345), .B2(G107), .ZN(new_n346));
  INV_X1    g160(.A(G101), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n346), .A2(new_n347), .A3(new_n339), .A4(new_n341), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n344), .A2(KEYINPUT4), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT66), .ZN(new_n350));
  INV_X1    g164(.A(G119), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G116), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n250), .A2(G119), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT2), .B(G113), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n350), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(G116), .B(G119), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT2), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n358), .A2(G113), .ZN(new_n359));
  INV_X1    g173(.A(G113), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(KEYINPUT2), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n357), .B(KEYINPUT66), .C1(new_n359), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n356), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n354), .A2(new_n355), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n347), .A2(KEYINPUT4), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n363), .A2(new_n364), .B1(new_n343), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n349), .A2(new_n366), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT5), .ZN(new_n368));
  OAI21_X1  g182(.A(G113), .B1(new_n352), .B2(KEYINPUT5), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT90), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n370), .A2(new_n371), .B1(new_n356), .B2(new_n362), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n256), .A2(G104), .ZN(new_n373));
  OAI21_X1  g187(.A(G101), .B1(new_n342), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT90), .B1(new_n368), .B2(new_n369), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n372), .A2(new_n348), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n367), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(G110), .B(G122), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n367), .A2(new_n378), .A3(new_n376), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(KEYINPUT6), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT6), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n377), .A2(new_n383), .A3(new_n379), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n260), .A2(KEYINPUT1), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n188), .A2(G143), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n206), .A2(G146), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n188), .A2(KEYINPUT64), .A3(G143), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT64), .B1(new_n188), .B2(G143), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n389), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n260), .B1(new_n386), .B2(KEYINPUT1), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n194), .B(new_n388), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n188), .A2(KEYINPUT64), .A3(G143), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT64), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n395), .B1(new_n206), .B2(G146), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n206), .A2(G146), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n394), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  AND2_X1   g212(.A1(KEYINPUT0), .A2(G128), .ZN(new_n399));
  NOR2_X1   g213(.A1(KEYINPUT0), .A2(G128), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n386), .A2(new_n387), .ZN(new_n402));
  AOI22_X1  g216(.A1(new_n398), .A2(new_n401), .B1(new_n402), .B2(new_n399), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n393), .B1(new_n194), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n202), .A2(G224), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n404), .B(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n382), .A2(new_n384), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n348), .A2(new_n374), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n409), .A2(new_n372), .A3(new_n375), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n378), .B(KEYINPUT8), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n357), .A2(KEYINPUT5), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT91), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n369), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n368), .A2(KEYINPUT91), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n414), .A2(new_n415), .B1(new_n356), .B2(new_n362), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n411), .B1(new_n416), .B2(new_n409), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n410), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT7), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n404), .B1(new_n419), .B2(new_n406), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n406), .A2(new_n419), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n393), .B(new_n421), .C1(new_n194), .C2(new_n403), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(G902), .B1(new_n424), .B2(new_n381), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n335), .B1(new_n408), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n408), .A2(new_n335), .A3(new_n425), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(KEYINPUT92), .A3(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(G214), .B1(G237), .B2(G902), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT92), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n429), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n334), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT22), .B(G137), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n202), .A2(G221), .A3(G234), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n435), .B(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n233), .A2(new_n191), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT24), .B(G110), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(KEYINPUT74), .B1(new_n260), .B2(G119), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT74), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(new_n351), .A3(G128), .ZN(new_n445));
  AOI22_X1  g259(.A1(new_n443), .A2(new_n445), .B1(G119), .B2(new_n260), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT75), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n446), .A2(KEYINPUT75), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n442), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OR2_X1    g265(.A1(new_n451), .A2(KEYINPUT79), .ZN(new_n452));
  INV_X1    g266(.A(G110), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n260), .A2(KEYINPUT23), .A3(G119), .ZN(new_n454));
  XOR2_X1   g268(.A(new_n454), .B(KEYINPUT76), .Z(new_n455));
  OR3_X1    g269(.A1(new_n351), .A2(KEYINPUT77), .A3(G128), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT77), .B1(new_n351), .B2(G128), .ZN(new_n457));
  OAI21_X1  g271(.A(KEYINPUT23), .B1(new_n260), .B2(G119), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n451), .A2(KEYINPUT79), .B1(new_n453), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n440), .B1(new_n452), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n449), .A2(new_n450), .A3(new_n442), .ZN(new_n463));
  OAI21_X1  g277(.A(G110), .B1(new_n455), .B2(new_n459), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n463), .B(new_n464), .C1(new_n232), .C2(new_n233), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n438), .B1(new_n462), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n450), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n446), .A2(KEYINPUT75), .ZN(new_n469));
  OAI211_X1 g283(.A(KEYINPUT79), .B(new_n441), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n460), .A2(new_n453), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n451), .A2(KEYINPUT79), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n439), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(new_n465), .A3(new_n437), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n467), .A2(new_n247), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT25), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n467), .A2(KEYINPUT25), .A3(new_n247), .A4(new_n475), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n284), .B1(G234), .B2(new_n247), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(G902), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n483), .B(KEYINPUT82), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT81), .ZN(new_n486));
  INV_X1    g300(.A(new_n475), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n437), .B1(new_n474), .B2(new_n465), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n467), .A2(KEYINPUT81), .A3(new_n475), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n485), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n482), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT28), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT11), .B1(new_n264), .B2(G137), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT11), .ZN(new_n496));
  INV_X1    g310(.A(G137), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n497), .A3(G134), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT65), .B1(new_n497), .B2(G134), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT65), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(new_n264), .A3(G137), .ZN(new_n502));
  AND4_X1   g316(.A1(new_n212), .A2(new_n499), .A3(new_n500), .A4(new_n502), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n500), .A2(new_n502), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n212), .B1(new_n504), .B2(new_n499), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n403), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n504), .A2(new_n212), .A3(new_n499), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n497), .A2(G134), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n264), .A2(G137), .ZN(new_n509));
  OAI21_X1  g323(.A(G131), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n390), .A2(new_n386), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n392), .B1(new_n511), .B2(new_n394), .ZN(new_n512));
  INV_X1    g326(.A(new_n388), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n507), .B(new_n510), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n506), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n356), .A2(new_n362), .B1(new_n354), .B2(new_n355), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n506), .A2(new_n516), .A3(new_n514), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n494), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n494), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n208), .A2(G210), .A3(new_n202), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT27), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT27), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n208), .A2(new_n526), .A3(G210), .A4(new_n202), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT26), .B(G101), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n528), .B1(new_n525), .B2(new_n527), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT29), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(G902), .B1(new_n523), .B2(new_n535), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n506), .A2(new_n516), .A3(new_n514), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n515), .A2(KEYINPUT30), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT30), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n506), .A2(new_n539), .A3(new_n514), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n537), .B1(new_n541), .B2(new_n517), .ZN(new_n542));
  OAI21_X1  g356(.A(KEYINPUT73), .B1(new_n542), .B2(new_n532), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n506), .A2(new_n539), .A3(new_n514), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n539), .B1(new_n506), .B2(new_n514), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n517), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n519), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT73), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n548), .A3(new_n533), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n543), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n516), .B1(new_n506), .B2(new_n514), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT28), .B1(new_n537), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT69), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n553), .B1(new_n530), .B2(new_n531), .ZN(new_n554));
  INV_X1    g368(.A(new_n531), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(KEYINPUT69), .A3(new_n529), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n552), .A2(new_n557), .A3(new_n521), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT72), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT72), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n552), .A2(new_n557), .A3(new_n560), .A4(new_n521), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n559), .A2(new_n534), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n536), .B1(new_n550), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(G472), .A2(G902), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n554), .A2(new_n556), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n566), .B1(new_n520), .B2(new_n522), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT68), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(KEYINPUT31), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n546), .A2(new_n519), .A3(new_n532), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n546), .A2(KEYINPUT68), .A3(new_n519), .A4(new_n532), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT31), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n565), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n563), .A2(G472), .B1(new_n575), .B2(KEYINPUT32), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n573), .A2(KEYINPUT31), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n564), .B1(new_n577), .B2(new_n571), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT70), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n574), .A2(new_n567), .A3(new_n570), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT70), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(new_n581), .A3(new_n564), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT71), .B(KEYINPUT32), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n579), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n493), .B1(new_n576), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(G221), .B1(new_n283), .B2(G902), .ZN(new_n586));
  XOR2_X1   g400(.A(new_n586), .B(KEYINPUT83), .Z(new_n587));
  INV_X1    g401(.A(G469), .ZN(new_n588));
  XNOR2_X1  g402(.A(G110), .B(G140), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n202), .A2(G227), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n503), .A2(new_n505), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n343), .A2(G101), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n341), .B1(new_n342), .B2(new_n340), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n339), .A2(new_n347), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT4), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n343), .A2(new_n365), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n403), .ZN(new_n599));
  OAI21_X1  g413(.A(KEYINPUT86), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n598), .A2(new_n403), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT86), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n602), .A3(new_n349), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n388), .B1(new_n402), .B2(new_n392), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n605), .B(new_n374), .C1(new_n594), .C2(new_n595), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT87), .B(KEYINPUT10), .Z(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n388), .B1(new_n391), .B2(new_n392), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n609), .A2(new_n348), .A3(KEYINPUT10), .A4(new_n374), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n592), .B1(new_n604), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n592), .ZN(new_n614));
  AOI211_X1 g428(.A(new_n614), .B(new_n611), .C1(new_n600), .C2(new_n603), .ZN(new_n615));
  OAI211_X1 g429(.A(KEYINPUT89), .B(new_n591), .C1(new_n613), .C2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n611), .B1(new_n600), .B2(new_n603), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n591), .B1(new_n617), .B2(new_n592), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n348), .A2(new_n374), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n606), .B1(new_n619), .B2(new_n609), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT88), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n620), .A2(new_n621), .A3(KEYINPUT12), .A4(new_n614), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n609), .B1(new_n348), .B2(new_n374), .ZN(new_n623));
  INV_X1    g437(.A(new_n606), .ZN(new_n624));
  OAI211_X1 g438(.A(KEYINPUT12), .B(new_n614), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(KEYINPUT88), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n620), .A2(new_n614), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n622), .B(new_n626), .C1(new_n627), .C2(KEYINPUT12), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n618), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n616), .A2(new_n629), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n601), .A2(new_n602), .A3(new_n349), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n602), .B1(new_n601), .B2(new_n349), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n612), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n614), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n617), .A2(new_n592), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(KEYINPUT89), .B1(new_n636), .B2(new_n591), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n588), .B(new_n247), .C1(new_n630), .C2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n628), .A2(new_n635), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n591), .B(KEYINPUT84), .ZN(new_n640));
  AOI22_X1  g454(.A1(new_n639), .A2(new_n640), .B1(new_n634), .B2(new_n618), .ZN(new_n641));
  OAI21_X1  g455(.A(G469), .B1(new_n641), .B2(G902), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n587), .B1(new_n638), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n434), .A2(new_n585), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G101), .ZN(G3));
  INV_X1    g459(.A(G475), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(new_n246), .B2(new_n247), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n324), .A2(new_n330), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n242), .B1(new_n322), .B2(KEYINPUT97), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n218), .B1(new_n306), .B2(new_n315), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT97), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(KEYINPUT99), .B1(new_n653), .B2(new_n245), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n648), .B1(new_n654), .B2(KEYINPUT20), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n647), .B1(new_n655), .B2(new_n332), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT102), .B(KEYINPUT33), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT33), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(KEYINPUT102), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n287), .A2(new_n288), .ZN(new_n660));
  MUX2_X1   g474(.A(new_n657), .B(new_n659), .S(new_n660), .Z(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(G478), .A3(new_n247), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n660), .A2(new_n247), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n290), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n408), .A2(new_n335), .A3(new_n425), .ZN(new_n667));
  OAI211_X1 g481(.A(new_n303), .B(new_n430), .C1(new_n667), .C2(new_n426), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n656), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n580), .A2(new_n247), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(G472), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n579), .A3(new_n582), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n493), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n669), .A2(new_n643), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT34), .B(G104), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G6));
  XNOR2_X1  g490(.A(KEYINPUT103), .B(KEYINPUT20), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n232), .A2(new_n233), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n221), .A2(new_n222), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n678), .B1(KEYINPUT17), .B2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n236), .A2(new_n237), .A3(new_n223), .A4(new_n225), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n318), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  AOI22_X1  g496(.A1(new_n649), .A2(new_n652), .B1(new_n682), .B2(new_n242), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n677), .B1(new_n683), .B2(new_n329), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n327), .A2(KEYINPUT103), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n324), .A2(new_n330), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n295), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n249), .A2(new_n684), .A3(new_n686), .A4(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n668), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n673), .A2(new_n689), .A3(new_n643), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT35), .B(G107), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G9));
  NAND2_X1  g506(.A1(new_n474), .A2(new_n465), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n438), .A2(KEYINPUT36), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(new_n695));
  AOI22_X1  g509(.A1(new_n480), .A2(new_n481), .B1(new_n484), .B2(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n672), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n434), .A2(new_n643), .A3(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT37), .B(G110), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G12));
  OAI21_X1  g514(.A(new_n430), .B1(new_n667), .B2(new_n426), .ZN(new_n701));
  AOI211_X1 g515(.A(new_n587), .B(new_n701), .C1(new_n638), .C2(new_n642), .ZN(new_n702));
  INV_X1    g516(.A(G900), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n299), .B1(new_n300), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n688), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n696), .B1(new_n576), .B2(new_n584), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n702), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G128), .ZN(G30));
  XOR2_X1   g522(.A(new_n704), .B(KEYINPUT39), .Z(new_n709));
  NAND2_X1  g523(.A1(new_n643), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT40), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT40), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n710), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(KEYINPUT105), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n429), .A2(new_n432), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(G472), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n542), .A2(new_n532), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n566), .B1(new_n537), .B2(new_n551), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n720), .B1(new_n723), .B2(new_n247), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n724), .B1(new_n575), .B2(KEYINPUT32), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n584), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n696), .A2(new_n687), .A3(new_n430), .ZN(new_n728));
  NOR4_X1   g542(.A1(new_n719), .A2(new_n727), .A3(new_n656), .A4(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n713), .A2(new_n716), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(KEYINPUT106), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT106), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n713), .A2(new_n716), .A3(new_n732), .A4(new_n729), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n206), .ZN(G45));
  NOR3_X1   g549(.A1(new_n656), .A2(new_n666), .A3(new_n704), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(new_n702), .A3(new_n706), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G146), .ZN(G48));
  OAI21_X1  g552(.A(new_n247), .B1(new_n630), .B2(new_n637), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(G469), .ZN(new_n740));
  INV_X1    g554(.A(new_n587), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n740), .A2(new_n741), .A3(new_n638), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n669), .A2(new_n742), .A3(new_n585), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(KEYINPUT107), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT107), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n669), .A2(new_n742), .A3(new_n585), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(KEYINPUT41), .B(G113), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(G15));
  NAND3_X1  g563(.A1(new_n742), .A2(new_n585), .A3(new_n689), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G116), .ZN(G18));
  INV_X1    g565(.A(new_n334), .ZN(new_n752));
  INV_X1    g566(.A(new_n701), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n742), .A2(new_n752), .A3(new_n706), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G119), .ZN(G21));
  OAI211_X1 g569(.A(new_n687), .B(new_n430), .C1(new_n667), .C2(new_n426), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n656), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n575), .B1(G472), .B2(new_n670), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n491), .B1(new_n480), .B2(new_n481), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n758), .A2(new_n759), .A3(new_n303), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n742), .A2(new_n757), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(KEYINPUT108), .B(G122), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n761), .B(new_n762), .ZN(G24));
  AND4_X1   g577(.A1(new_n741), .A2(new_n740), .A3(new_n638), .A4(new_n753), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n695), .A2(new_n484), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n482), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n758), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n764), .A2(new_n736), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G125), .ZN(G27));
  NAND2_X1  g584(.A1(new_n655), .A2(new_n332), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n249), .ZN(new_n772));
  INV_X1    g586(.A(new_n704), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n665), .A3(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n430), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n775), .B1(new_n429), .B2(new_n432), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n643), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n576), .B1(KEYINPUT32), .B2(new_n575), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n759), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n778), .A2(KEYINPUT42), .A3(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT109), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n783), .B1(new_n778), .B2(new_n585), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n643), .A2(new_n776), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n785), .A2(new_n783), .A3(new_n736), .A4(new_n585), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT42), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n782), .B1(new_n784), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(KEYINPUT110), .B(G131), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n789), .B(new_n790), .ZN(G33));
  NAND3_X1  g605(.A1(new_n785), .A2(new_n585), .A3(new_n705), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G134), .ZN(G36));
  INV_X1    g607(.A(new_n638), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT45), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n639), .A2(new_n640), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n613), .A2(new_n615), .A3(new_n591), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n641), .A2(KEYINPUT45), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(G469), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(G469), .A2(G902), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT46), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n794), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n800), .A2(KEYINPUT46), .A3(new_n801), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n741), .A3(new_n709), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT111), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n587), .B1(new_n804), .B2(new_n805), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT111), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(new_n810), .A3(new_n709), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n656), .A2(new_n665), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT43), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n813), .B(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n672), .A2(new_n766), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(KEYINPUT44), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT44), .B1(new_n815), .B2(new_n816), .ZN(new_n818));
  INV_X1    g632(.A(new_n776), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n812), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  XOR2_X1   g635(.A(KEYINPUT112), .B(G137), .Z(new_n822));
  XNOR2_X1  g636(.A(new_n821), .B(new_n822), .ZN(G39));
  XNOR2_X1  g637(.A(new_n809), .B(KEYINPUT47), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n576), .A2(new_n584), .ZN(new_n825));
  NOR4_X1   g639(.A1(new_n774), .A2(new_n819), .A3(new_n825), .A4(new_n759), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G140), .ZN(G42));
  INV_X1    g642(.A(new_n742), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n829), .A2(new_n819), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(new_n759), .A3(new_n299), .A4(new_n727), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n831), .A2(new_n772), .A3(new_n665), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT119), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n719), .B1(new_n833), .B2(KEYINPUT50), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n835), .B1(new_n829), .B2(new_n430), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n742), .A2(KEYINPUT118), .A3(new_n775), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n834), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n815), .A2(new_n299), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n758), .A2(new_n759), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n833), .A2(KEYINPUT50), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n832), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n839), .A2(new_n845), .A3(new_n830), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n815), .A2(new_n299), .ZN(new_n847));
  INV_X1    g661(.A(new_n830), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT120), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n768), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n809), .A2(KEYINPUT47), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n809), .A2(KEYINPUT47), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n740), .A2(new_n638), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n587), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  AOI22_X1  g671(.A1(new_n857), .A2(new_n776), .B1(new_n838), .B2(new_n842), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n839), .A2(new_n840), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n844), .B(new_n851), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT51), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n860), .A2(new_n861), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n850), .A2(new_n781), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n850), .A2(KEYINPUT121), .A3(new_n781), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n866), .A2(KEYINPUT48), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n839), .A2(new_n764), .A3(new_n840), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n666), .B1(new_n771), .B2(new_n249), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n869), .B(new_n296), .C1(new_n871), .C2(new_n831), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT121), .B1(new_n850), .B2(new_n781), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT48), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n862), .A2(new_n863), .A3(new_n868), .A4(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT53), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n754), .A2(new_n750), .A3(new_n761), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n878), .B1(new_n746), .B2(new_n744), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n663), .A2(new_n291), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n289), .A2(new_n292), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n880), .A2(KEYINPUT114), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT114), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n883), .B1(new_n293), .B2(new_n294), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n249), .B(new_n885), .C1(new_n331), .C2(new_n333), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n886), .B1(new_n656), .B2(new_n666), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n433), .A2(new_n302), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n887), .A2(new_n643), .A3(new_n673), .A4(new_n888), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n889), .A2(new_n644), .A3(new_n698), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n825), .A2(new_n643), .A3(new_n759), .A4(new_n776), .ZN(new_n891));
  INV_X1    g705(.A(new_n705), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n882), .A2(new_n884), .A3(new_n773), .ZN(new_n893));
  AND4_X1   g707(.A1(new_n249), .A2(new_n684), .A3(new_n893), .A4(new_n686), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n579), .A2(new_n582), .A3(new_n583), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n580), .A2(KEYINPUT32), .A3(new_n564), .ZN(new_n896));
  INV_X1    g710(.A(new_n536), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n559), .A2(new_n534), .A3(new_n561), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n548), .B1(new_n547), .B2(new_n533), .ZN(new_n899));
  AOI211_X1 g713(.A(KEYINPUT73), .B(new_n532), .C1(new_n546), .C2(new_n519), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n897), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n896), .B1(new_n902), .B2(new_n720), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n894), .B(new_n766), .C1(new_n895), .C2(new_n903), .ZN(new_n904));
  OAI22_X1  g718(.A1(new_n891), .A2(new_n892), .B1(new_n904), .B2(new_n777), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT115), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n870), .A2(new_n643), .A3(new_n773), .A4(new_n776), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n906), .B1(new_n907), .B2(new_n767), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n785), .A2(KEYINPUT115), .A3(new_n736), .A4(new_n768), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n789), .A2(new_n879), .A3(new_n890), .A4(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n766), .A2(new_n704), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n757), .A2(new_n726), .A3(new_n643), .A4(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n769), .A2(new_n737), .A3(new_n707), .A4(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(KEYINPUT52), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n706), .B(new_n702), .C1(new_n736), .C2(new_n705), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT52), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n916), .A2(new_n917), .A3(new_n769), .A4(new_n913), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n877), .B1(new_n911), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT54), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT117), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n915), .A2(KEYINPUT117), .A3(new_n918), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n878), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n890), .A2(new_n926), .A3(new_n747), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n927), .A2(KEYINPUT53), .A3(new_n789), .A4(new_n910), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n920), .B(new_n921), .C1(new_n925), .C2(new_n928), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n911), .A2(new_n877), .A3(new_n919), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n915), .A2(KEYINPUT117), .A3(new_n918), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT117), .B1(new_n915), .B2(new_n918), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n910), .A2(new_n747), .A3(new_n890), .A4(new_n926), .ZN(new_n934));
  INV_X1    g748(.A(new_n782), .ZN(new_n935));
  INV_X1    g749(.A(new_n788), .ZN(new_n936));
  INV_X1    g750(.A(new_n585), .ZN(new_n937));
  OAI21_X1  g751(.A(KEYINPUT109), .B1(new_n907), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n935), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(KEYINPUT116), .B1(new_n934), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT116), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n927), .A2(new_n941), .A3(new_n789), .A4(new_n910), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n933), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n930), .B1(new_n943), .B2(new_n877), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n929), .B1(new_n944), .B2(new_n921), .ZN(new_n945));
  OAI22_X1  g759(.A1(new_n876), .A2(new_n945), .B1(G952), .B2(G953), .ZN(new_n946));
  NOR4_X1   g760(.A1(new_n813), .A2(new_n493), .A3(new_n587), .A4(new_n775), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT49), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n947), .B1(new_n948), .B2(new_n855), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT113), .Z(new_n950));
  NAND2_X1  g764(.A1(new_n855), .A2(new_n948), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n719), .A2(new_n951), .A3(new_n727), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n946), .B1(new_n950), .B2(new_n952), .ZN(G75));
  NOR2_X1   g767(.A1(new_n202), .A2(G952), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n925), .A2(new_n928), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n934), .A2(new_n939), .ZN(new_n957));
  INV_X1    g771(.A(new_n919), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT53), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n960), .A2(new_n247), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT56), .B1(new_n961), .B2(G210), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n382), .A2(new_n384), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(new_n407), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT55), .Z(new_n965));
  OAI21_X1  g779(.A(new_n955), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n920), .B1(new_n925), .B2(new_n928), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT122), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n967), .A2(new_n968), .A3(G902), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n968), .B1(new_n967), .B2(G902), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n335), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT56), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n965), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n966), .B1(new_n973), .B2(new_n975), .ZN(G51));
  NOR2_X1   g790(.A1(new_n630), .A2(new_n637), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n967), .A2(KEYINPUT54), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n929), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n801), .B(KEYINPUT57), .Z(new_n980));
  AOI21_X1  g794(.A(new_n977), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT123), .ZN(new_n982));
  INV_X1    g796(.A(new_n800), .ZN(new_n983));
  AOI22_X1  g797(.A1(new_n981), .A2(new_n982), .B1(new_n971), .B2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n980), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n985), .B1(new_n978), .B2(new_n929), .ZN(new_n986));
  OAI21_X1  g800(.A(KEYINPUT123), .B1(new_n986), .B2(new_n977), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n954), .B1(new_n984), .B2(new_n987), .ZN(G54));
  INV_X1    g802(.A(new_n970), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n967), .A2(new_n968), .A3(G902), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n989), .A2(KEYINPUT58), .A3(G475), .A4(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n683), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n971), .A2(KEYINPUT58), .A3(G475), .A4(new_n324), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n992), .A2(new_n993), .A3(new_n955), .ZN(G60));
  NAND2_X1  g808(.A1(G478), .A2(G902), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT59), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n661), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n954), .B1(new_n979), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n661), .B1(new_n945), .B2(new_n996), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n998), .B1(new_n999), .B2(KEYINPUT124), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT124), .ZN(new_n1001));
  AOI211_X1 g815(.A(new_n1001), .B(new_n661), .C1(new_n945), .C2(new_n996), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n1000), .A2(new_n1002), .ZN(G63));
  INV_X1    g817(.A(KEYINPUT125), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT61), .ZN(new_n1005));
  NAND2_X1  g819(.A1(G217), .A2(G902), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(KEYINPUT60), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n967), .A2(new_n695), .A3(new_n1008), .ZN(new_n1009));
  AND2_X1   g823(.A1(new_n1009), .A2(new_n955), .ZN(new_n1010));
  OAI211_X1 g824(.A(new_n490), .B(new_n489), .C1(new_n960), .C2(new_n1007), .ZN(new_n1011));
  AOI211_X1 g825(.A(new_n1004), .B(new_n1005), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1011), .A2(new_n955), .A3(new_n1009), .ZN(new_n1013));
  AOI21_X1  g827(.A(KEYINPUT61), .B1(new_n1013), .B2(KEYINPUT125), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1012), .A2(new_n1014), .ZN(G66));
  INV_X1    g829(.A(new_n301), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n202), .B1(new_n1016), .B2(G224), .ZN(new_n1017));
  INV_X1    g831(.A(new_n927), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1017), .B1(new_n1018), .B2(new_n202), .ZN(new_n1019));
  INV_X1    g833(.A(G898), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n963), .B1(new_n1020), .B2(G953), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1019), .B(new_n1021), .ZN(G69));
  INV_X1    g836(.A(KEYINPUT127), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n781), .A2(new_n757), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1023), .B1(new_n812), .B2(new_n1025), .ZN(new_n1026));
  AOI211_X1 g840(.A(KEYINPUT127), .B(new_n1024), .C1(new_n808), .C2(new_n811), .ZN(new_n1027));
  OR2_X1    g841(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AND2_X1   g842(.A1(new_n916), .A2(new_n769), .ZN(new_n1029));
  AND2_X1   g843(.A1(new_n1029), .A2(new_n792), .ZN(new_n1030));
  AND3_X1   g844(.A1(new_n827), .A2(new_n789), .A3(new_n1030), .ZN(new_n1031));
  NAND4_X1  g845(.A1(new_n1028), .A2(new_n1031), .A3(new_n202), .A4(new_n821), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n541), .B(new_n320), .ZN(new_n1033));
  NAND2_X1  g847(.A1(G900), .A2(G953), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1035), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1032), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g851(.A(KEYINPUT126), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n887), .A2(new_n709), .ZN(new_n1039));
  NOR2_X1   g853(.A1(new_n1039), .A2(new_n891), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1040), .B1(new_n824), .B2(new_n826), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1041), .A2(new_n821), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n731), .A2(new_n1029), .A3(new_n733), .ZN(new_n1043));
  AOI21_X1  g857(.A(new_n1042), .B1(KEYINPUT62), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g858(.A(KEYINPUT62), .ZN(new_n1045));
  NAND4_X1  g859(.A1(new_n731), .A2(new_n1029), .A3(new_n1045), .A4(new_n733), .ZN(new_n1046));
  AOI21_X1  g860(.A(G953), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g861(.A(new_n1037), .B(new_n1038), .C1(new_n1047), .C2(new_n1033), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n1043), .A2(KEYINPUT62), .ZN(new_n1049));
  AND2_X1   g863(.A1(new_n1041), .A2(new_n821), .ZN(new_n1050));
  NAND3_X1  g864(.A1(new_n1049), .A2(new_n1050), .A3(new_n1046), .ZN(new_n1051));
  AOI21_X1  g865(.A(new_n1033), .B1(new_n1051), .B2(new_n202), .ZN(new_n1052));
  NOR2_X1   g866(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1053));
  NAND4_X1  g867(.A1(new_n821), .A2(new_n789), .A3(new_n827), .A4(new_n1030), .ZN(new_n1054));
  NOR2_X1   g868(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g869(.A(new_n1035), .B1(new_n1055), .B2(new_n202), .ZN(new_n1056));
  OAI21_X1  g870(.A(KEYINPUT126), .B1(new_n1052), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n1048), .A2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g872(.A(new_n202), .B1(G227), .B2(G900), .ZN(new_n1059));
  INV_X1    g873(.A(new_n1059), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g875(.A1(new_n1048), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n1061), .A2(new_n1062), .ZN(G72));
  NAND2_X1  g877(.A1(G472), .A2(G902), .ZN(new_n1064));
  XOR2_X1   g878(.A(new_n1064), .B(KEYINPUT63), .Z(new_n1065));
  INV_X1    g879(.A(new_n1065), .ZN(new_n1066));
  AOI211_X1 g880(.A(new_n1066), .B(new_n944), .C1(new_n901), .C2(new_n721), .ZN(new_n1067));
  NAND3_X1  g881(.A1(new_n1044), .A2(new_n927), .A3(new_n1046), .ZN(new_n1068));
  AOI211_X1 g882(.A(new_n542), .B(new_n533), .C1(new_n1068), .C2(new_n1065), .ZN(new_n1069));
  NOR3_X1   g883(.A1(new_n1053), .A2(new_n1054), .A3(new_n1018), .ZN(new_n1070));
  OAI211_X1 g884(.A(new_n542), .B(new_n533), .C1(new_n1070), .C2(new_n1066), .ZN(new_n1071));
  NAND2_X1  g885(.A1(new_n1071), .A2(new_n955), .ZN(new_n1072));
  NOR3_X1   g886(.A1(new_n1067), .A2(new_n1069), .A3(new_n1072), .ZN(G57));
endmodule


