//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 0 1 1 1 1 1 1 1 0 1 1 1 0 0 0 1 1 1 0 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(G137), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT11), .A3(G134), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n190), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G131), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n189), .A2(new_n192), .A3(new_n195), .A4(new_n190), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n194), .A2(KEYINPUT67), .A3(new_n196), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  AND2_X1   g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT0), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  XOR2_X1   g022(.A(KEYINPUT0), .B(G128), .Z(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(new_n205), .B2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n199), .A2(new_n200), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT68), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT69), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n207), .A2(KEYINPUT1), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(new_n202), .A3(new_n204), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n207), .A2(new_n201), .A3(G143), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n203), .B(G146), .C1(new_n207), .C2(KEYINPUT1), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n190), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n188), .A2(G137), .ZN(new_n221));
  OAI21_X1  g035(.A(G131), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n196), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n214), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n225), .A2(KEYINPUT69), .A3(new_n196), .A4(new_n222), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n199), .A2(KEYINPUT68), .A3(new_n200), .A4(new_n210), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n213), .A2(KEYINPUT30), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT2), .ZN(new_n230));
  INV_X1    g044(.A(G113), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT65), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT65), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(KEYINPUT2), .A3(G113), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n230), .A2(new_n231), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT66), .ZN(new_n238));
  INV_X1    g052(.A(G116), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n238), .B1(new_n239), .B2(G119), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(G119), .ZN(new_n241));
  INV_X1    g055(.A(G119), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(KEYINPUT66), .A3(G116), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n240), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n237), .A2(new_n244), .ZN(new_n245));
  AND2_X1   g059(.A1(new_n240), .A2(new_n243), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n246), .A2(new_n236), .A3(new_n235), .A4(new_n241), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT64), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n223), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n222), .A2(KEYINPUT64), .A3(new_n196), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(new_n225), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n210), .A2(new_n197), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT30), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n249), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n229), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n213), .A2(new_n249), .A3(new_n227), .A4(new_n228), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n260), .B(G101), .ZN(new_n261));
  NOR2_X1   g075(.A1(G237), .A2(G953), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G210), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n261), .B(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT31), .B1(new_n258), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n259), .A2(new_n264), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT31), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n229), .A2(new_n257), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n264), .B(KEYINPUT71), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT28), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n255), .A2(new_n248), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n274), .B1(new_n259), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n219), .A2(new_n223), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n199), .A2(new_n200), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n277), .B1(new_n278), .B2(new_n210), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT28), .B1(new_n279), .B2(new_n249), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n273), .B1(new_n276), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n271), .A2(new_n259), .A3(new_n264), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(KEYINPUT70), .A3(KEYINPUT31), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n268), .A2(new_n272), .A3(new_n281), .A4(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(G472), .A2(G902), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(KEYINPUT32), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n213), .A2(new_n227), .A3(new_n228), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n248), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n259), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n280), .B1(new_n291), .B2(KEYINPUT28), .ZN(new_n292));
  INV_X1    g106(.A(new_n264), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT29), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(G902), .B1(new_n292), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n271), .A2(new_n259), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n293), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n276), .A2(new_n280), .A3(new_n273), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n298), .B1(new_n299), .B2(KEYINPUT72), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n259), .A2(new_n275), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT28), .ZN(new_n302));
  INV_X1    g116(.A(new_n280), .ZN(new_n303));
  INV_X1    g117(.A(new_n273), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n302), .A2(KEYINPUT72), .A3(new_n303), .A4(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n294), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n296), .B1(new_n300), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G472), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT32), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n281), .A2(new_n272), .ZN(new_n310));
  AOI211_X1 g124(.A(new_n267), .B(new_n270), .C1(new_n269), .C2(new_n271), .ZN(new_n311));
  AOI21_X1  g125(.A(KEYINPUT70), .B1(new_n282), .B2(KEYINPUT31), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n285), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n309), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n284), .A2(KEYINPUT73), .A3(KEYINPUT32), .A4(new_n285), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n288), .A2(new_n308), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(G214), .B1(G237), .B2(G902), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(G210), .B1(G237), .B2(G902), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n208), .B(G125), .C1(new_n205), .C2(new_n209), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT83), .ZN(new_n323));
  INV_X1    g137(.A(G125), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n219), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT83), .B1(new_n225), .B2(G125), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n322), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  OR2_X1    g141(.A1(new_n327), .A2(KEYINPUT84), .ZN(new_n328));
  INV_X1    g142(.A(G953), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G224), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n330), .B(KEYINPUT85), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n327), .A2(KEYINPUT84), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n328), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n331), .B1(new_n328), .B2(new_n332), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G104), .ZN(new_n336));
  OAI21_X1  g150(.A(KEYINPUT3), .B1(new_n336), .B2(G107), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT3), .ZN(new_n338));
  INV_X1    g152(.A(G107), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n339), .A3(G104), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n336), .A2(G107), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n337), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT77), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT77), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n337), .A2(new_n340), .A3(new_n344), .A4(new_n341), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n343), .A2(G101), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G101), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n337), .A2(new_n340), .A3(new_n347), .A4(new_n341), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(KEYINPUT4), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n343), .A2(new_n350), .A3(G101), .A4(new_n345), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n351), .A2(new_n352), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n248), .B(new_n349), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n341), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n336), .A2(G107), .ZN(new_n357));
  OAI21_X1  g171(.A(G101), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n240), .A2(new_n243), .A3(KEYINPUT5), .A4(new_n241), .ZN(new_n359));
  OR3_X1    g173(.A1(new_n239), .A2(KEYINPUT5), .A3(G119), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(G113), .A3(new_n360), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n247), .A2(new_n348), .A3(new_n358), .A4(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n355), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(G110), .B(G122), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n365), .A2(KEYINPUT82), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n367), .B1(new_n355), .B2(new_n362), .ZN(new_n368));
  AOI22_X1  g182(.A1(new_n364), .A2(new_n365), .B1(new_n368), .B2(KEYINPUT6), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n368), .A2(KEYINPUT6), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n335), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT86), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n355), .A2(new_n362), .A3(new_n365), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n331), .A2(KEYINPUT7), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n327), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n322), .A2(new_n325), .A3(new_n326), .A4(new_n375), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n247), .A2(new_n361), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n358), .A2(new_n348), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n362), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n365), .B(KEYINPUT8), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n377), .A2(new_n378), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n374), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G902), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n373), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI211_X1 g201(.A(KEYINPUT86), .B(G902), .C1(new_n374), .C2(new_n384), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n321), .B1(new_n372), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(G902), .B1(new_n374), .B2(new_n384), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(new_n373), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n368), .A2(KEYINPUT6), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n374), .ZN(new_n394));
  OAI22_X1  g208(.A1(new_n394), .A2(new_n370), .B1(new_n333), .B2(new_n334), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n392), .A2(new_n395), .A3(new_n320), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n319), .B1(new_n390), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(G234), .A2(G237), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(G902), .A3(G953), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n399), .B(KEYINPUT96), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT21), .B(G898), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n398), .A2(G952), .A3(new_n329), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(G113), .B(G122), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT90), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n405), .B(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(new_n336), .ZN(new_n408));
  INV_X1    g222(.A(G140), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n324), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(G125), .A2(G140), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n201), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n410), .A2(G146), .A3(new_n411), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT87), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT87), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n413), .A2(new_n417), .A3(new_n414), .ZN(new_n418));
  INV_X1    g232(.A(G237), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(new_n329), .A3(G214), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n203), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n262), .A2(G143), .A3(G214), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT88), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT18), .ZN(new_n425));
  OAI22_X1  g239(.A1(new_n423), .A2(new_n424), .B1(new_n425), .B2(new_n195), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n425), .A2(new_n195), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n421), .A2(KEYINPUT88), .A3(new_n427), .A4(new_n422), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n416), .A2(new_n418), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n423), .A2(KEYINPUT17), .A3(G131), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n412), .A2(KEYINPUT16), .ZN(new_n432));
  NOR3_X1   g246(.A1(new_n324), .A2(KEYINPUT16), .A3(G140), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(G146), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT16), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n436), .B1(new_n410), .B2(new_n411), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n437), .A2(new_n201), .A3(new_n433), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT92), .ZN(new_n439));
  NOR3_X1   g253(.A1(new_n435), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n432), .A2(G146), .A3(new_n434), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n201), .B1(new_n437), .B2(new_n433), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT92), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n431), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n422), .ZN(new_n445));
  AOI21_X1  g259(.A(G143), .B1(new_n262), .B2(G214), .ZN(new_n446));
  OAI21_X1  g260(.A(G131), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT17), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n421), .A2(new_n195), .A3(new_n422), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT93), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n447), .A2(KEYINPUT93), .A3(new_n448), .A4(new_n449), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n408), .B(new_n430), .C1(new_n444), .C2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n416), .A2(new_n418), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n426), .A2(new_n428), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n437), .A2(new_n433), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n447), .A2(new_n449), .B1(new_n458), .B2(G146), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n412), .A2(KEYINPUT89), .A3(KEYINPUT19), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT19), .B1(new_n412), .B2(KEYINPUT89), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n201), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n456), .A2(new_n457), .B1(new_n459), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT91), .B1(new_n464), .B2(new_n408), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT91), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n407), .B(G104), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n459), .A2(new_n463), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n466), .B(new_n467), .C1(new_n468), .C2(new_n429), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n455), .A2(new_n465), .A3(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(G475), .A2(G902), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT20), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n455), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n439), .B1(new_n435), .B2(new_n438), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n441), .A2(new_n442), .A3(KEYINPUT92), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n478), .A2(new_n431), .A3(new_n452), .A4(new_n453), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n408), .B1(new_n479), .B2(new_n430), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n386), .B1(new_n475), .B2(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT94), .B(G475), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n470), .A2(KEYINPUT20), .A3(new_n471), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n474), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(G116), .B(G122), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n339), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n239), .A2(KEYINPUT14), .A3(G122), .ZN(new_n488));
  INV_X1    g302(.A(new_n486), .ZN(new_n489));
  OAI211_X1 g303(.A(G107), .B(new_n488), .C1(new_n489), .C2(KEYINPUT14), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n207), .A2(G143), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n203), .A2(G128), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT95), .ZN(new_n494));
  XNOR2_X1  g308(.A(G128), .B(G143), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT95), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n494), .A2(new_n497), .A3(new_n188), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n188), .B1(new_n494), .B2(new_n497), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n487), .B(new_n490), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n495), .A2(KEYINPUT13), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n501), .B(G134), .C1(KEYINPUT13), .C2(new_n492), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n486), .B(new_n339), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n494), .A2(new_n497), .A3(new_n188), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  XOR2_X1   g320(.A(KEYINPUT9), .B(G234), .Z(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(G217), .A3(new_n329), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n508), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n500), .A2(new_n505), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n386), .ZN(new_n513));
  INV_X1    g327(.A(G478), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(KEYINPUT15), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n512), .B(new_n386), .C1(KEYINPUT15), .C2(new_n514), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n485), .A2(new_n518), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n397), .A2(new_n404), .A3(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(G217), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n521), .B1(G234), .B2(new_n386), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n242), .A2(G128), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n524), .A2(KEYINPUT23), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(KEYINPUT23), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n525), .B(new_n526), .C1(G119), .C2(new_n207), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n527), .A2(G110), .ZN(new_n528));
  XNOR2_X1  g342(.A(G119), .B(G128), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(KEYINPUT74), .ZN(new_n530));
  XOR2_X1   g344(.A(KEYINPUT24), .B(G110), .Z(new_n531));
  NOR2_X1   g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n441), .B(new_n413), .C1(new_n528), .C2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n530), .A2(new_n531), .ZN(new_n534));
  XOR2_X1   g348(.A(new_n534), .B(KEYINPUT75), .Z(new_n535));
  NAND2_X1  g349(.A1(new_n527), .A2(G110), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n536), .B1(new_n435), .B2(new_n438), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n533), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n329), .A2(G221), .A3(G234), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT22), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(G137), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n533), .B(new_n541), .C1(new_n535), .C2(new_n537), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n386), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT25), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n543), .A2(KEYINPUT25), .A3(new_n386), .A4(new_n544), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n523), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n545), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n549), .B1(new_n523), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n507), .ZN(new_n552));
  OAI21_X1  g366(.A(G221), .B1(new_n552), .B2(G902), .ZN(new_n553));
  XNOR2_X1  g367(.A(G110), .B(G140), .ZN(new_n554));
  INV_X1    g368(.A(G227), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(G953), .ZN(new_n556));
  XOR2_X1   g370(.A(new_n554), .B(new_n556), .Z(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n210), .B(new_n349), .C1(new_n353), .C2(new_n354), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n199), .A2(new_n200), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n219), .A2(new_n380), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT10), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n561), .B(new_n562), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n559), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n560), .B1(new_n559), .B2(new_n563), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n558), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT81), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n559), .A2(new_n560), .A3(new_n563), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n557), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n219), .B(new_n380), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n278), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT79), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT12), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n380), .B(new_n225), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n575), .B1(new_n577), .B2(new_n560), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT79), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n572), .A2(KEYINPUT12), .A3(new_n197), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n571), .A2(new_n582), .ZN(new_n583));
  OAI211_X1 g397(.A(KEYINPUT81), .B(new_n558), .C1(new_n564), .C2(new_n565), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n568), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(G469), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n586), .A3(new_n386), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT80), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n570), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n565), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n569), .A2(KEYINPUT80), .A3(new_n557), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  XOR2_X1   g407(.A(new_n557), .B(KEYINPUT76), .Z(new_n594));
  INV_X1    g408(.A(new_n581), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n595), .B1(new_n576), .B2(new_n579), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n594), .B1(new_n596), .B2(new_n564), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n593), .A2(new_n597), .A3(G469), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n586), .A2(new_n386), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n553), .B1(new_n588), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n317), .A2(new_n520), .A3(new_n551), .A4(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  AND3_X1   g419(.A1(new_n474), .A2(new_n483), .A3(new_n484), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n512), .A2(KEYINPUT33), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT33), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n509), .A2(new_n608), .A3(new_n511), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(G478), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n512), .A2(new_n514), .A3(new_n386), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n514), .A2(new_n386), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n606), .A2(new_n614), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n397), .A2(new_n404), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT97), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n617), .B(G472), .C1(new_n313), .C2(G902), .ZN(new_n618));
  OAI21_X1  g432(.A(KEYINPUT97), .B1(new_n313), .B2(new_n314), .ZN(new_n619));
  INV_X1    g433(.A(G472), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n284), .B2(new_n386), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n618), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n616), .A2(new_n622), .A3(new_n603), .A4(new_n551), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT34), .B(G104), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G6));
  AND2_X1   g439(.A1(new_n397), .A2(new_n404), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n474), .A2(new_n483), .A3(new_n518), .A4(new_n484), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n629), .A2(new_n551), .A3(new_n603), .A4(new_n622), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT35), .B(G107), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT98), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n630), .B(new_n632), .ZN(G9));
  NOR2_X1   g447(.A1(new_n542), .A2(KEYINPUT36), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n538), .B(new_n634), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n635), .A2(new_n386), .A3(new_n523), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n549), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(KEYINPUT99), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT99), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n639), .B1(new_n549), .B2(new_n636), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n520), .A2(new_n622), .A3(new_n603), .A4(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT37), .ZN(new_n643));
  XOR2_X1   g457(.A(new_n643), .B(G110), .Z(G12));
  NAND2_X1  g458(.A1(new_n317), .A2(new_n641), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n390), .A2(new_n396), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n318), .ZN(new_n648));
  INV_X1    g462(.A(G900), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n400), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n403), .B(KEYINPUT100), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n606), .A2(KEYINPUT101), .A3(new_n518), .A4(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT101), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n655), .B1(new_n627), .B2(new_n652), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n602), .A2(new_n648), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n646), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G128), .ZN(G30));
  XOR2_X1   g474(.A(new_n652), .B(KEYINPUT39), .Z(new_n661));
  NAND2_X1  g475(.A1(new_n603), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(KEYINPUT40), .ZN(new_n663));
  AOI22_X1  g477(.A1(new_n273), .A2(new_n291), .B1(new_n269), .B2(new_n271), .ZN(new_n664));
  OAI21_X1  g478(.A(G472), .B1(new_n664), .B2(G902), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n288), .A2(new_n315), .A3(new_n316), .A4(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n663), .A2(new_n637), .A3(new_n666), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n485), .A2(new_n518), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n318), .B(new_n668), .C1(new_n662), .C2(KEYINPUT40), .ZN(new_n669));
  XOR2_X1   g483(.A(new_n647), .B(KEYINPUT38), .Z(new_n670));
  NOR3_X1   g484(.A1(new_n667), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(new_n203), .ZN(G45));
  INV_X1    g486(.A(new_n614), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n485), .A2(new_n673), .A3(new_n653), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n675), .B(new_n553), .C1(new_n588), .C2(new_n601), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n648), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n646), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G146), .ZN(G48));
  AND2_X1   g493(.A1(new_n317), .A2(new_n551), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n585), .A2(new_n386), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(G469), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n682), .A2(new_n553), .A3(new_n587), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT102), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT102), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n682), .A2(new_n685), .A3(new_n553), .A4(new_n587), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n680), .A2(new_n616), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT41), .B(G113), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G15));
  NAND4_X1  g504(.A1(new_n317), .A2(new_n551), .A3(new_n684), .A4(new_n686), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n626), .A2(new_n628), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n239), .ZN(G18));
  NAND3_X1  g508(.A1(new_n646), .A2(new_n520), .A3(new_n687), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G119), .ZN(G21));
  INV_X1    g510(.A(new_n272), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n266), .B1(new_n292), .B2(new_n304), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n697), .B1(new_n698), .B2(KEYINPUT103), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT103), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n700), .B(new_n266), .C1(new_n292), .C2(new_n304), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n314), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT104), .B(G472), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n705), .B1(new_n284), .B2(new_n386), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n626), .A2(new_n703), .A3(new_n551), .A4(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n684), .A2(new_n668), .A3(new_n686), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  NOR4_X1   g525(.A1(new_n702), .A2(new_n706), .A3(new_n637), .A4(new_n674), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n712), .A2(new_n397), .A3(new_n686), .A4(new_n684), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G125), .ZN(G27));
  NOR2_X1   g528(.A1(new_n647), .A2(new_n319), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n676), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n315), .A2(new_n308), .A3(new_n286), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n718), .A2(KEYINPUT105), .A3(new_n551), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT105), .B1(new_n718), .B2(new_n551), .ZN(new_n720));
  OAI211_X1 g534(.A(KEYINPUT42), .B(new_n717), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n676), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n317), .A2(new_n722), .A3(new_n551), .A4(new_n715), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT42), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G131), .ZN(G33));
  AND3_X1   g541(.A1(new_n317), .A2(new_n551), .A3(new_n715), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n728), .A2(new_n603), .A3(new_n656), .A4(new_n654), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G134), .ZN(G36));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n598), .B1(new_n731), .B2(new_n586), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT106), .ZN(new_n733));
  OR2_X1    g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n593), .A2(KEYINPUT45), .A3(new_n597), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n732), .A2(new_n733), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n600), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT46), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n737), .A2(KEYINPUT46), .A3(new_n600), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n740), .A2(new_n587), .A3(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n553), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n622), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n485), .A2(new_n614), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT43), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n745), .B(new_n747), .C1(new_n549), .C2(new_n636), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n716), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n748), .A2(new_n749), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n744), .A2(new_n661), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G137), .ZN(G39));
  INV_X1    g567(.A(KEYINPUT47), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n754), .B1(new_n742), .B2(new_n743), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n740), .A2(new_n587), .A3(new_n741), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(KEYINPUT47), .A3(new_n553), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n317), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n551), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n758), .A2(new_n759), .A3(new_n675), .A4(new_n715), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G140), .ZN(G42));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n317), .B(new_n641), .C1(new_n658), .C2(new_n677), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n397), .A2(new_n653), .A3(new_n668), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n666), .A2(new_n764), .A3(new_n603), .A4(new_n637), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(new_n713), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n763), .A2(new_n713), .A3(KEYINPUT52), .A4(new_n765), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT109), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n604), .A2(new_n623), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT108), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT108), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n604), .A2(new_n623), .A3(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n773), .A2(new_n630), .A3(new_n642), .A4(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n680), .A2(new_n629), .A3(new_n687), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n695), .A2(new_n710), .A3(new_n688), .A4(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n702), .A2(new_n637), .A3(new_n706), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n675), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n519), .A2(new_n653), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n781), .B1(new_n645), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n603), .A3(new_n715), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n726), .A2(new_n729), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n771), .B1(new_n779), .B2(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n775), .A2(new_n630), .ZN(new_n787));
  INV_X1    g601(.A(new_n616), .ZN(new_n788));
  OAI22_X1  g602(.A1(new_n691), .A2(new_n788), .B1(new_n708), .B2(new_n709), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n693), .ZN(new_n790));
  INV_X1    g604(.A(new_n642), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n791), .B1(new_n772), .B2(KEYINPUT108), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n787), .A2(new_n790), .A3(new_n695), .A4(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n726), .A2(new_n784), .A3(new_n729), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n793), .A2(KEYINPUT109), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n770), .B1(new_n786), .B2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n793), .A2(new_n797), .A3(new_n794), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n768), .A2(KEYINPUT110), .A3(new_n769), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT110), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n766), .A2(new_n801), .A3(new_n767), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT112), .B1(new_n799), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n775), .A2(new_n630), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n774), .B1(new_n604), .B2(new_n623), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n805), .A2(new_n791), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n778), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n785), .A2(new_n807), .A3(KEYINPUT53), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n800), .A2(new_n802), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT112), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n804), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n798), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n796), .A2(KEYINPUT53), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n779), .A2(new_n771), .A3(new_n785), .ZN(new_n817));
  OAI21_X1  g631(.A(KEYINPUT109), .B1(new_n793), .B2(new_n794), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT53), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n803), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n816), .A2(KEYINPUT54), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n762), .B1(new_n815), .B2(new_n821), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n796), .A2(KEYINPUT53), .B1(new_n819), .B2(new_n803), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT111), .B1(new_n823), .B2(KEYINPUT54), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n687), .A2(new_n715), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT114), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT114), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n687), .A2(new_n827), .A3(new_n715), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n747), .A2(new_n651), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n719), .A2(new_n720), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OR2_X1    g647(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n834));
  NAND2_X1  g648(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n831), .A2(KEYINPUT117), .A3(KEYINPUT48), .A4(new_n832), .ZN(new_n837));
  AND4_X1   g651(.A1(new_n551), .A2(new_n830), .A3(new_n703), .A4(new_n707), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n397), .A3(new_n687), .ZN(new_n839));
  INV_X1    g653(.A(G952), .ZN(new_n840));
  OR3_X1    g654(.A1(new_n840), .A2(KEYINPUT116), .A3(G953), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT116), .B1(new_n840), .B2(G953), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n837), .A2(new_n839), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n403), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n666), .A2(new_n759), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n829), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT115), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n829), .A2(KEYINPUT115), .A3(new_n844), .A4(new_n845), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n843), .B1(new_n615), .B2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n848), .A2(new_n606), .A3(new_n614), .A4(new_n849), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n682), .A2(new_n587), .ZN(new_n853));
  XOR2_X1   g667(.A(new_n853), .B(KEYINPUT107), .Z(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n743), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n755), .A2(new_n757), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(new_n715), .A3(new_n838), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n670), .A2(new_n319), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n838), .A2(new_n687), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT50), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n838), .A2(KEYINPUT50), .A3(new_n687), .A4(new_n858), .ZN(new_n862));
  AOI22_X1  g676(.A1(new_n831), .A2(new_n780), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n852), .A2(new_n857), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT113), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n864), .A2(new_n865), .A3(KEYINPUT51), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT51), .B1(new_n864), .B2(new_n865), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n836), .B(new_n851), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n822), .A2(new_n824), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(G952), .A2(G953), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n746), .A2(new_n553), .A3(new_n318), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n854), .B(KEYINPUT49), .ZN(new_n872));
  INV_X1    g686(.A(new_n666), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n872), .A2(new_n551), .A3(new_n670), .A4(new_n873), .ZN(new_n874));
  OAI22_X1  g688(.A1(new_n869), .A2(new_n870), .B1(new_n871), .B2(new_n874), .ZN(G75));
  NOR2_X1   g689(.A1(new_n394), .A2(new_n370), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n335), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n395), .ZN(new_n878));
  XNOR2_X1  g692(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n878), .B(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n386), .B1(new_n798), .B2(new_n813), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(G210), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT56), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI211_X1 g699(.A(KEYINPUT56), .B(new_n880), .C1(new_n882), .C2(G210), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n329), .A2(G952), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(G51));
  OR2_X1    g702(.A1(new_n600), .A2(KEYINPUT57), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n600), .A2(KEYINPUT57), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n814), .B1(new_n798), .B2(new_n813), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n817), .A2(new_n818), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT53), .B1(new_n892), .B2(new_n770), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n799), .A2(new_n803), .A3(KEYINPUT112), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n811), .B1(new_n809), .B2(new_n810), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n893), .A2(new_n896), .A3(KEYINPUT54), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n889), .B(new_n890), .C1(new_n891), .C2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n585), .ZN(new_n899));
  INV_X1    g713(.A(new_n737), .ZN(new_n900));
  OAI211_X1 g714(.A(G902), .B(new_n900), .C1(new_n893), .C2(new_n896), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT119), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n901), .B(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n887), .B1(new_n899), .B2(new_n903), .ZN(G54));
  NAND3_X1  g718(.A1(new_n882), .A2(KEYINPUT58), .A3(G475), .ZN(new_n905));
  INV_X1    g719(.A(new_n470), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n905), .A2(new_n906), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n907), .A2(new_n908), .A3(new_n887), .ZN(G60));
  AND2_X1   g723(.A1(new_n607), .A2(new_n609), .ZN(new_n910));
  XNOR2_X1  g724(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n613), .B(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n913), .B1(new_n891), .B2(new_n897), .ZN(new_n914));
  INV_X1    g728(.A(new_n887), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n912), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n917), .B1(new_n822), .B2(new_n824), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n916), .B1(new_n918), .B2(new_n910), .ZN(G63));
  NAND2_X1  g733(.A1(G217), .A2(G902), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT60), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n635), .B(KEYINPUT121), .Z(new_n923));
  OAI211_X1 g737(.A(new_n922), .B(new_n923), .C1(new_n893), .C2(new_n896), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n921), .B1(new_n798), .B2(new_n813), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n543), .A2(new_n544), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n915), .B(new_n924), .C1(new_n925), .C2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT61), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n928), .A2(KEYINPUT122), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(KEYINPUT122), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n927), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n922), .B1(new_n893), .B2(new_n896), .ZN(new_n932));
  INV_X1    g746(.A(new_n926), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n887), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n934), .A2(KEYINPUT122), .A3(new_n928), .A4(new_n924), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n931), .A2(new_n935), .ZN(G66));
  INV_X1    g750(.A(G224), .ZN(new_n937));
  OAI21_X1  g751(.A(G953), .B1(new_n401), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n938), .B1(new_n779), .B2(G953), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n876), .B1(G898), .B2(new_n329), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT123), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n939), .B(new_n941), .ZN(G69));
  NAND2_X1  g756(.A1(G900), .A2(G953), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n397), .A2(new_n668), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n744), .A2(new_n661), .A3(new_n832), .A4(new_n944), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n752), .A2(new_n945), .A3(new_n729), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n763), .A2(new_n713), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n946), .A2(new_n760), .A3(new_n726), .A4(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n943), .B1(new_n949), .B2(G953), .ZN(new_n950));
  INV_X1    g764(.A(new_n255), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n229), .B1(KEYINPUT30), .B2(new_n951), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT124), .Z(new_n953));
  OR2_X1    g767(.A1(new_n461), .A2(new_n462), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n953), .B(new_n954), .Z(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n950), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n671), .A2(new_n947), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT62), .ZN(new_n959));
  INV_X1    g773(.A(new_n662), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n728), .B(new_n960), .C1(new_n615), .C2(new_n628), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT125), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n752), .A2(new_n962), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n963), .A2(KEYINPUT126), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n963), .A2(KEYINPUT126), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n760), .B(new_n959), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n955), .B1(new_n966), .B2(new_n329), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(G953), .B1(new_n555), .B2(new_n649), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(KEYINPUT127), .ZN(new_n970));
  OR2_X1    g784(.A1(new_n969), .A2(KEYINPUT127), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n957), .A2(new_n968), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n950), .A2(new_n956), .ZN(new_n973));
  OAI211_X1 g787(.A(KEYINPUT127), .B(new_n969), .C1(new_n973), .C2(new_n967), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n972), .A2(new_n974), .ZN(G72));
  NAND2_X1  g789(.A1(G472), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT63), .Z(new_n977));
  OAI21_X1  g791(.A(new_n977), .B1(new_n966), .B2(new_n793), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n978), .A2(new_n264), .A3(new_n297), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n298), .A2(new_n282), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n823), .A2(new_n977), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n977), .B1(new_n949), .B2(new_n793), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n982), .A2(new_n259), .A3(new_n293), .A4(new_n271), .ZN(new_n983));
  AND4_X1   g797(.A1(new_n915), .A2(new_n979), .A3(new_n981), .A4(new_n983), .ZN(G57));
endmodule


