//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n558, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n612, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1161;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT66), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT67), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT68), .B(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G238), .A3(G237), .A4(G235), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT70), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT71), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OR2_X1    g036(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT72), .B(G2105), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(new_n469), .A3(G137), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n468), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n471));
  OAI211_X1 g046(.A(new_n467), .B(new_n470), .C1(new_n471), .C2(new_n469), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  OAI221_X1 g048(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n469), .C2(G112), .ZN(new_n474));
  INV_X1    g049(.A(G124), .ZN(new_n475));
  INV_X1    g050(.A(new_n469), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n468), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n474), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT73), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n479), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G2105), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n468), .A2(KEYINPUT73), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n478), .B1(G136), .B2(new_n487), .ZN(G162));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT74), .ZN(new_n491));
  OAI21_X1  g066(.A(G2105), .B1(new_n491), .B2(G114), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(KEYINPUT74), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n490), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n480), .A2(new_n482), .A3(G126), .A4(G2105), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n485), .A2(KEYINPUT72), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT72), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n480), .A2(new_n482), .A3(new_n498), .A4(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G138), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT4), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n468), .A2(new_n469), .A3(new_n504), .A4(G138), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n497), .B1(new_n503), .B2(new_n505), .ZN(G164));
  XNOR2_X1  g081(.A(KEYINPUT5), .B(G543), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT75), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  XOR2_X1   g085(.A(KEYINPUT6), .B(G651), .Z(new_n511));
  AOI22_X1  g086(.A1(new_n507), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR3_X1   g088(.A1(new_n508), .A2(KEYINPUT75), .A3(new_n509), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(G166));
  INV_X1    g090(.A(G51), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT77), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OR2_X1    g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(KEYINPUT77), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT78), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n520), .A2(KEYINPUT78), .A3(new_n523), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n516), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  XOR2_X1   g103(.A(KEYINPUT5), .B(G543), .Z(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n511), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G89), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n529), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n507), .A2(KEYINPUT76), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(G63), .A2(G651), .ZN(new_n538));
  OAI211_X1 g113(.A(new_n531), .B(new_n533), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n528), .A2(new_n539), .ZN(G168));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G64), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  XNOR2_X1  g118(.A(KEYINPUT79), .B(G90), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n543), .A2(G651), .B1(new_n530), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n526), .A2(new_n527), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G52), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n545), .A2(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n537), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n552), .A2(G651), .B1(G81), .B2(new_n530), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n546), .A2(G43), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n529), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n565), .A2(G651), .B1(new_n530), .B2(G91), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n520), .A2(KEYINPUT9), .A3(G53), .A4(new_n523), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n520), .A2(G53), .A3(new_n523), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n566), .A2(new_n567), .A3(new_n570), .ZN(G299));
  INV_X1    g146(.A(G168), .ZN(G286));
  OR2_X1    g147(.A1(new_n513), .A2(new_n514), .ZN(G303));
  NAND3_X1  g148(.A1(new_n520), .A2(G49), .A3(new_n523), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n530), .A2(G87), .ZN(new_n575));
  AOI21_X1  g150(.A(G74), .B1(new_n535), .B2(new_n536), .ZN(new_n576));
  OAI211_X1 g151(.A(new_n574), .B(new_n575), .C1(new_n576), .C2(new_n509), .ZN(G288));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  XOR2_X1   g153(.A(new_n578), .B(KEYINPUT81), .Z(new_n579));
  INV_X1    g154(.A(KEYINPUT80), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n507), .A2(new_n580), .A3(G61), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n580), .B1(new_n507), .B2(G61), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n507), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n585), .A2(new_n511), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT82), .ZN(G305));
  NAND2_X1  g163(.A1(G72), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G60), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n537), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(G85), .B2(new_n530), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n546), .A2(G47), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(new_n530), .A2(G92), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n530), .A2(KEYINPUT10), .A3(G92), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  XNOR2_X1  g174(.A(KEYINPUT83), .B(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n529), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n597), .A2(new_n598), .B1(G651), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n546), .A2(G54), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G171), .B2(new_n605), .ZN(G284));
  XNOR2_X1  g182(.A(G284), .B(KEYINPUT84), .ZN(G321));
  NAND2_X1  g183(.A1(G299), .A2(new_n605), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G168), .B2(new_n605), .ZN(G297));
  OAI21_X1  g185(.A(new_n609), .B1(G168), .B2(new_n605), .ZN(G280));
  INV_X1    g186(.A(new_n604), .ZN(new_n612));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n555), .A2(new_n605), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n604), .A2(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(new_n605), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g193(.A1(new_n485), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2100), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n487), .A2(G135), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT85), .ZN(new_n624));
  INV_X1    g199(.A(new_n477), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n469), .A2(G111), .ZN(new_n626));
  OAI21_X1  g201(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  AOI22_X1  g203(.A1(new_n625), .A2(G123), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(G2096), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n622), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n633), .B1(new_n632), .B2(new_n631), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT86), .ZN(G156));
  INV_X1    g210(.A(KEYINPUT14), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2427), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n636), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(new_n639), .B2(new_n638), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n641), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  AND3_X1   g224(.A1(new_n648), .A2(G14), .A3(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT87), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT88), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n652), .A2(new_n654), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(new_n657), .A3(KEYINPUT17), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT18), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g235(.A1(G2072), .A2(G2078), .ZN(new_n661));
  OAI22_X1  g236(.A1(new_n655), .A2(new_n659), .B1(new_n442), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n660), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2096), .B(G2100), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1956), .B(G2474), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT20), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n668), .A2(new_n669), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n667), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n667), .B2(new_n673), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1991), .B(G1996), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G229));
  INV_X1    g257(.A(G16), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G22), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(G166), .B2(new_n683), .ZN(new_n685));
  INV_X1    g260(.A(G1971), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n683), .A2(G23), .ZN(new_n688));
  INV_X1    g263(.A(G288), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n688), .B1(new_n689), .B2(new_n683), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT33), .B(G1976), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n687), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT32), .B(G1981), .Z(new_n694));
  OR2_X1    g269(.A1(G6), .A2(G16), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G305), .B2(new_n683), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n693), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(new_n694), .B2(new_n696), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n698), .A2(KEYINPUT34), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(KEYINPUT34), .ZN(new_n700));
  INV_X1    g275(.A(G25), .ZN(new_n701));
  OR3_X1    g276(.A1(new_n701), .A2(KEYINPUT89), .A3(G29), .ZN(new_n702));
  OAI21_X1  g277(.A(KEYINPUT89), .B1(new_n701), .B2(G29), .ZN(new_n703));
  OAI221_X1 g278(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n469), .C2(G107), .ZN(new_n704));
  INV_X1    g279(.A(G119), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(new_n705), .B2(new_n477), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G131), .B2(new_n487), .ZN(new_n707));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n702), .B(new_n703), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT35), .B(G1991), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(G16), .A2(G24), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G290), .B2(new_n683), .ZN(new_n713));
  INV_X1    g288(.A(G1986), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n711), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n714), .B2(new_n713), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n699), .A2(new_n700), .A3(new_n716), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT36), .Z(new_n718));
  NAND3_X1  g293(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT25), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G139), .B2(new_n487), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT92), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n723), .A2(new_n469), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  MUX2_X1   g300(.A(G33), .B(new_n725), .S(G29), .Z(new_n726));
  NOR2_X1   g301(.A1(new_n726), .A2(G2072), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT93), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n683), .A2(G20), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT23), .ZN(new_n730));
  INV_X1    g305(.A(G299), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(new_n683), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G1956), .ZN(new_n733));
  NAND2_X1  g308(.A1(G168), .A2(G16), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT96), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n734), .B(new_n735), .C1(G16), .C2(G21), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n735), .B2(new_n734), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1966), .ZN(new_n738));
  AOI211_X1 g313(.A(new_n733), .B(new_n738), .C1(G2072), .C2(new_n726), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n487), .A2(G141), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT95), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n625), .A2(G129), .ZN(new_n742));
  NAND3_X1  g317(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT26), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n745), .A2(new_n746), .B1(G105), .B2(new_n466), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n742), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n741), .A2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(new_n708), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n708), .B2(G32), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT27), .B(G1996), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n683), .A2(G4), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n612), .B2(new_n683), .ZN(new_n755));
  OAI22_X1  g330(.A1(new_n752), .A2(new_n753), .B1(G1348), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n683), .A2(G19), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n556), .B2(new_n683), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n756), .B1(G1341), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(G171), .A2(new_n683), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G5), .B2(new_n683), .ZN(new_n761));
  INV_X1    g336(.A(G1961), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n752), .A2(new_n753), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n755), .A2(G1348), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n761), .A2(new_n762), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n763), .A2(new_n764), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n708), .A2(G26), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n487), .A2(G140), .ZN(new_n771));
  OAI21_X1  g346(.A(G2104), .B1(new_n469), .B2(G116), .ZN(new_n772));
  NOR2_X1   g347(.A1(G104), .A2(G2105), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT90), .Z(new_n774));
  INV_X1    g349(.A(G128), .ZN(new_n775));
  OAI22_X1  g350(.A1(new_n772), .A2(new_n774), .B1(new_n477), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n771), .A2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n770), .B1(new_n778), .B2(G29), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G2067), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n708), .A2(G35), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G162), .B2(new_n708), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT29), .B(G2090), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT31), .B(G11), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT97), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT30), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n787), .A2(G28), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n708), .B1(new_n787), .B2(G28), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT24), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n708), .B1(new_n790), .B2(G34), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n791), .A2(KEYINPUT94), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n790), .A2(G34), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n791), .B2(KEYINPUT94), .ZN(new_n794));
  OAI22_X1  g369(.A1(new_n472), .A2(new_n708), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(G2084), .ZN(new_n796));
  OAI221_X1 g371(.A(new_n786), .B1(new_n788), .B2(new_n789), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n796), .B2(new_n795), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n780), .A2(new_n784), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(G27), .A2(G29), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G164), .B2(G29), .ZN(new_n801));
  INV_X1    g376(.A(G2078), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  OAI221_X1 g378(.A(new_n803), .B1(new_n708), .B2(new_n630), .C1(new_n758), .C2(G1341), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n767), .A2(new_n799), .A3(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n728), .A2(new_n739), .A3(new_n759), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n718), .A2(new_n806), .ZN(G311));
  OR2_X1    g382(.A1(new_n718), .A2(new_n806), .ZN(G150));
  NAND2_X1  g383(.A1(G80), .A2(G543), .ZN(new_n809));
  INV_X1    g384(.A(G67), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n537), .B2(new_n810), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n811), .A2(G651), .B1(G93), .B2(new_n530), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n546), .A2(G55), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G860), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT37), .Z(new_n816));
  NOR2_X1   g391(.A1(new_n604), .A2(new_n613), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT98), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT38), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n555), .A2(new_n814), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n553), .A2(new_n812), .A3(new_n554), .A4(new_n813), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n819), .B(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n824), .A2(KEYINPUT39), .ZN(new_n825));
  INV_X1    g400(.A(G860), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n824), .B2(KEYINPUT39), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n816), .B1(new_n825), .B2(new_n827), .ZN(G145));
  NAND2_X1  g403(.A1(new_n750), .A2(G164), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n503), .A2(new_n505), .ZN(new_n830));
  INV_X1    g405(.A(new_n497), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n749), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(new_n777), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n829), .A2(new_n778), .A3(new_n833), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT100), .ZN(new_n838));
  OAI21_X1  g413(.A(KEYINPUT99), .B1(new_n725), .B2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT99), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n722), .A2(new_n840), .A3(KEYINPUT100), .A4(new_n724), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n837), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n835), .A2(new_n839), .A3(new_n841), .A4(new_n836), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI221_X1 g420(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n469), .C2(G118), .ZN(new_n846));
  INV_X1    g421(.A(G130), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n846), .B1(new_n847), .B2(new_n477), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(G142), .B2(new_n487), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n620), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(new_n707), .Z(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n845), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n843), .A2(new_n844), .A3(new_n851), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(G162), .B(new_n472), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n631), .ZN(new_n857));
  AOI21_X1  g432(.A(G37), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n851), .B1(new_n845), .B2(KEYINPUT101), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT102), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT101), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n843), .A2(new_n861), .A3(new_n844), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n857), .ZN(new_n864));
  AND2_X1   g439(.A1(new_n854), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n860), .B1(new_n859), .B2(new_n862), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n858), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g444(.A(new_n822), .B(KEYINPUT103), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(new_n616), .Z(new_n871));
  AOI21_X1  g446(.A(G299), .B1(new_n602), .B2(new_n603), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n602), .A2(new_n603), .A3(G299), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n873), .A2(KEYINPUT41), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT104), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n874), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n878), .A2(new_n872), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n879), .A2(KEYINPUT104), .A3(KEYINPUT41), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT41), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(new_n878), .B2(new_n872), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n877), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n871), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(KEYINPUT105), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT105), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n871), .A2(new_n886), .A3(new_n883), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n871), .A2(new_n879), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n885), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(G305), .B(G288), .ZN(new_n890));
  XNOR2_X1  g465(.A(G290), .B(G303), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n890), .B(new_n891), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n892), .B(KEYINPUT42), .Z(new_n893));
  AND2_X1   g468(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n889), .A2(new_n893), .ZN(new_n895));
  OAI21_X1  g470(.A(G868), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n814), .A2(new_n605), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(G295));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n897), .ZN(G331));
  NAND3_X1  g474(.A1(new_n820), .A2(G301), .A3(new_n821), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(G301), .B1(new_n820), .B2(new_n821), .ZN(new_n902));
  OAI21_X1  g477(.A(G286), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n902), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(G168), .A3(new_n900), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n883), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(KEYINPUT106), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT106), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n883), .A2(new_n903), .A3(new_n905), .A4(new_n908), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n901), .A2(G286), .A3(new_n902), .ZN(new_n910));
  AOI21_X1  g485(.A(G168), .B1(new_n904), .B2(new_n900), .ZN(new_n911));
  OAI22_X1  g486(.A1(new_n910), .A2(new_n911), .B1(new_n872), .B2(new_n878), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n907), .A2(new_n892), .A3(new_n909), .A4(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(G37), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n918));
  INV_X1    g493(.A(new_n892), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n903), .A2(new_n905), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n920), .B1(new_n875), .B2(new_n882), .ZN(new_n921));
  INV_X1    g496(.A(new_n912), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n919), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n916), .A2(new_n917), .A3(new_n918), .A4(new_n923), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n923), .A2(new_n913), .A3(new_n918), .A4(new_n914), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT107), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n912), .A2(new_n909), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n892), .B1(new_n927), .B2(new_n907), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT43), .B1(new_n928), .B2(new_n915), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n924), .A2(new_n926), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n927), .A2(new_n907), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n919), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n916), .A2(new_n934), .A3(new_n918), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n916), .A2(new_n934), .A3(KEYINPUT108), .A4(new_n918), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n923), .A2(new_n913), .A3(new_n914), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n931), .B1(new_n939), .B2(KEYINPUT43), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n937), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n932), .A2(new_n941), .ZN(G397));
  INV_X1    g517(.A(KEYINPUT120), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n944));
  INV_X1    g519(.A(G40), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT110), .B1(new_n472), .B2(new_n945), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n468), .A2(G125), .ZN(new_n947));
  AND2_X1   g522(.A1(G113), .A2(G2104), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n476), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n470), .A2(new_n467), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT110), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n949), .A2(new_n950), .A3(new_n951), .A4(G40), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n944), .A2(new_n946), .A3(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G2090), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT50), .ZN(new_n955));
  INV_X1    g530(.A(G1384), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n832), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n953), .A2(KEYINPUT111), .A3(new_n954), .A4(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT111), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n957), .A2(new_n944), .A3(new_n946), .A4(new_n952), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n959), .B1(new_n960), .B2(G2090), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n832), .A2(KEYINPUT45), .A3(new_n956), .ZN(new_n962));
  XNOR2_X1  g537(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n963), .B1(G164), .B2(G1384), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n962), .A2(new_n964), .A3(new_n946), .A4(new_n952), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n686), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n958), .A2(new_n961), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT112), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT112), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n958), .A2(new_n961), .A3(new_n969), .A4(new_n966), .ZN(new_n970));
  XNOR2_X1  g545(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n971));
  NAND3_X1  g546(.A1(G303), .A2(G8), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT114), .ZN(new_n973));
  INV_X1    g548(.A(new_n971), .ZN(new_n974));
  INV_X1    g549(.A(G8), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n974), .B1(G166), .B2(new_n975), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n972), .A2(new_n973), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n973), .B1(new_n972), .B2(new_n976), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n968), .A2(G8), .A3(new_n970), .A4(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n946), .A2(new_n952), .A3(new_n956), .A4(new_n832), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(new_n975), .ZN(new_n984));
  INV_X1    g559(.A(G1981), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n584), .A2(new_n985), .A3(new_n586), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT49), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n985), .B1(new_n584), .B2(new_n586), .ZN(new_n989));
  OR3_X1    g564(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n988), .B1(new_n987), .B2(new_n989), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n984), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n689), .A2(G1976), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n993), .A2(new_n982), .A3(G8), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT52), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT116), .ZN(new_n997));
  INV_X1    g572(.A(G1976), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT52), .B1(G288), .B2(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n999), .B(KEYINPUT115), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n997), .B1(new_n1000), .B2(new_n994), .ZN(new_n1001));
  XOR2_X1   g576(.A(new_n999), .B(KEYINPUT115), .Z(new_n1002));
  INV_X1    g577(.A(new_n994), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(KEYINPUT116), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n996), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n981), .A2(new_n1005), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n992), .A2(new_n998), .A3(new_n689), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n986), .B(KEYINPUT117), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n984), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n980), .A2(new_n1005), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n946), .A2(new_n952), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1013), .A2(new_n954), .A3(new_n957), .A4(new_n944), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n966), .A2(new_n1014), .A3(KEYINPUT118), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT118), .B1(new_n966), .B2(new_n1014), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n1015), .A2(new_n1016), .A3(new_n975), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n972), .A2(new_n976), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT119), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1016), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n966), .A2(new_n1014), .A3(KEYINPUT118), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(G8), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT119), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1023), .A2(new_n1024), .A3(new_n1018), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1012), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1966), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT45), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(G164), .B2(G1384), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1029), .A2(new_n946), .A3(new_n952), .ZN(new_n1030));
  NOR3_X1   g605(.A1(G164), .A2(G1384), .A3(new_n963), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1027), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1013), .A2(new_n796), .A3(new_n957), .A4(new_n944), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(G8), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1035), .A2(G286), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT63), .B1(new_n1026), .B2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n960), .A2(G2090), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1038), .A2(KEYINPUT111), .B1(new_n686), .B2(new_n965), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n969), .B1(new_n1039), .B2(new_n961), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n970), .A2(G8), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1018), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT63), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1035), .A2(new_n1043), .A3(G286), .ZN(new_n1044));
  AND4_X1   g619(.A1(new_n980), .A2(new_n1042), .A3(new_n1005), .A4(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n943), .B(new_n1011), .C1(new_n1037), .C2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1020), .A2(new_n1025), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n980), .A2(new_n1005), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1047), .A2(new_n1048), .A3(new_n1036), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1045), .B1(new_n1049), .B2(new_n1043), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT120), .B1(new_n1050), .B2(new_n1010), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT122), .ZN(new_n1052));
  AND3_X1   g627(.A1(G299), .A2(new_n1052), .A3(KEYINPUT57), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT57), .B1(G299), .B2(new_n1052), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g630(.A(KEYINPUT56), .B(G2072), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1013), .A2(new_n964), .A3(new_n962), .A4(new_n1056), .ZN(new_n1057));
  XOR2_X1   g632(.A(KEYINPUT121), .B(G1956), .Z(new_n1058));
  NAND2_X1  g633(.A1(new_n960), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1055), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1055), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1061));
  OR2_X1    g636(.A1(new_n982), .A2(G2067), .ZN(new_n1062));
  INV_X1    g637(.A(G1348), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n960), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n604), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1060), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT61), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1061), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1067), .B1(new_n1068), .B2(new_n1060), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1059), .A2(new_n1057), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1071), .A2(KEYINPUT61), .A3(new_n1061), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1062), .A2(new_n1064), .A3(new_n604), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT60), .B1(new_n1073), .B2(new_n1065), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1069), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g650(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT58), .B(G1341), .ZN(new_n1078));
  OAI22_X1  g653(.A1(new_n983), .A2(new_n1078), .B1(new_n965), .B2(G1996), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1077), .B1(new_n1080), .B2(new_n555), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1079), .A2(new_n556), .A3(new_n1076), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n604), .A2(KEYINPUT60), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1062), .A2(new_n1064), .A3(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1081), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1066), .B1(new_n1075), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT124), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g663(.A(KEYINPUT124), .B(new_n1066), .C1(new_n1075), .C2(new_n1085), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n962), .A2(new_n964), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1093), .A2(new_n802), .A3(new_n1013), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT127), .B(KEYINPUT53), .Z(new_n1095));
  AOI22_X1  g670(.A1(new_n1094), .A2(new_n1095), .B1(new_n762), .B2(new_n960), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1097), .A2(KEYINPUT53), .A3(new_n802), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(G301), .B(KEYINPUT54), .ZN(new_n1100));
  AND4_X1   g675(.A1(KEYINPUT53), .A2(G160), .A3(G40), .A4(new_n802), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1100), .B1(new_n1093), .B2(new_n1101), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1099), .A2(new_n1100), .B1(new_n1102), .B2(new_n1096), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n975), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1104));
  NOR2_X1   g679(.A1(G168), .A2(new_n975), .ZN(new_n1105));
  NOR3_X1   g680(.A1(new_n1104), .A2(KEYINPUT51), .A3(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(G286), .A2(KEYINPUT125), .A3(G8), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT125), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(G168), .B2(new_n975), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT51), .B1(new_n1104), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(KEYINPUT126), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT126), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1113), .B(KEYINPUT51), .C1(new_n1104), .C2(new_n1110), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1106), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1034), .A2(new_n1105), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1103), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1091), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1106), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1035), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1113), .B1(new_n1122), .B2(KEYINPUT51), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1114), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1120), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1125), .A2(KEYINPUT62), .A3(new_n1116), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT62), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(G301), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1047), .A2(new_n1048), .A3(new_n1130), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1090), .A2(new_n1119), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1046), .A2(new_n1051), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n946), .A2(new_n952), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1134), .A2(new_n964), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n777), .B(G2067), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n750), .A2(G1996), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n750), .A2(G1996), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1136), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n707), .A2(new_n710), .ZN(new_n1141));
  OR2_X1    g716(.A1(new_n707), .A2(new_n710), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g718(.A(G290), .B(G1986), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1135), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1133), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1136), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1135), .B1(new_n1147), .B2(new_n749), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n1134), .A2(G1996), .A3(new_n964), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1148), .B1(KEYINPUT46), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1150), .B1(KEYINPUT46), .B2(new_n1149), .ZN(new_n1151));
  XOR2_X1   g726(.A(new_n1151), .B(KEYINPUT47), .Z(new_n1152));
  NAND2_X1  g727(.A1(new_n1143), .A2(new_n1135), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1135), .A2(new_n714), .A3(new_n593), .A4(new_n592), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT48), .ZN(new_n1155));
  OAI22_X1  g730(.A1(new_n1139), .A2(new_n1141), .B1(G2067), .B2(new_n778), .ZN(new_n1156));
  AOI22_X1  g731(.A1(new_n1153), .A2(new_n1155), .B1(new_n1135), .B2(new_n1156), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1152), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1146), .A2(new_n1158), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g734(.A1(G229), .A2(new_n463), .A3(G401), .A4(G227), .ZN(new_n1161));
  NAND3_X1  g735(.A1(new_n930), .A2(new_n868), .A3(new_n1161), .ZN(G225));
  INV_X1    g736(.A(G225), .ZN(G308));
endmodule


