//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 0 0 1 0 1 0 1 1 1 1 1 1 0 0 0 0 0 1 0 1 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  OR2_X1    g001(.A1(KEYINPUT69), .A2(G116), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT69), .A2(G116), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(G119), .A3(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT68), .B1(new_n191), .B2(G119), .ZN(new_n192));
  OR3_X1    g006(.A1(new_n191), .A2(KEYINPUT68), .A3(G119), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT2), .B(G113), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n195), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n197), .A2(new_n190), .A3(new_n192), .A4(new_n193), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n200));
  INV_X1    g014(.A(G137), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G134), .ZN(new_n202));
  NOR2_X1   g016(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n200), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G131), .ZN(new_n205));
  INV_X1    g019(.A(G134), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G137), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n201), .A2(KEYINPUT64), .A3(KEYINPUT11), .A4(G134), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n204), .A2(new_n205), .A3(new_n207), .A4(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n205), .B1(new_n202), .B2(new_n207), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(KEYINPUT66), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n212));
  AOI211_X1 g026(.A(new_n212), .B(new_n205), .C1(new_n202), .C2(new_n207), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n209), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G128), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n216));
  INV_X1    g030(.A(G143), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G146), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G143), .ZN(new_n220));
  OAI22_X1  g034(.A1(new_n216), .A2(new_n218), .B1(new_n220), .B2(G128), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n216), .A2(new_n220), .A3(new_n218), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(G143), .B(G146), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(KEYINPUT67), .A3(new_n216), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n221), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n214), .A2(new_n227), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n220), .A2(new_n218), .A3(KEYINPUT0), .A4(G128), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT0), .B(G128), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n229), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(KEYINPUT65), .A2(G131), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n200), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n206), .A2(G137), .ZN(new_n235));
  OR2_X1    g049(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n208), .A2(new_n207), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n233), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n201), .A2(G134), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n240), .B1(new_n234), .B2(new_n235), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(new_n232), .A3(new_n204), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n231), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  NOR3_X1   g057(.A1(new_n228), .A2(KEYINPUT30), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT30), .ZN(new_n245));
  INV_X1    g059(.A(new_n221), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT67), .B1(new_n225), .B2(new_n216), .ZN(new_n247));
  AND4_X1   g061(.A1(KEYINPUT67), .A2(new_n216), .A3(new_n220), .A4(new_n218), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n210), .A2(KEYINPUT66), .ZN(new_n250));
  XNOR2_X1  g064(.A(G134), .B(G137), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n212), .B1(new_n251), .B2(new_n205), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n249), .A2(new_n209), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n231), .ZN(new_n255));
  NOR3_X1   g069(.A1(new_n237), .A2(new_n238), .A3(new_n233), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n232), .B1(new_n241), .B2(new_n204), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n245), .B1(new_n254), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n199), .B1(new_n244), .B2(new_n259), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n196), .A2(new_n198), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n254), .A2(new_n261), .A3(new_n258), .ZN(new_n262));
  NOR2_X1   g076(.A1(G237), .A2(G953), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G210), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(KEYINPUT27), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT26), .B(G101), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n265), .B(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT70), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n262), .A2(new_n270), .A3(new_n267), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n260), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(KEYINPUT71), .A3(KEYINPUT31), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT31), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n260), .A2(new_n269), .A3(new_n274), .A4(new_n271), .ZN(new_n275));
  INV_X1    g089(.A(new_n267), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT28), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n199), .B1(new_n228), .B2(new_n243), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n277), .B1(new_n278), .B2(new_n262), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n262), .A2(new_n277), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n276), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n273), .A2(new_n275), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT71), .B1(new_n272), .B2(KEYINPUT31), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n187), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT32), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT72), .ZN(new_n288));
  OAI211_X1 g102(.A(KEYINPUT32), .B(new_n187), .C1(new_n283), .C2(new_n284), .ZN(new_n289));
  INV_X1    g103(.A(new_n259), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n254), .A2(new_n245), .A3(new_n258), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n261), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n262), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n276), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n279), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(new_n267), .A3(new_n280), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT29), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n294), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G902), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n299), .B1(new_n296), .B2(new_n297), .ZN(new_n300));
  OAI21_X1  g114(.A(G472), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  AND2_X1   g115(.A1(new_n289), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n285), .A2(new_n303), .A3(new_n286), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n288), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G221), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT9), .B(G234), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n306), .B1(new_n308), .B2(new_n299), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n256), .A2(new_n257), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G101), .ZN(new_n313));
  INV_X1    g127(.A(G107), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G104), .ZN(new_n315));
  INV_X1    g129(.A(G104), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G107), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n313), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT79), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(new_n314), .A3(G104), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT3), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n319), .A2(new_n314), .A3(KEYINPUT3), .A4(G104), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT80), .B1(new_n314), .B2(G104), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT80), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(new_n316), .A3(G107), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n325), .A2(new_n327), .A3(new_n313), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n318), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n249), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT10), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n249), .A2(new_n329), .A3(KEYINPUT10), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n324), .A2(new_n328), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT4), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n325), .A2(new_n327), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n324), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G101), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n313), .B1(new_n324), .B2(new_n337), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT4), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n231), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n312), .B1(new_n334), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n341), .B1(KEYINPUT4), .B2(new_n335), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n341), .A2(KEYINPUT4), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n255), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n347), .A2(new_n311), .A3(new_n332), .A4(new_n333), .ZN(new_n348));
  XNOR2_X1  g162(.A(G110), .B(G140), .ZN(new_n349));
  INV_X1    g163(.A(G953), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n350), .A2(G227), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n349), .B(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n344), .A2(new_n348), .A3(new_n353), .ZN(new_n354));
  NOR3_X1   g168(.A1(new_n334), .A2(new_n343), .A3(new_n312), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT81), .B1(new_n249), .B2(new_n329), .ZN(new_n356));
  INV_X1    g170(.A(new_n318), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n335), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n359), .A3(new_n227), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n356), .A2(new_n360), .A3(new_n330), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n312), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT12), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n363), .B1(new_n311), .B2(KEYINPUT82), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n361), .A2(new_n312), .A3(new_n364), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n355), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI211_X1 g182(.A(G469), .B(new_n354), .C1(new_n368), .C2(new_n353), .ZN(new_n369));
  INV_X1    g183(.A(G469), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n370), .A2(new_n299), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n344), .A2(new_n348), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n352), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n361), .A2(new_n312), .A3(new_n364), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n364), .B1(new_n361), .B2(new_n312), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n353), .B(new_n348), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  AOI211_X1 g192(.A(G469), .B(G902), .C1(new_n375), .C2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n310), .B1(new_n373), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT83), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT83), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n382), .B(new_n310), .C1(new_n373), .C2(new_n379), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G217), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n385), .B1(G234), .B2(new_n299), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(G902), .ZN(new_n387));
  INV_X1    g201(.A(G119), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT74), .B1(new_n388), .B2(G128), .ZN(new_n389));
  OR2_X1    g203(.A1(new_n389), .A2(KEYINPUT23), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(G128), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(KEYINPUT23), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  OR2_X1    g207(.A1(new_n393), .A2(G110), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT73), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n395), .B1(new_n388), .B2(G128), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n215), .A2(KEYINPUT73), .A3(G119), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n391), .A3(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(KEYINPUT24), .B(G110), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT75), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT76), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n398), .A2(KEYINPUT75), .A3(new_n399), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n394), .A2(new_n402), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G125), .ZN(new_n406));
  NOR3_X1   g220(.A1(new_n406), .A2(KEYINPUT16), .A3(G140), .ZN(new_n407));
  XNOR2_X1  g221(.A(G125), .B(G140), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n407), .B1(new_n408), .B2(KEYINPUT16), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G146), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n402), .B(new_n404), .C1(new_n393), .C2(G110), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT76), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n408), .A2(new_n219), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n405), .A2(new_n410), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n393), .A2(G110), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n409), .A2(G146), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n409), .A2(G146), .ZN(new_n417));
  OAI221_X1 g231(.A(new_n415), .B1(new_n399), .B2(new_n398), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT22), .B(G137), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n350), .A2(G221), .A3(G234), .ZN(new_n421));
  XOR2_X1   g235(.A(new_n420), .B(new_n421), .Z(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n414), .A2(new_n418), .A3(new_n422), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT78), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n424), .A2(KEYINPUT78), .A3(new_n425), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n386), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT77), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT25), .ZN(new_n433));
  AOI21_X1  g247(.A(G902), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n424), .A2(new_n425), .A3(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n432), .A2(new_n433), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n431), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n436), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n424), .A2(new_n425), .A3(new_n438), .A4(new_n434), .ZN(new_n439));
  AOI22_X1  g253(.A1(new_n387), .A2(new_n430), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT93), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n441), .B1(new_n417), .B2(new_n416), .ZN(new_n442));
  OR2_X1    g256(.A1(new_n409), .A2(G146), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(KEYINPUT93), .A3(new_n410), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n263), .A2(G143), .A3(G214), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(G143), .B1(new_n263), .B2(G214), .ZN(new_n447));
  OAI21_X1  g261(.A(G131), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n263), .A2(G214), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n217), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(new_n205), .A3(new_n445), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT17), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n448), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  OR2_X1    g267(.A1(new_n448), .A2(new_n452), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n442), .A2(new_n444), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n450), .A2(KEYINPUT89), .A3(new_n445), .ZN(new_n456));
  NAND2_X1  g270(.A1(KEYINPUT18), .A2(G131), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n406), .A2(G140), .ZN(new_n459));
  INV_X1    g273(.A(G140), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(G125), .ZN(new_n461));
  OAI21_X1  g275(.A(G146), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n456), .A2(new_n458), .B1(new_n462), .B2(new_n413), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n450), .A2(KEYINPUT89), .A3(new_n457), .A4(new_n445), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  XOR2_X1   g279(.A(G113), .B(G122), .Z(new_n466));
  XOR2_X1   g280(.A(KEYINPUT92), .B(G104), .Z(new_n467));
  XOR2_X1   g281(.A(new_n466), .B(new_n467), .Z(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n455), .A2(new_n465), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n469), .B1(new_n455), .B2(new_n465), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n299), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G475), .ZN(new_n474));
  NOR2_X1   g288(.A1(G475), .A2(G902), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n448), .A2(new_n451), .B1(new_n409), .B2(G146), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n408), .A2(KEYINPUT90), .A3(KEYINPUT19), .ZN(new_n478));
  AOI21_X1  g292(.A(KEYINPUT19), .B1(new_n408), .B2(KEYINPUT90), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n219), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n465), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT91), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n477), .A2(new_n480), .B1(new_n463), .B2(new_n464), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT91), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n486), .A3(new_n468), .ZN(new_n487));
  AOI211_X1 g301(.A(KEYINPUT20), .B(new_n476), .C1(new_n487), .C2(new_n470), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT20), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n468), .B1(new_n485), .B2(KEYINPUT91), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n482), .A2(new_n483), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n470), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n489), .B1(new_n492), .B2(new_n475), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n474), .B1(new_n488), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(G128), .B(G143), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT13), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n215), .A2(KEYINPUT13), .A3(G143), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n497), .A2(new_n206), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n206), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n496), .A2(new_n498), .B1(new_n499), .B2(KEYINPUT94), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n499), .A2(KEYINPUT94), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n188), .A2(G122), .A3(new_n189), .ZN(new_n502));
  OR2_X1    g316(.A1(new_n191), .A2(G122), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n314), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n314), .B1(new_n502), .B2(new_n503), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n500), .B(new_n501), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n495), .B(new_n206), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n502), .A2(new_n503), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(KEYINPUT14), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT14), .ZN(new_n511));
  OAI21_X1  g325(.A(G107), .B1(new_n502), .B2(new_n511), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n508), .B(new_n504), .C1(new_n510), .C2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n507), .A2(new_n513), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n307), .A2(new_n385), .A3(G953), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT95), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n507), .A2(new_n513), .A3(new_n515), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n514), .A2(KEYINPUT95), .A3(new_n516), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n520), .A2(new_n299), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(G478), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n523), .A2(KEYINPUT15), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n524), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n520), .A2(new_n299), .A3(new_n521), .A4(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n350), .A2(G952), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n529), .B1(G234), .B2(G237), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT21), .B(G898), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(KEYINPUT96), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  AOI211_X1 g347(.A(new_n299), .B(new_n350), .C1(G234), .C2(G237), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n530), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OR3_X1    g349(.A1(new_n494), .A2(new_n528), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(G210), .B1(G237), .B2(G902), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(G110), .B(G122), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n261), .B1(new_n340), .B2(new_n342), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n190), .A2(new_n193), .A3(KEYINPUT5), .A4(new_n192), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n191), .A2(KEYINPUT5), .A3(G119), .ZN(new_n543));
  INV_X1    g357(.A(G113), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n198), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n547), .A2(new_n358), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n540), .B1(new_n541), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n199), .B1(new_n345), .B2(new_n346), .ZN(new_n550));
  INV_X1    g364(.A(new_n548), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n550), .A2(new_n551), .A3(new_n539), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n549), .A2(new_n552), .A3(KEYINPUT6), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n227), .A2(new_n406), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n231), .A2(G125), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n350), .A2(G224), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT6), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n559), .B(new_n540), .C1(new_n541), .C2(new_n548), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n553), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n556), .A2(KEYINPUT88), .A3(KEYINPUT7), .A4(new_n557), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n554), .A2(KEYINPUT87), .A3(new_n555), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n557), .A2(KEYINPUT7), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n563), .B(new_n564), .C1(KEYINPUT87), .C2(new_n554), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT86), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n198), .B(new_n546), .C1(new_n358), .C2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n547), .A2(KEYINPUT86), .A3(new_n329), .ZN(new_n568));
  XOR2_X1   g382(.A(KEYINPUT85), .B(KEYINPUT8), .Z(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(new_n539), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT88), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n554), .A2(new_n555), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n572), .B1(new_n573), .B2(new_n564), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n562), .A2(new_n565), .A3(new_n571), .A4(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n552), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n299), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n538), .B1(new_n561), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n577), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n553), .A2(new_n558), .A3(new_n560), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n537), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(G214), .B1(G237), .B2(G902), .ZN(new_n583));
  XOR2_X1   g397(.A(new_n583), .B(KEYINPUT84), .Z(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n536), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n305), .A2(new_n384), .A3(new_n440), .A4(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(G101), .ZN(G3));
  NAND2_X1  g403(.A1(new_n272), .A2(KEYINPUT31), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT71), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n275), .A2(new_n282), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n273), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n299), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(G472), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n596), .A2(new_n285), .A3(new_n440), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n522), .A2(new_n523), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT33), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n520), .A2(new_n599), .A3(new_n521), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n517), .A2(KEYINPUT33), .A3(new_n519), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n299), .A2(G478), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n598), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n494), .A2(new_n604), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n586), .A2(new_n535), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n597), .A2(new_n384), .A3(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(KEYINPUT97), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT34), .B(G104), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G6));
  AND2_X1   g424(.A1(new_n455), .A2(new_n465), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n469), .B1(new_n482), .B2(new_n483), .ZN(new_n612));
  AOI22_X1  g426(.A1(new_n611), .A2(new_n469), .B1(new_n612), .B2(new_n486), .ZN(new_n613));
  OAI21_X1  g427(.A(KEYINPUT20), .B1(new_n613), .B2(new_n476), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT98), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n492), .A2(new_n489), .A3(new_n475), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n493), .A2(KEYINPUT98), .B1(new_n473), .B2(G475), .ZN(new_n618));
  XOR2_X1   g432(.A(new_n535), .B(KEYINPUT99), .Z(new_n619));
  NAND4_X1  g433(.A1(new_n617), .A2(new_n618), .A3(new_n528), .A4(new_n619), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n620), .A2(KEYINPUT100), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n620), .A2(KEYINPUT100), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n621), .A2(new_n622), .A3(new_n586), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(new_n384), .A3(new_n597), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT35), .B(G107), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G9));
  NAND2_X1  g440(.A1(new_n596), .A2(new_n285), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n437), .A2(new_n439), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n423), .A2(KEYINPUT36), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n419), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n387), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n634), .A2(new_n384), .A3(new_n587), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT37), .B(G110), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G12));
  AOI21_X1  g451(.A(new_n584), .B1(new_n578), .B2(new_n581), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(G900), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n530), .B1(new_n534), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n617), .A2(new_n618), .A3(new_n528), .A4(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n305), .A2(new_n644), .A3(new_n384), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT101), .B(G128), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G30));
  INV_X1    g461(.A(new_n272), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n278), .A2(new_n262), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n648), .B1(new_n276), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(G472), .B1(new_n650), .B2(G902), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n289), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n288), .A2(new_n652), .A3(new_n304), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n632), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT38), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n582), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n578), .A2(new_n581), .A3(KEYINPUT38), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n494), .A2(new_n528), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n659), .A2(new_n584), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n655), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(KEYINPUT102), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n641), .B(KEYINPUT39), .Z(new_n665));
  NAND2_X1  g479(.A1(new_n384), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n666), .B(KEYINPUT40), .Z(new_n667));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n655), .A2(new_n668), .A3(new_n662), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n664), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G143), .ZN(G45));
  NAND3_X1  g485(.A1(new_n494), .A2(new_n604), .A3(new_n642), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n494), .A2(new_n604), .A3(KEYINPUT103), .A4(new_n642), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n639), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n677), .A2(new_n305), .A3(new_n384), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G146), .ZN(G48));
  NAND2_X1  g493(.A1(new_n375), .A2(new_n378), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n370), .B1(new_n680), .B2(new_n299), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n680), .A2(new_n370), .A3(new_n299), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n682), .A2(new_n310), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT104), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n685), .A2(new_n305), .A3(new_n440), .A4(new_n606), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT41), .B(G113), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G15));
  NAND4_X1  g502(.A1(new_n685), .A2(new_n623), .A3(new_n305), .A4(new_n440), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT105), .B(G116), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G18));
  NOR2_X1   g505(.A1(new_n681), .A2(new_n379), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n638), .A2(new_n692), .A3(new_n310), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n693), .A2(new_n536), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n305), .A2(new_n694), .A3(new_n632), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G119), .ZN(G21));
  NOR2_X1   g510(.A1(new_n661), .A2(new_n586), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n697), .A2(new_n619), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n700), .B1(new_n590), .B2(new_n282), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n590), .A2(new_n700), .A3(new_n282), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n702), .A2(new_n275), .A3(new_n703), .ZN(new_n704));
  AOI22_X1  g518(.A1(new_n704), .A2(new_n187), .B1(new_n595), .B2(G472), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n699), .B1(new_n705), .B2(new_n440), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n703), .A2(new_n275), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n187), .B1(new_n707), .B2(new_n701), .ZN(new_n708));
  AND4_X1   g522(.A1(new_n699), .A2(new_n596), .A3(new_n440), .A4(new_n708), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n698), .B(new_n685), .C1(new_n706), .C2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  NAND3_X1  g525(.A1(new_n596), .A2(new_n708), .A3(new_n632), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n712), .A2(new_n676), .A3(new_n693), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT108), .B(G125), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G27));
  NAND2_X1  g529(.A1(new_n302), .A2(new_n287), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n674), .A2(new_n675), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n717), .A3(new_n440), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT109), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n719), .B1(new_n373), .B2(new_n379), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n683), .A2(KEYINPUT109), .A3(new_n372), .A4(new_n369), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n720), .A2(new_n310), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n578), .A2(new_n581), .A3(new_n585), .ZN(new_n723));
  OR2_X1    g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g538(.A(KEYINPUT42), .B1(new_n718), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n676), .A2(KEYINPUT42), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n722), .A2(new_n723), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n726), .A2(new_n727), .A3(new_n305), .A4(new_n440), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(new_n205), .ZN(G33));
  INV_X1    g544(.A(new_n643), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n727), .A2(new_n305), .A3(new_n440), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G134), .ZN(G36));
  INV_X1    g547(.A(new_n494), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n604), .ZN(new_n735));
  XOR2_X1   g549(.A(new_n735), .B(KEYINPUT43), .Z(new_n736));
  AND3_X1   g550(.A1(new_n736), .A2(new_n627), .A3(new_n632), .ZN(new_n737));
  OR2_X1    g551(.A1(new_n737), .A2(KEYINPUT44), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n723), .B1(new_n737), .B2(KEYINPUT44), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n348), .B1(new_n376), .B2(new_n377), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n355), .A2(new_n352), .ZN(new_n741));
  AOI22_X1  g555(.A1(new_n352), .A2(new_n740), .B1(new_n741), .B2(new_n344), .ZN(new_n742));
  OAI21_X1  g556(.A(G469), .B1(new_n742), .B2(KEYINPUT45), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n743), .B1(KEYINPUT45), .B2(new_n742), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n371), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(KEYINPUT46), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n379), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(KEYINPUT46), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n309), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n738), .A2(new_n739), .A3(new_n665), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G137), .ZN(G39));
  NAND2_X1  g565(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  NOR4_X1   g567(.A1(new_n305), .A2(new_n440), .A3(new_n676), .A4(new_n723), .ZN(new_n754));
  XOR2_X1   g568(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n755));
  OAI211_X1 g569(.A(new_n753), .B(new_n754), .C1(new_n749), .C2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G140), .ZN(G42));
  NAND2_X1  g571(.A1(new_n734), .A2(new_n528), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n605), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n638), .A2(new_n619), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n597), .A2(new_n384), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n588), .A2(new_n635), .A3(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT112), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n588), .A2(new_n635), .A3(new_n761), .A4(KEYINPUT112), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n710), .A2(new_n686), .A3(new_n689), .A4(new_n695), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n725), .A2(new_n728), .A3(new_n732), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n724), .A2(new_n676), .A3(new_n712), .ZN(new_n770));
  INV_X1    g584(.A(new_n723), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n525), .A2(new_n527), .A3(new_n642), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n617), .A2(new_n772), .A3(new_n618), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n771), .A2(KEYINPUT113), .A3(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n617), .A2(new_n772), .A3(new_n618), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n775), .B1(new_n723), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n778), .A2(new_n305), .A3(new_n384), .A4(new_n632), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI22_X1  g595(.A1(new_n774), .A2(new_n777), .B1(new_n381), .B2(new_n383), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n782), .A2(KEYINPUT114), .A3(new_n305), .A4(new_n632), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n770), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n766), .A2(new_n768), .A3(new_n769), .A4(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n638), .A2(new_n660), .A3(new_n642), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n722), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n653), .A3(new_n633), .ZN(new_n792));
  INV_X1    g606(.A(new_n693), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n717), .A2(new_n793), .A3(new_n705), .A4(new_n632), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n678), .A2(new_n792), .A3(new_n645), .A4(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n795), .A2(KEYINPUT115), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(KEYINPUT115), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n789), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n795), .A2(KEYINPUT52), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n788), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI211_X1 g614(.A(KEYINPUT72), .B(KEYINPUT32), .C1(new_n594), .C2(new_n187), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n303), .B1(new_n285), .B2(new_n286), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI22_X1  g617(.A1(new_n803), .A2(new_n302), .B1(new_n383), .B2(new_n381), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n713), .B1(new_n804), .B2(new_n644), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n805), .A2(new_n806), .A3(new_n678), .A4(new_n792), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n795), .A2(KEYINPUT115), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT52), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n799), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n809), .A2(KEYINPUT116), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n787), .B1(new_n800), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n769), .A2(new_n784), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n767), .B1(new_n764), .B2(new_n765), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n807), .A2(new_n808), .A3(KEYINPUT52), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n798), .A2(new_n814), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n786), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n812), .A2(new_n813), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n798), .A2(new_n788), .A3(new_n799), .ZN(new_n820));
  OAI21_X1  g634(.A(KEYINPUT116), .B1(new_n809), .B2(new_n810), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n785), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  MUX2_X1   g636(.A(new_n817), .B(new_n822), .S(new_n786), .Z(new_n823));
  OAI21_X1  g637(.A(new_n819), .B1(new_n823), .B2(new_n813), .ZN(new_n824));
  INV_X1    g638(.A(new_n684), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(KEYINPUT118), .A3(new_n771), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n827), .B1(new_n684), .B2(new_n723), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n826), .A2(new_n530), .A3(new_n828), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n829), .A2(new_n440), .A3(new_n654), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n494), .A2(new_n604), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n829), .A2(new_n736), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n832), .B1(new_n712), .B2(new_n833), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n706), .A2(new_n709), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n835), .A2(new_n530), .A3(new_n736), .ZN(new_n836));
  INV_X1    g650(.A(new_n659), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(new_n585), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n836), .A2(new_n825), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT50), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n836), .A2(KEYINPUT50), .A3(new_n825), .A4(new_n838), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n834), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n692), .A2(new_n309), .ZN(new_n844));
  INV_X1    g658(.A(new_n753), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n749), .A2(new_n755), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n836), .A2(new_n771), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n843), .A2(new_n849), .A3(KEYINPUT51), .ZN(new_n850));
  AND4_X1   g664(.A1(new_n440), .A2(new_n829), .A3(new_n716), .A4(new_n736), .ZN(new_n851));
  XOR2_X1   g665(.A(new_n851), .B(KEYINPUT48), .Z(new_n852));
  NAND3_X1  g666(.A1(new_n836), .A2(new_n638), .A3(new_n825), .ZN(new_n853));
  INV_X1    g667(.A(new_n605), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n529), .B1(new_n830), .B2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n850), .A2(new_n852), .A3(new_n853), .A4(new_n855), .ZN(new_n856));
  XOR2_X1   g670(.A(new_n844), .B(KEYINPUT117), .Z(new_n857));
  OAI21_X1  g671(.A(new_n857), .B1(new_n845), .B2(new_n846), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n848), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT51), .B1(new_n843), .B2(new_n859), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  OAI22_X1  g675(.A1(new_n824), .A2(new_n861), .B1(G952), .B2(G953), .ZN(new_n862));
  INV_X1    g676(.A(new_n735), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n863), .A2(new_n440), .A3(new_n310), .A4(new_n585), .ZN(new_n864));
  INV_X1    g678(.A(new_n692), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n864), .B1(KEYINPUT49), .B2(new_n865), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n866), .B(KEYINPUT111), .Z(new_n867));
  OAI21_X1  g681(.A(new_n659), .B1(KEYINPUT49), .B2(new_n865), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n868), .A2(new_n653), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n862), .B1(new_n867), .B2(new_n869), .ZN(G75));
  AOI21_X1  g684(.A(new_n299), .B1(new_n812), .B2(new_n818), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(G210), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT56), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n558), .B(KEYINPUT120), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT55), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n553), .A2(new_n560), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n877), .B(KEYINPUT119), .Z(new_n878));
  XNOR2_X1  g692(.A(new_n876), .B(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n874), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n350), .A2(G952), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n879), .B1(new_n872), .B2(new_n873), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(G51));
  NAND2_X1  g698(.A1(new_n812), .A2(new_n818), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(new_n813), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n371), .B(KEYINPUT57), .Z(new_n887));
  OAI21_X1  g701(.A(new_n680), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n871), .A2(new_n744), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n882), .B1(new_n888), .B2(new_n889), .ZN(G54));
  NAND3_X1  g704(.A1(new_n871), .A2(KEYINPUT58), .A3(G475), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n891), .A2(new_n613), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n891), .A2(new_n613), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n892), .A2(new_n893), .A3(new_n882), .ZN(G60));
  NAND2_X1  g708(.A1(G478), .A2(G902), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT59), .Z(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  AOI22_X1  g711(.A1(new_n824), .A2(new_n897), .B1(new_n600), .B2(new_n601), .ZN(new_n898));
  INV_X1    g712(.A(new_n882), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n600), .A2(new_n601), .A3(new_n897), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n899), .B1(new_n886), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n898), .A2(new_n901), .ZN(G63));
  INV_X1    g716(.A(KEYINPUT61), .ZN(new_n903));
  NAND2_X1  g717(.A1(G217), .A2(G902), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT60), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(new_n812), .B2(new_n818), .ZN(new_n906));
  OAI211_X1 g720(.A(KEYINPUT121), .B(new_n899), .C1(new_n906), .C2(new_n430), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n630), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n905), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n785), .A2(new_n809), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT53), .B1(new_n911), .B2(new_n816), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n814), .A2(new_n815), .A3(KEYINPUT53), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n913), .B1(new_n820), .B2(new_n821), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n910), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n430), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT121), .B1(new_n917), .B2(new_n899), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n903), .B1(new_n909), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n430), .B1(new_n885), .B2(new_n910), .ZN(new_n920));
  OR2_X1    g734(.A1(new_n920), .A2(KEYINPUT122), .ZN(new_n921));
  AOI211_X1 g735(.A(new_n903), .B(new_n882), .C1(new_n906), .C2(new_n630), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n920), .A2(KEYINPUT122), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n919), .A2(new_n924), .ZN(G66));
  AOI21_X1  g739(.A(new_n350), .B1(new_n532), .B2(G224), .ZN(new_n926));
  INV_X1    g740(.A(new_n815), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n926), .B1(new_n927), .B2(new_n350), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n878), .B1(G898), .B2(new_n350), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT123), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n928), .B(new_n930), .ZN(G69));
  NAND2_X1  g745(.A1(new_n756), .A2(new_n750), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n805), .A2(new_n678), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n933), .B1(new_n670), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n305), .A2(new_n440), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n759), .A2(new_n771), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n936), .A2(new_n666), .A3(new_n937), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n932), .A2(new_n935), .A3(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n670), .A2(new_n933), .A3(new_n934), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT124), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n939), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n290), .A2(new_n291), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n478), .A2(new_n479), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n944), .A2(new_n350), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n769), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n749), .A2(new_n665), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n716), .A2(new_n440), .A3(new_n697), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n934), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OR3_X1    g766(.A1(new_n932), .A2(new_n949), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n350), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n947), .B1(new_n640), .B2(G953), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n350), .B1(G227), .B2(G900), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT125), .ZN(new_n958));
  AOI22_X1  g772(.A1(new_n948), .A2(new_n956), .B1(KEYINPUT126), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n958), .A2(KEYINPUT126), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(G72));
  NAND2_X1  g775(.A1(G472), .A2(G902), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT63), .Z(new_n963));
  OAI21_X1  g777(.A(new_n963), .B1(new_n944), .B2(new_n927), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT127), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n292), .A2(new_n293), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  OAI211_X1 g782(.A(KEYINPUT127), .B(new_n963), .C1(new_n944), .C2(new_n927), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n966), .A2(new_n267), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n963), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n294), .A2(new_n272), .ZN(new_n972));
  OR3_X1    g786(.A1(new_n823), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n963), .B1(new_n953), .B2(new_n927), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n968), .A2(new_n267), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n882), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n970), .A2(new_n973), .A3(new_n976), .ZN(G57));
endmodule


