//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 0 0 1 1 0 1 1 1 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n553, new_n554, new_n555, new_n556, new_n559, new_n560, new_n561,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n571,
    new_n572, new_n573, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n590, new_n591, new_n592, new_n593, new_n594, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170, new_n1171, new_n1172;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  AND2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n461), .A2(G137), .B1(G101), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n458), .B2(new_n459), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(KEYINPUT67), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n470));
  AOI211_X1 g045(.A(new_n470), .B(new_n465), .C1(new_n466), .C2(new_n467), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n464), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  OAI21_X1  g048(.A(G2104), .B1(new_n465), .B2(G112), .ZN(new_n474));
  OR3_X1    g049(.A1(KEYINPUT68), .A2(G100), .A3(G2105), .ZN(new_n475));
  OAI21_X1  g050(.A(KEYINPUT68), .B1(G100), .B2(G2105), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n460), .A2(new_n465), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  AOI211_X1 g055(.A(new_n477), .B(new_n480), .C1(G136), .C2(new_n461), .ZN(G162));
  OR2_X1    g056(.A1(G102), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G114), .C2(new_n465), .ZN(new_n483));
  OAI211_X1 g058(.A(G126), .B(G2105), .C1(new_n458), .C2(new_n459), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT69), .ZN(new_n487));
  OAI211_X1 g062(.A(G138), .B(new_n465), .C1(new_n458), .C2(new_n459), .ZN(new_n488));
  OR2_X1    g063(.A1(new_n488), .A2(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n485), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n487), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G164));
  INV_X1    g070(.A(KEYINPUT5), .ZN(new_n496));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(KEYINPUT70), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(KEYINPUT5), .A3(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n501), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  OR3_X1    g078(.A1(new_n502), .A2(KEYINPUT71), .A3(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT71), .B1(new_n502), .B2(new_n503), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(new_n503), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n498), .A2(new_n500), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n497), .B1(new_n507), .B2(new_n508), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n509), .A2(G88), .B1(new_n510), .B2(G50), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n504), .A2(new_n505), .A3(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G166));
  NAND2_X1  g088(.A1(new_n509), .A2(G89), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n501), .A2(G63), .A3(G651), .ZN(new_n515));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT7), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n510), .A2(G51), .ZN(new_n518));
  AND4_X1   g093(.A1(new_n514), .A2(new_n515), .A3(new_n517), .A4(new_n518), .ZN(G168));
  AOI22_X1  g094(.A1(new_n509), .A2(G90), .B1(new_n510), .B2(G52), .ZN(new_n520));
  INV_X1    g095(.A(G64), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n521), .B1(new_n498), .B2(new_n500), .ZN(new_n522));
  AND2_X1   g097(.A1(G77), .A2(G543), .ZN(new_n523));
  OAI21_X1  g098(.A(G651), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(G171));
  AND3_X1   g101(.A1(new_n499), .A2(KEYINPUT5), .A3(G543), .ZN(new_n527));
  AOI21_X1  g102(.A(KEYINPUT5), .B1(new_n499), .B2(G543), .ZN(new_n528));
  OAI21_X1  g103(.A(G56), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(G68), .A2(G543), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n503), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT6), .B(G651), .ZN(new_n532));
  OAI211_X1 g107(.A(new_n532), .B(G81), .C1(new_n527), .C2(new_n528), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n532), .A2(G43), .A3(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G860), .ZN(G153));
  NAND4_X1  g112(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g113(.A1(G1), .A2(G3), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT8), .ZN(new_n540));
  NAND4_X1  g115(.A1(G319), .A2(G483), .A3(G661), .A4(new_n540), .ZN(G188));
  NAND2_X1  g116(.A1(new_n510), .A2(G53), .ZN(new_n542));
  AND2_X1   g117(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n510), .A2(G53), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n501), .A2(G65), .ZN(new_n548));
  AND2_X1   g123(.A1(G78), .A2(G543), .ZN(new_n549));
  OAI21_X1  g124(.A(G651), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n509), .A2(G91), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n547), .A2(new_n550), .A3(new_n551), .ZN(G299));
  NAND2_X1  g127(.A1(new_n525), .A2(KEYINPUT73), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT73), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n520), .A2(new_n554), .A3(new_n524), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(G301));
  INV_X1    g132(.A(G168), .ZN(G286));
  NAND2_X1  g133(.A1(new_n512), .A2(KEYINPUT74), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n504), .A2(new_n560), .A3(new_n505), .A4(new_n511), .ZN(new_n561));
  AND2_X1   g136(.A1(new_n559), .A2(new_n561), .ZN(G303));
  AOI22_X1  g137(.A1(new_n509), .A2(G87), .B1(new_n510), .B2(G49), .ZN(new_n563));
  OAI21_X1  g138(.A(G651), .B1(new_n501), .B2(G74), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(G288));
  AOI22_X1  g140(.A1(new_n501), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n566), .A2(new_n503), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n509), .A2(G86), .B1(new_n510), .B2(G48), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(G305));
  XOR2_X1   g145(.A(KEYINPUT75), .B(G85), .Z(new_n571));
  AOI22_X1  g146(.A1(new_n509), .A2(new_n571), .B1(new_n510), .B2(G47), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n501), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n503), .B2(new_n573), .ZN(G290));
  AOI21_X1  g149(.A(KEYINPUT10), .B1(new_n509), .B2(G92), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n509), .A2(KEYINPUT10), .A3(G92), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(G66), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(new_n498), .B2(new_n500), .ZN(new_n580));
  NAND2_X1  g155(.A1(G79), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n510), .A2(G54), .ZN(new_n584));
  AND3_X1   g159(.A1(new_n583), .A2(KEYINPUT76), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(KEYINPUT76), .B1(new_n583), .B2(new_n584), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n578), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  MUX2_X1   g162(.A(new_n587), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g163(.A(new_n587), .B(G301), .S(G868), .Z(G321));
  INV_X1    g164(.A(G868), .ZN(new_n590));
  NOR3_X1   g165(.A1(G168), .A2(KEYINPUT77), .A3(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT77), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(G286), .B2(G868), .ZN(new_n593));
  NAND2_X1  g168(.A1(G299), .A2(new_n590), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n591), .B1(new_n593), .B2(new_n594), .ZN(G297));
  AOI21_X1  g170(.A(new_n591), .B1(new_n593), .B2(new_n594), .ZN(G280));
  AND4_X1   g171(.A1(KEYINPUT10), .A2(new_n501), .A3(G92), .A4(new_n532), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(new_n575), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT76), .ZN(new_n599));
  OAI21_X1  g174(.A(G66), .B1(new_n527), .B2(new_n528), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n503), .B1(new_n600), .B2(new_n581), .ZN(new_n601));
  INV_X1    g176(.A(new_n584), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n599), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n583), .A2(KEYINPUT76), .A3(new_n584), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n598), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G860), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT78), .ZN(G148));
  NAND2_X1  g183(.A1(new_n605), .A2(new_n606), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G868), .B2(new_n536), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XOR2_X1   g187(.A(KEYINPUT79), .B(KEYINPUT12), .Z(new_n613));
  NAND3_X1  g188(.A1(new_n465), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT13), .ZN(new_n616));
  INV_X1    g191(.A(G2100), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n461), .A2(G135), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n478), .A2(G123), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n465), .A2(G111), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n620), .B(new_n621), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(G2096), .Z(new_n625));
  NAND3_X1  g200(.A1(new_n618), .A2(new_n619), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT80), .ZN(G156));
  XOR2_X1   g202(.A(KEYINPUT81), .B(KEYINPUT14), .Z(new_n628));
  XOR2_X1   g203(.A(KEYINPUT15), .B(G2435), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2438), .ZN(new_n630));
  XOR2_X1   g205(.A(G2427), .B(G2430), .Z(new_n631));
  AOI21_X1  g206(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(new_n630), .B2(new_n631), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XOR2_X1   g210(.A(G1341), .B(G1348), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n633), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G2443), .B(G2446), .Z(new_n639));
  OAI21_X1  g214(.A(G14), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n640), .B1(new_n639), .B2(new_n638), .ZN(G401));
  XOR2_X1   g216(.A(G2084), .B(G2090), .Z(new_n642));
  XNOR2_X1  g217(.A(G2067), .B(G2678), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  AOI21_X1  g220(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT82), .B(KEYINPUT17), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n645), .B(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n646), .B1(new_n648), .B2(new_n644), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT83), .Z(new_n650));
  INV_X1    g225(.A(new_n642), .ZN(new_n651));
  NOR3_X1   g226(.A1(new_n651), .A2(new_n644), .A3(new_n645), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT18), .Z(new_n653));
  NOR2_X1   g228(.A1(new_n651), .A2(new_n643), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n653), .B1(new_n648), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2096), .B(G2100), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1961), .B(G1966), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT84), .ZN(new_n660));
  XOR2_X1   g235(.A(G1956), .B(G2474), .Z(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n662), .A2(KEYINPUT85), .ZN(new_n663));
  XOR2_X1   g238(.A(G1971), .B(G1976), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(KEYINPUT85), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n663), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT20), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n660), .A2(new_n661), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n669), .B1(new_n662), .B2(new_n665), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n665), .A2(KEYINPUT86), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT87), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n673), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1991), .B(G1996), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1981), .B(G1986), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n681), .ZN(G229));
  INV_X1    g257(.A(G29), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G35), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(G162), .B2(new_n683), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT29), .Z(new_n686));
  INV_X1    g261(.A(G2090), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT102), .ZN(new_n689));
  INV_X1    g264(.A(G1348), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n605), .A2(G16), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(G4), .B2(G16), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n689), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(new_n690), .B2(new_n692), .ZN(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G20), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT23), .Z(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G299), .B2(G16), .ZN(new_n698));
  INV_X1    g273(.A(G1956), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n695), .A2(G19), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(new_n536), .B2(new_n695), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(G1341), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n683), .A2(G26), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT91), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n461), .A2(G140), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n478), .A2(G128), .ZN(new_n708));
  OR2_X1    g283(.A1(G104), .A2(G2105), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n709), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n707), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n706), .B1(new_n712), .B2(new_n683), .ZN(new_n713));
  INV_X1    g288(.A(G2067), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n703), .B(new_n715), .C1(new_n686), .C2(new_n687), .ZN(new_n716));
  NOR3_X1   g291(.A1(new_n694), .A2(new_n700), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n695), .A2(G21), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G168), .B2(new_n695), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT98), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n720), .A2(G1966), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n720), .A2(G1966), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT30), .B(G28), .ZN(new_n723));
  OR2_X1    g298(.A1(KEYINPUT31), .A2(G11), .ZN(new_n724));
  NAND2_X1  g299(.A1(KEYINPUT31), .A2(G11), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n723), .A2(new_n683), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n695), .A2(G5), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G171), .B2(new_n695), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G1961), .ZN(new_n730));
  OAI221_X1 g305(.A(new_n726), .B1(new_n683), .B2(new_n624), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  NOR3_X1   g306(.A1(new_n721), .A2(new_n722), .A3(new_n731), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT99), .Z(new_n733));
  NOR2_X1   g308(.A1(G29), .A2(G32), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n478), .A2(G129), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT95), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n461), .A2(G141), .ZN(new_n737));
  NAND3_X1  g312(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT26), .Z(new_n739));
  NAND2_X1  g314(.A1(new_n463), .A2(G105), .ZN(new_n740));
  NAND4_X1  g315(.A1(new_n736), .A2(new_n737), .A3(new_n739), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT96), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n734), .B1(new_n742), .B2(G29), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT27), .B(G1996), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n683), .A2(G27), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G164), .B2(new_n683), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT100), .B(G2078), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n730), .B2(new_n729), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT24), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n683), .B1(new_n752), .B2(G34), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(KEYINPUT93), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(KEYINPUT93), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n752), .B2(G34), .ZN(new_n756));
  AOI22_X1  g331(.A1(G160), .A2(G29), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT94), .Z(new_n758));
  INV_X1    g333(.A(G2084), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n746), .A2(new_n751), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n683), .A2(G33), .ZN(new_n762));
  NAND2_X1  g337(.A1(G115), .A2(G2104), .ZN(new_n763));
  INV_X1    g338(.A(G127), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n460), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n465), .B1(new_n765), .B2(KEYINPUT92), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(KEYINPUT92), .B2(new_n765), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT25), .ZN(new_n768));
  NAND2_X1  g343(.A1(G103), .A2(G2104), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n769), .B2(G2105), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n465), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n461), .A2(G139), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n767), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n762), .B1(new_n773), .B2(new_n683), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(G2072), .Z(new_n775));
  OAI221_X1 g350(.A(new_n775), .B1(new_n758), .B2(new_n759), .C1(new_n743), .C2(new_n745), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT97), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n761), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n733), .B(new_n778), .C1(new_n777), .C2(new_n776), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT101), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n461), .A2(G131), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n478), .A2(G119), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n465), .A2(G107), .ZN(new_n783));
  OAI21_X1  g358(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n781), .B(new_n782), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  MUX2_X1   g360(.A(G25), .B(new_n785), .S(G29), .Z(new_n786));
  XOR2_X1   g361(.A(KEYINPUT35), .B(G1991), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  MUX2_X1   g363(.A(G24), .B(G290), .S(G16), .Z(new_n789));
  XOR2_X1   g364(.A(KEYINPUT88), .B(G1986), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(G166), .A2(G16), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G16), .B2(G22), .ZN(new_n793));
  INV_X1    g368(.A(G1971), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  MUX2_X1   g370(.A(G6), .B(G305), .S(G16), .Z(new_n796));
  XOR2_X1   g371(.A(KEYINPUT32), .B(G1981), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n793), .A2(new_n794), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n695), .A2(G23), .ZN(new_n800));
  INV_X1    g375(.A(G288), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(new_n695), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT33), .B(G1976), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT89), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n802), .B(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n795), .A2(new_n798), .A3(new_n799), .A4(new_n805), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n788), .B(new_n791), .C1(new_n806), .C2(KEYINPUT34), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(KEYINPUT34), .B2(new_n806), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT90), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(KEYINPUT36), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n808), .B(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n717), .A2(new_n780), .A3(new_n811), .ZN(G150));
  INV_X1    g387(.A(G150), .ZN(G311));
  AOI22_X1  g388(.A1(new_n509), .A2(G93), .B1(new_n510), .B2(G55), .ZN(new_n814));
  INV_X1    g389(.A(G67), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n498), .B2(new_n500), .ZN(new_n816));
  NAND2_X1  g391(.A1(G80), .A2(G543), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(G651), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(KEYINPUT104), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT104), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n814), .A2(new_n822), .A3(new_n819), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(G860), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT37), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n605), .A2(G559), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT38), .Z(new_n829));
  INV_X1    g404(.A(new_n530), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(new_n501), .B2(G56), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n534), .B(new_n533), .C1(new_n831), .C2(new_n503), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n821), .A2(new_n832), .A3(new_n823), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n536), .A2(KEYINPUT103), .A3(new_n820), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT103), .ZN(new_n835));
  OAI21_X1  g410(.A(G67), .B1(new_n527), .B2(new_n528), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n503), .B1(new_n836), .B2(new_n817), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n532), .B(G93), .C1(new_n527), .C2(new_n528), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n532), .A2(G55), .A3(G543), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n835), .B1(new_n841), .B2(new_n832), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n833), .A2(new_n834), .A3(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n829), .B(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n825), .B1(new_n845), .B2(KEYINPUT39), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n827), .B1(new_n846), .B2(new_n847), .ZN(G145));
  NOR2_X1   g423(.A1(new_n741), .A2(new_n773), .ZN(new_n849));
  INV_X1    g424(.A(new_n742), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n849), .B1(new_n850), .B2(new_n773), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n485), .B1(new_n489), .B2(new_n490), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n785), .B(new_n615), .Z(new_n854));
  NAND2_X1  g429(.A1(new_n478), .A2(G130), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT105), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  INV_X1    g432(.A(G118), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n857), .B1(new_n858), .B2(G2105), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(new_n461), .B2(G142), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n854), .B(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(new_n711), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n862), .A2(new_n711), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n853), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n864), .A2(new_n853), .A3(new_n865), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n851), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  INV_X1    g445(.A(new_n851), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(new_n866), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n472), .B(new_n624), .Z(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(G162), .ZN(new_n875));
  AOI21_X1  g450(.A(G37), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n875), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n869), .A2(new_n872), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(KEYINPUT106), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n876), .A2(new_n881), .A3(new_n878), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n880), .A2(KEYINPUT40), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(KEYINPUT40), .B1(new_n880), .B2(new_n882), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(G395));
  OR2_X1    g460(.A1(new_n824), .A2(G868), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n843), .B(new_n609), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT107), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(new_n605), .B2(G299), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n605), .A2(G299), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n547), .A2(new_n550), .A3(new_n551), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n587), .A2(new_n891), .A3(KEYINPUT107), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n887), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(KEYINPUT41), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT41), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n889), .A2(new_n892), .A3(new_n896), .A4(new_n890), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n894), .B1(new_n887), .B2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(G305), .B(KEYINPUT108), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n512), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT108), .ZN(new_n902));
  XNOR2_X1  g477(.A(G305), .B(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(G166), .ZN(new_n904));
  XNOR2_X1  g479(.A(G290), .B(G288), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n901), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n905), .B1(new_n901), .B2(new_n904), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n899), .B(new_n908), .ZN(new_n909));
  XOR2_X1   g484(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n910));
  XNOR2_X1  g485(.A(new_n909), .B(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n886), .B1(new_n911), .B2(new_n590), .ZN(G295));
  OAI21_X1  g487(.A(new_n886), .B1(new_n911), .B2(new_n590), .ZN(G331));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n520), .A2(new_n554), .A3(new_n524), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n554), .B1(new_n520), .B2(new_n524), .ZN(new_n916));
  OAI21_X1  g491(.A(G168), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n515), .A2(new_n518), .A3(new_n517), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n918), .A2(new_n514), .B1(new_n524), .B2(new_n520), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  NOR3_X1   g496(.A1(new_n841), .A2(new_n832), .A3(new_n835), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT103), .B1(new_n536), .B2(new_n820), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(new_n924), .A3(new_n833), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n919), .B1(new_n556), .B2(G168), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n843), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n895), .A2(new_n928), .A3(new_n897), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n893), .A2(new_n925), .A3(new_n927), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT110), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n893), .A2(new_n925), .A3(new_n927), .A4(KEYINPUT110), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n929), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  OR2_X1    g509(.A1(new_n934), .A2(new_n908), .ZN(new_n935));
  INV_X1    g510(.A(G37), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n929), .A2(new_n930), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(new_n908), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n935), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n914), .B1(new_n939), .B2(KEYINPUT43), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n934), .A2(new_n908), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT111), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n941), .A2(new_n942), .A3(new_n936), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n935), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n942), .B1(new_n941), .B2(new_n936), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n940), .B1(new_n946), .B2(KEYINPUT43), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT43), .B1(new_n944), .B2(new_n945), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n935), .A2(new_n949), .A3(new_n936), .A4(new_n938), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT112), .B1(new_n951), .B2(new_n914), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT112), .ZN(new_n953));
  AOI211_X1 g528(.A(new_n953), .B(KEYINPUT44), .C1(new_n948), .C2(new_n950), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n947), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT113), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI211_X1 g532(.A(KEYINPUT113), .B(new_n947), .C1(new_n952), .C2(new_n954), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(G397));
  XNOR2_X1  g534(.A(new_n711), .B(G2067), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n960), .B1(G1996), .B2(new_n741), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(new_n850), .B2(G1996), .ZN(new_n962));
  INV_X1    g537(.A(new_n787), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n785), .B(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT114), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G1384), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n853), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT45), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI211_X1 g545(.A(G40), .B(new_n464), .C1(new_n469), .C2(new_n471), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n966), .A2(new_n973), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n973), .A2(G1986), .A3(G290), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n975), .B(KEYINPUT48), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n972), .B1(new_n960), .B2(new_n741), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n973), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT46), .ZN(new_n980));
  INV_X1    g555(.A(G1996), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n980), .B1(new_n972), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n978), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  XOR2_X1   g558(.A(new_n983), .B(KEYINPUT47), .Z(new_n984));
  OR2_X1    g559(.A1(new_n785), .A2(new_n963), .ZN(new_n985));
  OAI22_X1  g560(.A1(new_n962), .A2(new_n985), .B1(G2067), .B2(new_n711), .ZN(new_n986));
  AOI211_X1 g561(.A(new_n977), .B(new_n984), .C1(new_n972), .C2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT127), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT63), .ZN(new_n989));
  INV_X1    g564(.A(G1976), .ZN(new_n990));
  OAI221_X1 g565(.A(G8), .B1(new_n990), .B2(G288), .C1(new_n968), .C2(new_n971), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT52), .ZN(new_n992));
  INV_X1    g567(.A(new_n971), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n852), .A2(G1384), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G1981), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n568), .A2(new_n996), .A3(new_n569), .ZN(new_n997));
  INV_X1    g572(.A(new_n569), .ZN(new_n998));
  OAI21_X1  g573(.A(G1981), .B1(new_n998), .B2(new_n567), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT116), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT49), .ZN(new_n1001));
  OAI211_X1 g576(.A(G8), .B(new_n995), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n992), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT52), .B1(G288), .B2(new_n990), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT115), .B1(new_n991), .B2(new_n1006), .ZN(new_n1007));
  OR3_X1    g582(.A1(new_n991), .A2(KEYINPUT115), .A3(new_n1006), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1004), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G8), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n971), .B1(new_n968), .B2(KEYINPUT50), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n494), .A2(new_n1012), .A3(new_n967), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1011), .A2(new_n687), .A3(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n969), .A2(G1384), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n853), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n993), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT45), .B1(new_n494), .B2(new_n967), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n794), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1010), .B1(new_n1014), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n559), .A2(G8), .A3(new_n561), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n559), .A2(KEYINPUT55), .A3(G8), .A4(new_n561), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1021), .A2(new_n1027), .A3(KEYINPUT117), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1029), .B1(new_n1020), .B2(new_n1026), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1012), .B1(new_n494), .B2(new_n967), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n852), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n1031), .A2(new_n1032), .A3(new_n971), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n687), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1010), .B1(new_n1034), .B2(new_n1019), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n1026), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1009), .A2(new_n1028), .A3(new_n1030), .A4(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n971), .B1(new_n968), .B2(new_n969), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n494), .A2(new_n1015), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT118), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n494), .A2(new_n1041), .A3(new_n1015), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1038), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1966), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1033), .A2(new_n759), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1010), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(G168), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n989), .B1(new_n1037), .B2(new_n1048), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1009), .A2(new_n1036), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1035), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n989), .B1(new_n1051), .B2(new_n1027), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1050), .A2(G168), .A3(new_n1047), .A4(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n968), .A2(new_n971), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n990), .B(new_n801), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1056));
  AOI211_X1 g631(.A(new_n1010), .B(new_n1055), .C1(new_n1056), .C2(new_n997), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1036), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1057), .B1(new_n1058), .B2(new_n1009), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1054), .A2(new_n1059), .ZN(new_n1060));
  AND3_X1   g635(.A1(G299), .A2(KEYINPUT119), .A3(KEYINPUT57), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT57), .B1(G299), .B2(KEYINPUT119), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1018), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n971), .B1(new_n853), .B2(new_n1015), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT56), .B(G2072), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(G1956), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1064), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1033), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1071), .A2(new_n690), .B1(new_n714), .B2(new_n1055), .ZN(new_n1072));
  OR2_X1    g647(.A1(new_n1072), .A2(new_n587), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n993), .B1(new_n1012), .B2(new_n994), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1013), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n699), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1076), .A2(new_n1063), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1070), .B1(new_n1073), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1070), .A2(KEYINPUT61), .A3(new_n1078), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1072), .A2(KEYINPUT60), .ZN(new_n1082));
  OAI221_X1 g657(.A(KEYINPUT60), .B1(G2067), .B2(new_n995), .C1(new_n1033), .C2(G1348), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n605), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1081), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  NOR3_X1   g660(.A1(new_n1017), .A2(new_n1018), .A3(G1996), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT58), .B(G1341), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1055), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n536), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OAI211_X1 g666(.A(KEYINPUT59), .B(new_n536), .C1(new_n1086), .C2(new_n1088), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1091), .B(new_n1092), .C1(new_n605), .C2(new_n1083), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1085), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1095), .B1(new_n1096), .B2(new_n1064), .ZN(new_n1097));
  AOI211_X1 g672(.A(KEYINPUT120), .B(new_n1063), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1078), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT61), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1080), .B1(new_n1094), .B2(new_n1101), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1103));
  INV_X1    g678(.A(G2078), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1065), .A2(new_n1104), .A3(new_n1066), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1106), .A2(G2078), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1038), .A2(new_n1040), .A3(new_n1042), .A4(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n993), .B1(new_n968), .B2(KEYINPUT50), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n730), .B1(new_n1110), .B2(new_n1031), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1107), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT126), .B1(new_n1112), .B2(new_n556), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n1071), .A2(new_n730), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT126), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1114), .A2(new_n1115), .A3(G301), .A4(new_n1109), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n464), .A2(G40), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1118), .A2(new_n468), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n970), .A2(KEYINPUT125), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT125), .B1(new_n970), .B2(new_n1119), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1016), .B(new_n1108), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n1114), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(G171), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT54), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1050), .B(new_n1103), .C1(new_n1117), .C2(new_n1126), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1112), .A2(KEYINPUT124), .A3(new_n556), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT124), .B1(new_n1112), .B2(new_n556), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1123), .A2(new_n1114), .A3(G301), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT54), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1102), .A2(new_n1127), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n1134));
  NAND2_X1  g709(.A1(G286), .A2(G8), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1135), .B(KEYINPUT121), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT122), .B1(new_n1047), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1043), .A2(new_n1044), .B1(new_n1033), .B2(new_n759), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1139), .B(new_n1136), .C1(new_n1140), .C2(new_n1010), .ZN(new_n1141));
  AND3_X1   g716(.A1(new_n1138), .A2(KEYINPUT51), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT51), .ZN(new_n1143));
  OAI211_X1 g718(.A(KEYINPUT122), .B(new_n1143), .C1(new_n1047), .C2(new_n1137), .ZN(new_n1144));
  OR2_X1    g719(.A1(new_n1140), .A2(new_n1136), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1134), .B1(new_n1142), .B2(new_n1146), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1138), .A2(KEYINPUT51), .A3(new_n1141), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1148), .A2(KEYINPUT123), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1060), .B1(new_n1133), .B2(new_n1151), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1142), .A2(new_n1134), .A3(new_n1146), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT123), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT62), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT62), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1147), .A2(new_n1156), .A3(new_n1150), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1037), .A2(new_n1130), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1155), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1152), .A2(new_n1159), .ZN(new_n1160));
  XOR2_X1   g735(.A(G290), .B(G1986), .Z(new_n1161));
  NAND2_X1  g736(.A1(new_n966), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(new_n972), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n988), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1163), .ZN(new_n1165));
  AOI211_X1 g740(.A(KEYINPUT127), .B(new_n1165), .C1(new_n1152), .C2(new_n1159), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n987), .B1(new_n1164), .B2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g742(.A(G319), .ZN(new_n1169));
  NOR3_X1   g743(.A1(G401), .A2(G227), .A3(new_n1169), .ZN(new_n1170));
  NAND3_X1  g744(.A1(new_n680), .A2(new_n681), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g745(.A(new_n1171), .B1(new_n880), .B2(new_n882), .ZN(new_n1172));
  NAND2_X1  g746(.A1(new_n1172), .A2(new_n951), .ZN(G225));
  INV_X1    g747(.A(G225), .ZN(G308));
endmodule


