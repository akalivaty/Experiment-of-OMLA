

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589;

  NOR2_X1 U321 ( .A1(n486), .A2(n485), .ZN(n567) );
  NOR2_X1 U322 ( .A1(n491), .A2(n421), .ZN(n422) );
  XNOR2_X1 U323 ( .A(n475), .B(KEYINPUT48), .ZN(n476) );
  XNOR2_X1 U324 ( .A(KEYINPUT38), .B(n460), .ZN(n508) );
  XOR2_X1 U325 ( .A(KEYINPUT28), .B(n482), .Z(n529) );
  XOR2_X1 U326 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n289) );
  XOR2_X1 U327 ( .A(G22GAT), .B(n329), .Z(n290) );
  NOR2_X1 U328 ( .A1(n533), .A2(n360), .ZN(n361) );
  XNOR2_X1 U329 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U330 ( .A(n456), .B(n455), .ZN(n458) );
  XNOR2_X1 U331 ( .A(n477), .B(n476), .ZN(n546) );
  XOR2_X1 U332 ( .A(n439), .B(n438), .Z(n575) );
  XOR2_X1 U333 ( .A(KEYINPUT41), .B(n578), .Z(n554) );
  XOR2_X1 U334 ( .A(n320), .B(n311), .Z(n533) );
  XNOR2_X1 U335 ( .A(KEYINPUT98), .B(n372), .ZN(n547) );
  XNOR2_X1 U336 ( .A(n487), .B(G176GAT), .ZN(n488) );
  XNOR2_X1 U337 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n461) );
  XNOR2_X1 U338 ( .A(n489), .B(n488), .ZN(G1349GAT) );
  XNOR2_X1 U339 ( .A(n462), .B(n461), .ZN(G1330GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT18), .B(KEYINPUT90), .Z(n292) );
  XNOR2_X1 U341 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n291) );
  XNOR2_X1 U342 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U343 ( .A(G169GAT), .B(n293), .Z(n320) );
  XOR2_X1 U344 ( .A(KEYINPUT91), .B(KEYINPUT87), .Z(n295) );
  XNOR2_X1 U345 ( .A(G71GAT), .B(G183GAT), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U347 ( .A(KEYINPUT88), .B(G176GAT), .Z(n297) );
  XNOR2_X1 U348 ( .A(KEYINPUT20), .B(KEYINPUT92), .ZN(n296) );
  XNOR2_X1 U349 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U350 ( .A(n299), .B(n298), .Z(n310) );
  XOR2_X1 U351 ( .A(G120GAT), .B(KEYINPUT89), .Z(n301) );
  XNOR2_X1 U352 ( .A(G15GAT), .B(G113GAT), .ZN(n300) );
  XNOR2_X1 U353 ( .A(n301), .B(n300), .ZN(n308) );
  XOR2_X1 U354 ( .A(KEYINPUT0), .B(G127GAT), .Z(n346) );
  XOR2_X1 U355 ( .A(G134GAT), .B(G190GAT), .Z(n303) );
  XNOR2_X1 U356 ( .A(G43GAT), .B(G99GAT), .ZN(n302) );
  XNOR2_X1 U357 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U358 ( .A(n346), .B(n304), .Z(n306) );
  NAND2_X1 U359 ( .A1(G227GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U360 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U361 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U362 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U363 ( .A(KEYINPUT27), .B(KEYINPUT100), .ZN(n327) );
  XNOR2_X1 U364 ( .A(G8GAT), .B(G183GAT), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n312), .B(KEYINPUT80), .ZN(n401) );
  XOR2_X1 U366 ( .A(G36GAT), .B(G190GAT), .Z(n377) );
  XOR2_X1 U367 ( .A(n401), .B(n377), .Z(n314) );
  NAND2_X1 U368 ( .A1(G226GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U369 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U370 ( .A(n315), .B(KEYINPUT99), .Z(n318) );
  XNOR2_X1 U371 ( .A(G176GAT), .B(G92GAT), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n316), .B(G64GAT), .ZN(n440) );
  XNOR2_X1 U373 ( .A(G204GAT), .B(n440), .ZN(n317) );
  XNOR2_X1 U374 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n326) );
  XNOR2_X1 U376 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n321) );
  XNOR2_X1 U377 ( .A(n321), .B(KEYINPUT93), .ZN(n322) );
  XOR2_X1 U378 ( .A(n322), .B(KEYINPUT94), .Z(n324) );
  XNOR2_X1 U379 ( .A(G197GAT), .B(G218GAT), .ZN(n323) );
  XOR2_X1 U380 ( .A(n324), .B(n323), .Z(n338) );
  INV_X1 U381 ( .A(n338), .ZN(n325) );
  XOR2_X1 U382 ( .A(n326), .B(n325), .Z(n478) );
  INV_X1 U383 ( .A(n478), .ZN(n524) );
  XOR2_X1 U384 ( .A(n327), .B(n524), .Z(n367) );
  XNOR2_X1 U385 ( .A(KEYINPUT23), .B(KEYINPUT96), .ZN(n328) );
  XNOR2_X1 U386 ( .A(n289), .B(n328), .ZN(n329) );
  NAND2_X1 U387 ( .A1(G228GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U388 ( .A(n290), .B(n330), .ZN(n331) );
  XOR2_X1 U389 ( .A(n331), .B(KEYINPUT95), .Z(n336) );
  XOR2_X1 U390 ( .A(KEYINPUT2), .B(G162GAT), .Z(n333) );
  XNOR2_X1 U391 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n332) );
  XNOR2_X1 U392 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U393 ( .A(G141GAT), .B(n334), .Z(n353) );
  XNOR2_X1 U394 ( .A(G50GAT), .B(n353), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U396 ( .A(n338), .B(n337), .Z(n343) );
  XOR2_X1 U397 ( .A(KEYINPUT72), .B(KEYINPUT71), .Z(n340) );
  XNOR2_X1 U398 ( .A(G78GAT), .B(G148GAT), .ZN(n339) );
  XNOR2_X1 U399 ( .A(n340), .B(n339), .ZN(n342) );
  XOR2_X1 U400 ( .A(G106GAT), .B(G204GAT), .Z(n341) );
  XNOR2_X1 U401 ( .A(n342), .B(n341), .ZN(n457) );
  XNOR2_X1 U402 ( .A(n343), .B(n457), .ZN(n482) );
  INV_X1 U403 ( .A(n529), .ZN(n358) );
  XOR2_X1 U404 ( .A(KEYINPUT97), .B(KEYINPUT6), .Z(n345) );
  XNOR2_X1 U405 ( .A(G148GAT), .B(G85GAT), .ZN(n344) );
  XNOR2_X1 U406 ( .A(n345), .B(n344), .ZN(n357) );
  XOR2_X1 U407 ( .A(G120GAT), .B(G57GAT), .Z(n447) );
  XOR2_X1 U408 ( .A(G29GAT), .B(G134GAT), .Z(n382) );
  XOR2_X1 U409 ( .A(n447), .B(n382), .Z(n348) );
  XOR2_X1 U410 ( .A(G113GAT), .B(G1GAT), .Z(n430) );
  XNOR2_X1 U411 ( .A(n430), .B(n346), .ZN(n347) );
  XNOR2_X1 U412 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U413 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n350) );
  NAND2_X1 U414 ( .A1(G225GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U415 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U416 ( .A(n352), .B(n351), .Z(n355) );
  XNOR2_X1 U417 ( .A(n353), .B(KEYINPUT5), .ZN(n354) );
  XNOR2_X1 U418 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U419 ( .A(n357), .B(n356), .Z(n372) );
  NAND2_X1 U420 ( .A1(n358), .A2(n547), .ZN(n359) );
  NOR2_X1 U421 ( .A1(n367), .A2(n359), .ZN(n532) );
  XNOR2_X1 U422 ( .A(KEYINPUT101), .B(n532), .ZN(n360) );
  XNOR2_X1 U423 ( .A(n361), .B(KEYINPUT102), .ZN(n374) );
  NAND2_X1 U424 ( .A1(n533), .A2(n524), .ZN(n362) );
  NAND2_X1 U425 ( .A1(n482), .A2(n362), .ZN(n363) );
  XNOR2_X1 U426 ( .A(KEYINPUT25), .B(n363), .ZN(n370) );
  NOR2_X1 U427 ( .A1(n533), .A2(n482), .ZN(n365) );
  XNOR2_X1 U428 ( .A(KEYINPUT104), .B(KEYINPUT26), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U430 ( .A(KEYINPUT103), .B(n366), .Z(n573) );
  INV_X1 U431 ( .A(n367), .ZN(n368) );
  NAND2_X1 U432 ( .A1(n573), .A2(n368), .ZN(n545) );
  XNOR2_X1 U433 ( .A(KEYINPUT105), .B(n545), .ZN(n369) );
  NOR2_X1 U434 ( .A1(n370), .A2(n369), .ZN(n371) );
  NOR2_X1 U435 ( .A1(n372), .A2(n371), .ZN(n373) );
  NOR2_X1 U436 ( .A1(n374), .A2(n373), .ZN(n491) );
  INV_X1 U437 ( .A(KEYINPUT36), .ZN(n395) );
  XOR2_X1 U438 ( .A(KEYINPUT76), .B(KEYINPUT10), .Z(n376) );
  XNOR2_X1 U439 ( .A(G106GAT), .B(KEYINPUT77), .ZN(n375) );
  XNOR2_X1 U440 ( .A(n376), .B(n375), .ZN(n394) );
  XOR2_X1 U441 ( .A(n377), .B(KEYINPUT78), .Z(n379) );
  NAND2_X1 U442 ( .A1(G232GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U443 ( .A(n379), .B(n378), .ZN(n387) );
  XOR2_X1 U444 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n381) );
  XNOR2_X1 U445 ( .A(G92GAT), .B(KEYINPUT79), .ZN(n380) );
  XNOR2_X1 U446 ( .A(n381), .B(n380), .ZN(n383) );
  XNOR2_X1 U447 ( .A(n383), .B(n382), .ZN(n385) );
  XOR2_X1 U448 ( .A(G218GAT), .B(G162GAT), .Z(n384) );
  XNOR2_X1 U449 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U450 ( .A(n387), .B(n386), .Z(n392) );
  XOR2_X1 U451 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n389) );
  XNOR2_X1 U452 ( .A(G50GAT), .B(G43GAT), .ZN(n388) );
  XNOR2_X1 U453 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U454 ( .A(KEYINPUT7), .B(n390), .Z(n427) );
  XOR2_X1 U455 ( .A(G99GAT), .B(G85GAT), .Z(n449) );
  XNOR2_X1 U456 ( .A(n427), .B(n449), .ZN(n391) );
  XNOR2_X1 U457 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U458 ( .A(n394), .B(n393), .Z(n560) );
  NAND2_X1 U459 ( .A1(n395), .A2(n560), .ZN(n398) );
  INV_X1 U460 ( .A(n560), .ZN(n396) );
  NAND2_X1 U461 ( .A1(KEYINPUT36), .A2(n396), .ZN(n397) );
  NAND2_X1 U462 ( .A1(n398), .A2(n397), .ZN(n467) );
  XOR2_X1 U463 ( .A(KEYINPUT13), .B(KEYINPUT69), .Z(n400) );
  XNOR2_X1 U464 ( .A(G71GAT), .B(KEYINPUT70), .ZN(n399) );
  XNOR2_X1 U465 ( .A(n400), .B(n399), .ZN(n450) );
  XNOR2_X1 U466 ( .A(n450), .B(n401), .ZN(n420) );
  XOR2_X1 U467 ( .A(KEYINPUT14), .B(G64GAT), .Z(n403) );
  XNOR2_X1 U468 ( .A(G1GAT), .B(G57GAT), .ZN(n402) );
  XNOR2_X1 U469 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U470 ( .A(KEYINPUT86), .B(KEYINPUT15), .Z(n405) );
  XNOR2_X1 U471 ( .A(KEYINPUT12), .B(KEYINPUT81), .ZN(n404) );
  XNOR2_X1 U472 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U473 ( .A(n407), .B(n406), .Z(n418) );
  XOR2_X1 U474 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n409) );
  XNOR2_X1 U475 ( .A(KEYINPUT83), .B(KEYINPUT82), .ZN(n408) );
  XNOR2_X1 U476 ( .A(n409), .B(n408), .ZN(n416) );
  XOR2_X1 U477 ( .A(G15GAT), .B(G22GAT), .Z(n431) );
  XOR2_X1 U478 ( .A(G155GAT), .B(G78GAT), .Z(n411) );
  XNOR2_X1 U479 ( .A(G127GAT), .B(G211GAT), .ZN(n410) );
  XNOR2_X1 U480 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U481 ( .A(n431), .B(n412), .Z(n414) );
  NAND2_X1 U482 ( .A1(G231GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U483 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U484 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U485 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U486 ( .A(n420), .B(n419), .Z(n565) );
  INV_X1 U487 ( .A(n565), .ZN(n583) );
  NAND2_X1 U488 ( .A1(n467), .A2(n583), .ZN(n421) );
  XNOR2_X1 U489 ( .A(n422), .B(KEYINPUT108), .ZN(n423) );
  XNOR2_X1 U490 ( .A(n423), .B(KEYINPUT37), .ZN(n521) );
  XOR2_X1 U491 ( .A(G8GAT), .B(G141GAT), .Z(n425) );
  XNOR2_X1 U492 ( .A(G169GAT), .B(G197GAT), .ZN(n424) );
  XNOR2_X1 U493 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U494 ( .A(n427), .B(n426), .ZN(n439) );
  XOR2_X1 U495 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n429) );
  XNOR2_X1 U496 ( .A(KEYINPUT67), .B(KEYINPUT30), .ZN(n428) );
  XNOR2_X1 U497 ( .A(n429), .B(n428), .ZN(n435) );
  XOR2_X1 U498 ( .A(G29GAT), .B(G36GAT), .Z(n433) );
  XNOR2_X1 U499 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U500 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U501 ( .A(n435), .B(n434), .Z(n437) );
  NAND2_X1 U502 ( .A1(G229GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U503 ( .A(n437), .B(n436), .ZN(n438) );
  NAND2_X1 U504 ( .A1(n440), .A2(KEYINPUT32), .ZN(n444) );
  INV_X1 U505 ( .A(n440), .ZN(n442) );
  INV_X1 U506 ( .A(KEYINPUT32), .ZN(n441) );
  NAND2_X1 U507 ( .A1(n442), .A2(n441), .ZN(n443) );
  NAND2_X1 U508 ( .A1(n444), .A2(n443), .ZN(n446) );
  AND2_X1 U509 ( .A1(G230GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U510 ( .A(n446), .B(n445), .ZN(n448) );
  XNOR2_X1 U511 ( .A(n448), .B(n447), .ZN(n456) );
  XOR2_X1 U512 ( .A(n450), .B(n449), .Z(n454) );
  XOR2_X1 U513 ( .A(KEYINPUT73), .B(KEYINPUT31), .Z(n452) );
  XNOR2_X1 U514 ( .A(KEYINPUT33), .B(KEYINPUT74), .ZN(n451) );
  XNOR2_X1 U515 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U516 ( .A(n458), .B(n457), .Z(n578) );
  NOR2_X1 U517 ( .A1(n575), .A2(n578), .ZN(n459) );
  XNOR2_X1 U518 ( .A(n459), .B(KEYINPUT75), .ZN(n494) );
  NOR2_X1 U519 ( .A1(n521), .A2(n494), .ZN(n460) );
  NAND2_X1 U520 ( .A1(n508), .A2(n533), .ZN(n462) );
  INV_X1 U521 ( .A(KEYINPUT54), .ZN(n480) );
  INV_X1 U522 ( .A(n575), .ZN(n563) );
  NAND2_X1 U523 ( .A1(n563), .A2(n554), .ZN(n463) );
  XNOR2_X1 U524 ( .A(n463), .B(KEYINPUT46), .ZN(n465) );
  NOR2_X1 U525 ( .A1(n396), .A2(n565), .ZN(n464) );
  AND2_X1 U526 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U527 ( .A(KEYINPUT47), .B(n466), .ZN(n474) );
  NAND2_X1 U528 ( .A1(n467), .A2(n565), .ZN(n468) );
  XNOR2_X1 U529 ( .A(n468), .B(KEYINPUT45), .ZN(n469) );
  XOR2_X1 U530 ( .A(KEYINPUT65), .B(n469), .Z(n470) );
  NOR2_X1 U531 ( .A1(n578), .A2(n470), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n471), .B(KEYINPUT114), .ZN(n472) );
  NAND2_X1 U533 ( .A1(n472), .A2(n575), .ZN(n473) );
  NAND2_X1 U534 ( .A1(n474), .A2(n473), .ZN(n477) );
  XNOR2_X1 U535 ( .A(KEYINPUT64), .B(KEYINPUT115), .ZN(n475) );
  NOR2_X1 U536 ( .A1(n546), .A2(n478), .ZN(n479) );
  XNOR2_X1 U537 ( .A(n480), .B(n479), .ZN(n481) );
  NOR2_X1 U538 ( .A1(n547), .A2(n481), .ZN(n574) );
  NAND2_X1 U539 ( .A1(n574), .A2(n482), .ZN(n484) );
  XOR2_X1 U540 ( .A(KEYINPUT122), .B(KEYINPUT55), .Z(n483) );
  XNOR2_X1 U541 ( .A(n484), .B(n483), .ZN(n486) );
  INV_X1 U542 ( .A(n533), .ZN(n485) );
  NAND2_X1 U543 ( .A1(n567), .A2(n554), .ZN(n489) );
  XOR2_X1 U544 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n487) );
  NOR2_X1 U545 ( .A1(n583), .A2(n396), .ZN(n490) );
  XNOR2_X1 U546 ( .A(n490), .B(KEYINPUT16), .ZN(n493) );
  INV_X1 U547 ( .A(n491), .ZN(n492) );
  NAND2_X1 U548 ( .A1(n493), .A2(n492), .ZN(n510) );
  NOR2_X1 U549 ( .A1(n494), .A2(n510), .ZN(n501) );
  NAND2_X1 U550 ( .A1(n547), .A2(n501), .ZN(n495) );
  XNOR2_X1 U551 ( .A(n495), .B(KEYINPUT34), .ZN(n496) );
  XNOR2_X1 U552 ( .A(G1GAT), .B(n496), .ZN(G1324GAT) );
  NAND2_X1 U553 ( .A1(n501), .A2(n524), .ZN(n497) );
  XNOR2_X1 U554 ( .A(n497), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT35), .B(KEYINPUT106), .Z(n499) );
  NAND2_X1 U556 ( .A1(n501), .A2(n533), .ZN(n498) );
  XNOR2_X1 U557 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U558 ( .A(G15GAT), .B(n500), .ZN(G1326GAT) );
  XOR2_X1 U559 ( .A(G22GAT), .B(KEYINPUT107), .Z(n503) );
  NAND2_X1 U560 ( .A1(n501), .A2(n529), .ZN(n502) );
  XNOR2_X1 U561 ( .A(n503), .B(n502), .ZN(G1327GAT) );
  XOR2_X1 U562 ( .A(G29GAT), .B(KEYINPUT39), .Z(n505) );
  NAND2_X1 U563 ( .A1(n508), .A2(n547), .ZN(n504) );
  XNOR2_X1 U564 ( .A(n505), .B(n504), .ZN(G1328GAT) );
  XOR2_X1 U565 ( .A(G36GAT), .B(KEYINPUT109), .Z(n507) );
  NAND2_X1 U566 ( .A1(n524), .A2(n508), .ZN(n506) );
  XNOR2_X1 U567 ( .A(n507), .B(n506), .ZN(G1329GAT) );
  NAND2_X1 U568 ( .A1(n508), .A2(n529), .ZN(n509) );
  XNOR2_X1 U569 ( .A(n509), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT42), .B(KEYINPUT110), .Z(n512) );
  NAND2_X1 U571 ( .A1(n554), .A2(n575), .ZN(n520) );
  NOR2_X1 U572 ( .A1(n520), .A2(n510), .ZN(n517) );
  NAND2_X1 U573 ( .A1(n517), .A2(n547), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U575 ( .A(G57GAT), .B(n513), .Z(G1332GAT) );
  XOR2_X1 U576 ( .A(G64GAT), .B(KEYINPUT111), .Z(n515) );
  NAND2_X1 U577 ( .A1(n517), .A2(n524), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n515), .B(n514), .ZN(G1333GAT) );
  NAND2_X1 U579 ( .A1(n517), .A2(n533), .ZN(n516) );
  XNOR2_X1 U580 ( .A(n516), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U581 ( .A(G78GAT), .B(KEYINPUT43), .Z(n519) );
  NAND2_X1 U582 ( .A1(n517), .A2(n529), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  XNOR2_X1 U584 ( .A(G85GAT), .B(KEYINPUT112), .ZN(n523) );
  NOR2_X1 U585 ( .A1(n521), .A2(n520), .ZN(n528) );
  NAND2_X1 U586 ( .A1(n528), .A2(n547), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n523), .B(n522), .ZN(G1336GAT) );
  NAND2_X1 U588 ( .A1(n528), .A2(n524), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n525), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U590 ( .A(G99GAT), .B(KEYINPUT113), .Z(n527) );
  NAND2_X1 U591 ( .A1(n528), .A2(n533), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(G1338GAT) );
  NAND2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n530), .B(KEYINPUT44), .ZN(n531) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  NAND2_X1 U596 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U597 ( .A1(n546), .A2(n534), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n541), .A2(n563), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n535), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .Z(n537) );
  NAND2_X1 U601 ( .A1(n541), .A2(n554), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n539) );
  NAND2_X1 U604 ( .A1(n541), .A2(n565), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U606 ( .A(G127GAT), .B(n540), .Z(G1342GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U608 ( .A1(n541), .A2(n396), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U610 ( .A(G134GAT), .B(n544), .Z(G1343GAT) );
  NOR2_X1 U611 ( .A1(n546), .A2(n545), .ZN(n548) );
  NAND2_X1 U612 ( .A1(n548), .A2(n547), .ZN(n559) );
  NOR2_X1 U613 ( .A1(n575), .A2(n559), .ZN(n550) );
  XNOR2_X1 U614 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U616 ( .A(G141GAT), .B(n551), .ZN(G1344GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT120), .B(KEYINPUT52), .Z(n553) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(n557) );
  INV_X1 U620 ( .A(n554), .ZN(n555) );
  NOR2_X1 U621 ( .A1(n555), .A2(n559), .ZN(n556) );
  XOR2_X1 U622 ( .A(n557), .B(n556), .Z(G1345GAT) );
  NOR2_X1 U623 ( .A1(n583), .A2(n559), .ZN(n558) );
  XOR2_X1 U624 ( .A(G155GAT), .B(n558), .Z(G1346GAT) );
  NOR2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n562) );
  XNOR2_X1 U626 ( .A(G162GAT), .B(KEYINPUT121), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n563), .A2(n567), .ZN(n564) );
  XNOR2_X1 U629 ( .A(G169GAT), .B(n564), .ZN(G1348GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n567), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U632 ( .A1(n567), .A2(n396), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n570), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT124), .B(KEYINPUT59), .Z(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n577) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n582) );
  NOR2_X1 U640 ( .A1(n575), .A2(n582), .ZN(n576) );
  XOR2_X1 U641 ( .A(n577), .B(n576), .Z(G1352GAT) );
  INV_X1 U642 ( .A(n582), .ZN(n585) );
  AND2_X1 U643 ( .A1(n578), .A2(n585), .ZN(n580) );
  XNOR2_X1 U644 ( .A(KEYINPUT125), .B(KEYINPUT61), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U646 ( .A(G204GAT), .B(n581), .Z(G1353GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(G211GAT), .B(n584), .Z(G1354GAT) );
  NAND2_X1 U649 ( .A1(n585), .A2(n467), .ZN(n586) );
  XNOR2_X1 U650 ( .A(n586), .B(KEYINPUT62), .ZN(n587) );
  XOR2_X1 U651 ( .A(n587), .B(KEYINPUT126), .Z(n589) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(G1355GAT) );
endmodule

