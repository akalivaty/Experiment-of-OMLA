//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 0 0 0 0 0 0 1 1 1 0 0 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n997, new_n998;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT26), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  AOI22_X1  g004(.A1(new_n205), .A2(KEYINPUT68), .B1(G183gat), .B2(G190gat), .ZN(new_n206));
  OR2_X1    g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT26), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT68), .ZN(new_n209));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  NAND4_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n204), .A4(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n206), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT69), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT69), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n206), .A2(new_n214), .A3(new_n211), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT67), .ZN(new_n218));
  INV_X1    g017(.A(G183gat), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT27), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n219), .A2(KEYINPUT27), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n217), .B(new_n220), .C1(new_n221), .C2(new_n218), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT28), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT27), .B(G183gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(KEYINPUT28), .A3(new_n217), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n216), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n202), .A2(KEYINPUT23), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT64), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n210), .A2(KEYINPUT23), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(new_n207), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(G183gat), .B2(G190gat), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n230), .B(new_n232), .C1(new_n233), .C2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT25), .ZN(new_n237));
  OAI22_X1  g036(.A1(new_n219), .A2(new_n217), .B1(KEYINPUT65), .B2(KEYINPUT24), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n238), .B1(KEYINPUT65), .B2(KEYINPUT24), .ZN(new_n239));
  OR2_X1    g038(.A1(new_n239), .A2(new_n235), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n232), .A2(KEYINPUT25), .A3(new_n229), .ZN(new_n241));
  AOI22_X1  g040(.A1(new_n236), .A2(new_n237), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n242), .A2(KEYINPUT66), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n236), .A2(new_n237), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n240), .A2(new_n241), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n244), .A2(KEYINPUT66), .A3(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n228), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G113gat), .B(G120gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT70), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT1), .ZN(new_n251));
  XNOR2_X1  g050(.A(G127gat), .B(G134gat), .ZN(new_n252));
  INV_X1    g051(.A(G113gat), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n253), .A2(KEYINPUT70), .A3(G120gat), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n250), .A2(new_n251), .A3(new_n252), .A4(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n252), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n256), .B1(KEYINPUT1), .B2(new_n248), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n247), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(G227gat), .ZN(new_n261));
  INV_X1    g060(.A(G233gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n258), .B(new_n228), .C1(new_n243), .C2(new_n246), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n260), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT32), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT33), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  XOR2_X1   g067(.A(G15gat), .B(G43gat), .Z(new_n269));
  XNOR2_X1  g068(.A(G71gat), .B(G99gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n266), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n271), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n265), .B(KEYINPUT32), .C1(new_n267), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n263), .B1(new_n260), .B2(new_n264), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT34), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n279), .B1(new_n276), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n260), .A2(new_n264), .ZN(new_n283));
  INV_X1    g082(.A(new_n263), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n280), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n285), .B1(new_n276), .B2(new_n278), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n286), .A2(new_n272), .A3(new_n274), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n288));
  INV_X1    g087(.A(G22gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(G197gat), .A2(G204gat), .ZN(new_n292));
  AND2_X1   g091(.A1(G197gat), .A2(G204gat), .ZN(new_n293));
  AND2_X1   g092(.A1(G211gat), .A2(G218gat), .ZN(new_n294));
  OAI22_X1  g093(.A1(new_n292), .A2(new_n293), .B1(new_n294), .B2(KEYINPUT22), .ZN(new_n295));
  XOR2_X1   g094(.A(G211gat), .B(G218gat), .Z(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  XOR2_X1   g096(.A(G155gat), .B(G162gat), .Z(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G155gat), .ZN(new_n300));
  INV_X1    g099(.A(G162gat), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT2), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  XOR2_X1   g101(.A(G141gat), .B(G148gat), .Z(new_n303));
  NAND3_X1  g102(.A1(new_n299), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n302), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(new_n298), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT3), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT29), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n297), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n312), .B1(G228gat), .B2(G233gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT84), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n297), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n295), .A2(new_n314), .A3(new_n296), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(new_n311), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n309), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  AND3_X1   g117(.A1(new_n304), .A2(new_n306), .A3(KEYINPUT77), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT77), .B1(new_n304), .B2(new_n306), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT85), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT85), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n318), .A2(new_n324), .A3(new_n321), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n313), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT3), .B1(new_n297), .B2(new_n311), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n327), .A2(new_n308), .ZN(new_n328));
  OAI211_X1 g127(.A(G228gat), .B(G233gat), .C1(new_n312), .C2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G78gat), .B(G106gat), .ZN(new_n330));
  INV_X1    g129(.A(G50gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(KEYINPUT83), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n326), .A2(new_n329), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n334), .B1(new_n326), .B2(new_n329), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n291), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n326), .A2(new_n329), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(new_n333), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n326), .A2(new_n329), .A3(new_n334), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(new_n290), .A3(new_n340), .ZN(new_n341));
  AND2_X1   g140(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n282), .A2(new_n287), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT88), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G1gat), .B(G29gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n346), .B(KEYINPUT0), .ZN(new_n347));
  XNOR2_X1  g146(.A(G57gat), .B(G85gat), .ZN(new_n348));
  XOR2_X1   g147(.A(new_n347), .B(new_n348), .Z(new_n349));
  NAND2_X1  g148(.A1(new_n307), .A2(KEYINPUT3), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n310), .A2(new_n258), .A3(new_n350), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n259), .B(KEYINPUT4), .C1(new_n319), .C2(new_n320), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n306), .A2(new_n304), .A3(new_n255), .A4(new_n257), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT4), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT5), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n351), .A2(new_n352), .A3(new_n355), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n307), .A2(new_n258), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n361), .A2(KEYINPUT78), .A3(new_n353), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT78), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n307), .A2(new_n258), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n358), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n360), .B1(new_n365), .B2(new_n356), .ZN(new_n366));
  INV_X1    g165(.A(new_n353), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT79), .B1(new_n367), .B2(new_n354), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n259), .B(new_n354), .C1(new_n319), .C2(new_n320), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT79), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n353), .A2(new_n370), .A3(KEYINPUT4), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n368), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT5), .B1(new_n372), .B2(new_n351), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n349), .B1(new_n366), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT80), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT6), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT80), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n377), .B(new_n349), .C1(new_n366), .C2(new_n373), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT81), .ZN(new_n380));
  OR2_X1    g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NOR3_X1   g180(.A1(new_n366), .A2(new_n373), .A3(new_n349), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n382), .B1(new_n379), .B2(new_n380), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(KEYINPUT6), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n297), .ZN(new_n387));
  AND2_X1   g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n388), .B(new_n228), .C1(new_n243), .C2(new_n246), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n244), .A2(new_n245), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT73), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n228), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n213), .A2(new_n215), .B1(new_n224), .B2(new_n226), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT73), .B1(new_n393), .B2(new_n242), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n388), .A2(KEYINPUT29), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n392), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n387), .B1(new_n389), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n392), .A2(new_n394), .ZN(new_n398));
  AOI22_X1  g197(.A1(new_n395), .A2(new_n247), .B1(new_n398), .B2(new_n388), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n397), .B1(new_n399), .B2(new_n387), .ZN(new_n400));
  XOR2_X1   g199(.A(G8gat), .B(G36gat), .Z(new_n401));
  XNOR2_X1  g200(.A(G64gat), .B(G92gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n404));
  XOR2_X1   g203(.A(new_n403), .B(new_n404), .Z(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n400), .A2(KEYINPUT30), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT76), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n247), .A2(new_n395), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n398), .A2(new_n388), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n410), .A3(new_n387), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n405), .B1(new_n412), .B2(new_n397), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n407), .A2(new_n408), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT30), .ZN(new_n415));
  INV_X1    g214(.A(new_n400), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n415), .B1(new_n416), .B2(new_n405), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n408), .B1(new_n407), .B2(new_n413), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n282), .A2(new_n287), .A3(new_n342), .A4(KEYINPUT88), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n345), .A2(new_n386), .A3(new_n420), .A4(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT35), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n417), .A2(new_n413), .A3(new_n407), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n282), .A2(new_n287), .A3(KEYINPUT72), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT72), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n286), .A2(new_n426), .A3(new_n272), .A4(new_n274), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n424), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n382), .ZN(new_n429));
  MUX2_X1   g228(.A(new_n376), .B(new_n379), .S(new_n429), .Z(new_n430));
  NAND2_X1  g229(.A1(new_n337), .A2(new_n341), .ZN(new_n431));
  NOR3_X1   g230(.A1(new_n430), .A2(KEYINPUT35), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT36), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n425), .A2(new_n434), .A3(new_n427), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n282), .A2(new_n287), .A3(KEYINPUT36), .ZN(new_n436));
  XNOR2_X1  g235(.A(KEYINPUT86), .B(KEYINPUT38), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n389), .A2(new_n396), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n297), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT37), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(new_n411), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n405), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n441), .B1(new_n440), .B2(new_n411), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n438), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT87), .ZN(new_n446));
  INV_X1    g245(.A(new_n443), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n441), .B1(new_n399), .B2(new_n297), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n439), .A2(new_n387), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n438), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n447), .A2(new_n450), .B1(new_n400), .B2(new_n406), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT87), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n452), .B(new_n438), .C1(new_n443), .C2(new_n444), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n446), .A2(new_n430), .A3(new_n451), .A4(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT40), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n356), .B1(new_n372), .B2(new_n351), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT39), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n349), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n362), .A2(new_n364), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT39), .B1(new_n461), .B2(new_n357), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n455), .B1(new_n459), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n429), .ZN(new_n465));
  NOR3_X1   g264(.A1(new_n459), .A2(new_n455), .A3(new_n463), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n431), .B1(new_n424), .B2(new_n467), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n435), .A2(new_n436), .B1(new_n454), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n419), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n470), .A2(new_n417), .A3(new_n414), .ZN(new_n471));
  AOI22_X1  g270(.A1(new_n381), .A2(new_n383), .B1(KEYINPUT6), .B2(new_n382), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n431), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n423), .A2(new_n433), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n289), .A2(G15gat), .ZN(new_n475));
  INV_X1    g274(.A(G15gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(G22gat), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT91), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n475), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(G1gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(G15gat), .B(G22gat), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n482), .A2(new_n478), .A3(G1gat), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT16), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(G8gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT92), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT92), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n486), .A2(new_n489), .A3(G8gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(G8gat), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n481), .A2(new_n483), .A3(new_n492), .A4(new_n485), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(KEYINPUT93), .ZN(new_n494));
  NAND2_X1  g293(.A1(KEYINPUT90), .A2(G36gat), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(KEYINPUT90), .A2(G36gat), .ZN(new_n497));
  OAI21_X1  g296(.A(G29gat), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT14), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n499), .B1(G29gat), .B2(G36gat), .ZN(new_n500));
  INV_X1    g299(.A(G29gat), .ZN(new_n501));
  INV_X1    g300(.A(G36gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT14), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n498), .A2(KEYINPUT15), .A3(new_n500), .A4(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G43gat), .B(G50gat), .ZN(new_n505));
  OR2_X1    g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT15), .ZN(new_n507));
  INV_X1    g306(.A(new_n497), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n501), .B1(new_n508), .B2(new_n495), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n503), .A2(new_n500), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n511), .A2(new_n504), .A3(new_n505), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT17), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n506), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n513), .B1(new_n506), .B2(new_n512), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n491), .B(new_n494), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n506), .A2(new_n512), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n486), .A2(new_n489), .A3(G8gat), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n489), .B1(new_n486), .B2(G8gat), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT93), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n493), .B(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n517), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(G229gat), .A2(G233gat), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n524), .B(KEYINPUT94), .Z(new_n525));
  NAND3_X1  g324(.A1(new_n516), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT18), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n516), .A2(new_n523), .A3(KEYINPUT18), .A4(new_n525), .ZN(new_n529));
  INV_X1    g328(.A(new_n517), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n491), .A2(new_n530), .A3(new_n494), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n523), .A2(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n525), .B(KEYINPUT13), .Z(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n528), .A2(new_n529), .A3(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G113gat), .B(G141gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  XOR2_X1   g337(.A(G169gat), .B(G197gat), .Z(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT12), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n535), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n528), .A2(new_n529), .A3(new_n534), .A4(new_n541), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n545), .B(KEYINPUT95), .Z(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n474), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT98), .ZN(new_n549));
  NAND2_X1  g348(.A1(G71gat), .A2(G78gat), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT9), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OR2_X1    g351(.A1(G57gat), .A2(G64gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(G57gat), .A2(G64gat), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT96), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n553), .A2(new_n556), .A3(new_n554), .ZN(new_n557));
  XNOR2_X1  g356(.A(G71gat), .B(G78gat), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n555), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AND2_X1   g358(.A1(G57gat), .A2(G64gat), .ZN(new_n560));
  NOR2_X1   g359(.A1(G57gat), .A2(G64gat), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g361(.A1(G71gat), .A2(G78gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(G71gat), .A2(G78gat), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n552), .B(new_n562), .C1(new_n565), .C2(new_n556), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n559), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n567), .A2(KEYINPUT21), .ZN(new_n568));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G127gat), .ZN(new_n571));
  AOI211_X1 g370(.A(new_n522), .B(new_n520), .C1(KEYINPUT21), .C2(new_n567), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(new_n300), .ZN(new_n575));
  XOR2_X1   g374(.A(G183gat), .B(G211gat), .Z(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n573), .B(new_n577), .Z(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G99gat), .A2(G106gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT8), .ZN(new_n581));
  NAND2_X1  g380(.A1(G85gat), .A2(G92gat), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT7), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(G85gat), .ZN(new_n585));
  INV_X1    g384(.A(G92gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n581), .A2(new_n584), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G99gat), .B(G106gat), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  AND3_X1   g391(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI22_X1  g394(.A1(KEYINPUT8), .A2(new_n580), .B1(new_n585), .B2(new_n586), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n590), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT41), .ZN(new_n600));
  NAND2_X1  g399(.A1(G232gat), .A2(G233gat), .ZN(new_n601));
  OAI22_X1  g400(.A1(new_n530), .A2(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n514), .A2(new_n515), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n602), .B1(new_n603), .B2(new_n599), .ZN(new_n604));
  XOR2_X1   g403(.A(G190gat), .B(G218gat), .Z(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n601), .A2(new_n600), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT97), .ZN(new_n608));
  XOR2_X1   g407(.A(G134gat), .B(G162gat), .Z(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n606), .B(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n549), .B1(new_n579), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n611), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n578), .A2(KEYINPUT98), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G230gat), .A2(G233gat), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n595), .A2(new_n590), .A3(new_n596), .ZN(new_n616));
  INV_X1    g415(.A(new_n597), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n567), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT10), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n566), .B(new_n559), .C1(new_n592), .C2(new_n597), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n621), .A2(KEYINPUT99), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT99), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n618), .A2(new_n620), .A3(new_n623), .A4(new_n619), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n598), .A2(KEYINPUT10), .A3(new_n567), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n615), .B1(new_n622), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n618), .A2(new_n620), .ZN(new_n629));
  INV_X1    g428(.A(new_n615), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(KEYINPUT100), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT100), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n629), .A2(new_n633), .A3(new_n630), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G120gat), .B(G148gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(G176gat), .B(G204gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n636), .B(new_n637), .Z(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NOR3_X1   g438(.A1(new_n628), .A2(new_n635), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n635), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n621), .A2(KEYINPUT99), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n642), .A2(new_n625), .A3(new_n624), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n643), .A2(KEYINPUT101), .A3(new_n615), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT101), .B1(new_n643), .B2(new_n615), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n641), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n640), .B1(new_n646), .B2(new_n639), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n612), .A2(new_n614), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n386), .B(KEYINPUT102), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n548), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g451(.A1(new_n548), .A2(new_n649), .ZN(new_n653));
  INV_X1    g452(.A(new_n424), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n655), .A2(new_n492), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n656), .A2(KEYINPUT103), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(KEYINPUT103), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT42), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT16), .B(G8gat), .Z(new_n660));
  AOI21_X1  g459(.A(new_n659), .B1(new_n655), .B2(new_n660), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n655), .A2(new_n659), .A3(new_n660), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n657), .B(new_n658), .C1(new_n661), .C2(new_n662), .ZN(G1325gat));
  NAND2_X1  g462(.A1(new_n435), .A2(new_n436), .ZN(new_n664));
  OAI21_X1  g463(.A(G15gat), .B1(new_n653), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n425), .A2(new_n427), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n548), .A2(new_n476), .A3(new_n666), .A4(new_n649), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(G1326gat));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n342), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT43), .B(G22gat), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  INV_X1    g470(.A(KEYINPUT45), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n579), .A2(new_n647), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n613), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n548), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n650), .A2(new_n501), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n672), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  OR3_X1    g476(.A1(new_n675), .A2(new_n672), .A3(new_n676), .ZN(new_n678));
  INV_X1    g477(.A(new_n545), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n681), .B1(new_n474), .B2(new_n613), .ZN(new_n682));
  NAND2_X1  g481(.A1(KEYINPUT104), .A2(KEYINPUT44), .ZN(new_n683));
  AOI22_X1  g482(.A1(new_n422), .A2(KEYINPUT35), .B1(new_n428), .B2(new_n432), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n454), .A2(new_n468), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n664), .A2(new_n473), .A3(new_n685), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n611), .B(new_n683), .C1(new_n684), .C2(new_n686), .ZN(new_n687));
  AOI211_X1 g486(.A(new_n679), .B(new_n673), .C1(new_n682), .C2(new_n687), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n688), .A2(new_n650), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n677), .B(new_n678), .C1(new_n689), .C2(new_n501), .ZN(G1328gat));
  NAND2_X1  g489(.A1(new_n508), .A2(new_n495), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n654), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT46), .B1(new_n675), .B2(new_n693), .ZN(new_n694));
  OR3_X1    g493(.A1(new_n675), .A2(KEYINPUT46), .A3(new_n693), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n688), .A2(new_n424), .ZN(new_n696));
  INV_X1    g495(.A(new_n691), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n694), .B(new_n695), .C1(new_n696), .C2(new_n697), .ZN(G1329gat));
  INV_X1    g497(.A(G43gat), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n548), .A2(new_n699), .A3(new_n666), .A4(new_n674), .ZN(new_n700));
  INV_X1    g499(.A(new_n664), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n688), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n700), .B1(new_n702), .B2(new_n699), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT47), .B1(new_n700), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  OAI221_X1 g505(.A(new_n700), .B1(new_n704), .B2(KEYINPUT47), .C1(new_n702), .C2(new_n699), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(G1330gat));
  AOI21_X1  g507(.A(new_n331), .B1(new_n688), .B2(new_n431), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT48), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n675), .A2(G50gat), .A3(new_n342), .ZN(new_n711));
  OR3_X1    g510(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n710), .B1(new_n709), .B2(new_n711), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(G1331gat));
  INV_X1    g513(.A(new_n474), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n646), .A2(new_n639), .ZN(new_n716));
  INV_X1    g515(.A(new_n640), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AND4_X1   g517(.A1(new_n679), .A2(new_n612), .A3(new_n614), .A4(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n650), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g522(.A1(new_n720), .A2(new_n654), .ZN(new_n724));
  NOR2_X1   g523(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n725));
  AND2_X1   g524(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(new_n724), .B2(new_n725), .ZN(G1333gat));
  OAI21_X1  g527(.A(G71gat), .B1(new_n720), .B2(new_n664), .ZN(new_n729));
  INV_X1    g528(.A(G71gat), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n666), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n720), .B2(new_n731), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g532(.A1(new_n721), .A2(new_n431), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g534(.A1(new_n474), .A2(new_n613), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n578), .A2(new_n545), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n736), .A2(KEYINPUT106), .A3(KEYINPUT51), .A4(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT106), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n611), .B(new_n737), .C1(new_n684), .C2(new_n686), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT51), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n740), .A2(new_n741), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n650), .A2(new_n585), .A3(new_n718), .ZN(new_n746));
  INV_X1    g545(.A(new_n737), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n747), .A2(new_n647), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n749), .B1(new_n682), .B2(new_n687), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n750), .A2(new_n650), .ZN(new_n751));
  OAI22_X1  g550(.A1(new_n745), .A2(new_n746), .B1(new_n585), .B2(new_n751), .ZN(G1336gat));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753));
  AOI211_X1 g552(.A(new_n654), .B(new_n749), .C1(new_n682), .C2(new_n687), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n753), .B1(new_n754), .B2(new_n586), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n424), .A2(new_n586), .A3(new_n718), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n756), .B1(new_n743), .B2(new_n744), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT108), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n755), .B2(new_n757), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n762));
  AND3_X1   g561(.A1(new_n740), .A2(new_n762), .A3(new_n741), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n762), .B1(new_n740), .B2(new_n741), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n756), .B1(new_n765), .B2(new_n743), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n754), .A2(new_n586), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT52), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n759), .A2(new_n761), .A3(new_n768), .ZN(G1337gat));
  AND2_X1   g568(.A1(new_n750), .A2(new_n701), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n770), .A2(KEYINPUT109), .ZN(new_n771));
  OAI21_X1  g570(.A(G99gat), .B1(new_n770), .B2(KEYINPUT109), .ZN(new_n772));
  INV_X1    g571(.A(G99gat), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n666), .A2(new_n773), .A3(new_n718), .ZN(new_n774));
  OAI22_X1  g573(.A1(new_n771), .A2(new_n772), .B1(new_n745), .B2(new_n774), .ZN(G1338gat));
  NAND2_X1  g574(.A1(new_n682), .A2(new_n687), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n776), .A2(new_n431), .A3(new_n748), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT53), .B1(new_n777), .B2(G106gat), .ZN(new_n778));
  INV_X1    g577(.A(G106gat), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n431), .A2(new_n779), .A3(new_n718), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n778), .B1(new_n745), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n780), .B1(new_n765), .B2(new_n743), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT110), .ZN(new_n783));
  AOI211_X1 g582(.A(new_n783), .B(new_n779), .C1(new_n750), .C2(new_n431), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT110), .B1(new_n777), .B2(G106gat), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n782), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n781), .B1(new_n786), .B2(new_n787), .ZN(G1339gat));
  XNOR2_X1  g587(.A(new_n472), .B(KEYINPUT102), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n790));
  INV_X1    g589(.A(new_n533), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n523), .A2(new_n531), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n525), .B1(new_n516), .B2(new_n523), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n792), .B1(new_n793), .B2(KEYINPUT112), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT112), .ZN(new_n795));
  AOI211_X1 g594(.A(new_n795), .B(new_n525), .C1(new_n516), .C2(new_n523), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n540), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n718), .A2(new_n790), .A3(new_n544), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n544), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT113), .B1(new_n799), .B2(new_n647), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n628), .A2(new_n803), .ZN(new_n804));
  OR2_X1    g603(.A1(new_n643), .A2(new_n615), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT101), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n627), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n643), .A2(KEYINPUT101), .A3(new_n615), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n808), .A2(new_n803), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT111), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n810), .A2(new_n811), .A3(new_n639), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n811), .B1(new_n810), .B2(new_n639), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n806), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n804), .A2(new_n805), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n644), .A2(new_n645), .A3(KEYINPUT54), .ZN(new_n817));
  OAI21_X1  g616(.A(KEYINPUT111), .B1(new_n817), .B2(new_n638), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n810), .A2(new_n811), .A3(new_n639), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n816), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n717), .B(new_n814), .C1(new_n820), .C2(KEYINPUT55), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n801), .B1(new_n821), .B2(new_n679), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n613), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n821), .A2(new_n613), .ZN(new_n824));
  INV_X1    g623(.A(new_n799), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n823), .A2(KEYINPUT114), .A3(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n818), .A2(new_n819), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n640), .B1(new_n829), .B2(new_n806), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n815), .B1(new_n812), .B2(new_n813), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n802), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n830), .A2(new_n832), .A3(new_n545), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n611), .B1(new_n833), .B2(new_n801), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n821), .A2(new_n613), .A3(new_n799), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n828), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n827), .A2(new_n579), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n649), .A2(new_n679), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n789), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n345), .A2(new_n421), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n840), .A2(new_n424), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(new_n253), .A3(new_n545), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n431), .B1(new_n837), .B2(new_n838), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n650), .A2(new_n428), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(G113gat), .B1(new_n846), .B2(new_n547), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  XOR2_X1   g647(.A(new_n848), .B(KEYINPUT115), .Z(G1340gat));
  INV_X1    g648(.A(G120gat), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n846), .A2(new_n850), .A3(new_n647), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n842), .A2(new_n718), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n852), .B2(new_n850), .ZN(G1341gat));
  INV_X1    g652(.A(G127gat), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n842), .A2(new_n854), .A3(new_n578), .ZN(new_n855));
  OAI21_X1  g654(.A(G127gat), .B1(new_n846), .B2(new_n579), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1342gat));
  NAND2_X1  g656(.A1(new_n654), .A2(new_n611), .ZN(new_n858));
  NOR4_X1   g657(.A1(new_n840), .A2(G134gat), .A3(new_n841), .A4(new_n858), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT56), .ZN(new_n860));
  OAI21_X1  g659(.A(G134gat), .B1(new_n846), .B2(new_n613), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(KEYINPUT116), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n861), .A2(KEYINPUT116), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n860), .B1(new_n862), .B2(new_n863), .ZN(G1343gat));
  INV_X1    g663(.A(KEYINPUT58), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n837), .A2(new_n838), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n867), .A3(new_n431), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n424), .B1(new_n435), .B2(new_n436), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n650), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT117), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n870), .B(new_n871), .ZN(new_n872));
  XNOR2_X1  g671(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n820), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n814), .A2(new_n717), .ZN(new_n876));
  OAI21_X1  g675(.A(KEYINPUT119), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n831), .A2(new_n873), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n830), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n877), .A2(new_n546), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n825), .A2(new_n718), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n611), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n579), .B1(new_n883), .B2(new_n835), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n342), .B1(new_n884), .B2(new_n838), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n868), .B(new_n872), .C1(new_n867), .C2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(G141gat), .B1(new_n886), .B2(new_n679), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n664), .A2(new_n431), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT120), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n547), .A2(G141gat), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n839), .A2(new_n889), .A3(new_n654), .A4(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n865), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n865), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n885), .A2(new_n867), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n894), .A2(new_n546), .A3(new_n868), .A4(new_n872), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n893), .B1(new_n895), .B2(G141gat), .ZN(new_n896));
  OAI21_X1  g695(.A(KEYINPUT121), .B1(new_n892), .B2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT121), .ZN(new_n898));
  OAI21_X1  g697(.A(G141gat), .B1(new_n886), .B2(new_n547), .ZN(new_n899));
  INV_X1    g698(.A(new_n893), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(new_n891), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n894), .A2(new_n545), .A3(new_n868), .A4(new_n872), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n903), .B2(G141gat), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n898), .B(new_n901), .C1(new_n904), .C2(new_n865), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n897), .A2(new_n905), .ZN(G1344gat));
  NAND2_X1  g705(.A1(new_n839), .A2(new_n889), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(new_n424), .ZN(new_n908));
  INV_X1    g707(.A(G148gat), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n909), .A3(new_n718), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n886), .A2(new_n647), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n911), .A2(KEYINPUT59), .A3(new_n909), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT59), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n866), .A2(new_n431), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT57), .ZN(new_n915));
  INV_X1    g714(.A(new_n883), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n799), .B1(new_n824), .B2(KEYINPUT122), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n917), .B1(KEYINPUT122), .B2(new_n824), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n578), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n648), .A2(new_n546), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n867), .B(new_n431), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n915), .A2(new_n921), .A3(new_n718), .A4(new_n872), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n913), .B1(new_n922), .B2(G148gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n910), .B1(new_n912), .B2(new_n923), .ZN(G1345gat));
  OAI21_X1  g723(.A(G155gat), .B1(new_n886), .B2(new_n579), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n908), .A2(new_n300), .A3(new_n578), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1346gat));
  OAI21_X1  g726(.A(G162gat), .B1(new_n886), .B2(new_n613), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n654), .A2(new_n301), .A3(new_n611), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n928), .B1(new_n907), .B2(new_n929), .ZN(G1347gat));
  NAND3_X1  g729(.A1(new_n789), .A2(new_n666), .A3(new_n424), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n866), .A2(new_n342), .A3(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT125), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n844), .A2(KEYINPUT125), .A3(new_n932), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(G169gat), .B1(new_n937), .B2(new_n547), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n650), .B1(new_n837), .B2(new_n838), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(KEYINPUT123), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n424), .B1(new_n939), .B2(KEYINPUT123), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n941), .A2(new_n942), .A3(new_n841), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n679), .A2(G169gat), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n944), .B1(new_n943), .B2(new_n945), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n938), .B1(new_n946), .B2(new_n947), .ZN(G1348gat));
  INV_X1    g747(.A(G176gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n943), .A2(new_n949), .A3(new_n718), .ZN(new_n950));
  OAI21_X1  g749(.A(G176gat), .B1(new_n937), .B2(new_n647), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(G1349gat));
  NAND3_X1  g751(.A1(new_n935), .A2(new_n578), .A3(new_n936), .ZN(new_n953));
  AOI22_X1  g752(.A1(new_n953), .A2(G183gat), .B1(KEYINPUT126), .B2(KEYINPUT60), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n578), .A2(new_n225), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n943), .A2(new_n955), .ZN(new_n956));
  OR2_X1    g755(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n954), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n954), .B2(new_n956), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n958), .A2(new_n959), .ZN(G1350gat));
  NAND3_X1  g759(.A1(new_n943), .A2(new_n217), .A3(new_n611), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n935), .A2(new_n611), .A3(new_n936), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n962), .A2(new_n963), .A3(G190gat), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n963), .B1(new_n962), .B2(G190gat), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n961), .B1(new_n964), .B2(new_n965), .ZN(G1351gat));
  NOR3_X1   g765(.A1(new_n650), .A2(new_n701), .A3(new_n654), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n915), .A2(new_n921), .A3(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(G197gat), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n968), .A2(new_n969), .A3(new_n547), .ZN(new_n970));
  NOR3_X1   g769(.A1(new_n941), .A2(new_n942), .A3(new_n888), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(new_n545), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n970), .B1(new_n969), .B2(new_n972), .ZN(G1352gat));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT127), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n647), .A2(G204gat), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n975), .B1(new_n971), .B2(new_n976), .ZN(new_n977));
  INV_X1    g776(.A(new_n939), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT123), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g779(.A(new_n888), .ZN(new_n981));
  NAND4_X1  g780(.A1(new_n980), .A2(new_n424), .A3(new_n981), .A4(new_n940), .ZN(new_n982));
  INV_X1    g781(.A(new_n976), .ZN(new_n983));
  NOR3_X1   g782(.A1(new_n982), .A2(KEYINPUT127), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n974), .B1(new_n977), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g784(.A(G204gat), .B1(new_n968), .B2(new_n647), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n971), .A2(new_n975), .A3(new_n976), .ZN(new_n987));
  OAI21_X1  g786(.A(KEYINPUT127), .B1(new_n982), .B2(new_n983), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n987), .A2(new_n988), .A3(KEYINPUT62), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n985), .A2(new_n986), .A3(new_n989), .ZN(G1353gat));
  OR3_X1    g789(.A1(new_n982), .A2(G211gat), .A3(new_n579), .ZN(new_n991));
  OR2_X1    g790(.A1(new_n968), .A2(new_n579), .ZN(new_n992));
  AOI21_X1  g791(.A(KEYINPUT63), .B1(new_n992), .B2(G211gat), .ZN(new_n993));
  OAI211_X1 g792(.A(KEYINPUT63), .B(G211gat), .C1(new_n968), .C2(new_n579), .ZN(new_n994));
  INV_X1    g793(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n991), .B1(new_n993), .B2(new_n995), .ZN(G1354gat));
  OAI21_X1  g795(.A(G218gat), .B1(new_n968), .B2(new_n613), .ZN(new_n997));
  OR2_X1    g796(.A1(new_n613), .A2(G218gat), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n997), .B1(new_n982), .B2(new_n998), .ZN(G1355gat));
endmodule


