//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 1 0 1 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 0 0 0 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 1 1 0 1 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1181, new_n1182, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT66), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G50), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  OAI22_X1  g0015(.A1(new_n213), .A2(KEYINPUT67), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n216), .B1(KEYINPUT67), .B2(new_n213), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G116), .ZN(new_n220));
  INV_X1    g0020(.A(G270), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AND2_X1   g0022(.A1(G77), .A2(G244), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n209), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OR2_X1    g0024(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT68), .Z(new_n226));
  NAND2_X1  g0026(.A1(new_n203), .A2(G50), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT65), .Z(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR3_X1   g0030(.A1(new_n229), .A2(new_n207), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n209), .A2(G13), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n232), .B(G250), .C1(G257), .C2(G264), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT0), .Z(new_n234));
  AND2_X1   g0034(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n235));
  NOR4_X1   g0035(.A1(new_n226), .A2(new_n231), .A3(new_n234), .A4(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n221), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n214), .ZN(new_n246));
  INV_X1    g0046(.A(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  INV_X1    g0049(.A(G107), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(new_n220), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n248), .B(new_n252), .ZN(G351));
  NAND3_X1  g0053(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(G50), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n230), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n206), .A2(G20), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n256), .B1(new_n261), .B2(G50), .ZN(new_n262));
  XOR2_X1   g0062(.A(new_n262), .B(KEYINPUT70), .Z(new_n263));
  XOR2_X1   g0063(.A(KEYINPUT8), .B(G58), .Z(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(G20), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G150), .ZN(new_n269));
  NOR2_X1   g0069(.A1(G20), .A2(G33), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  OAI22_X1  g0071(.A1(new_n265), .A2(new_n268), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n201), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n207), .B1(new_n273), .B2(new_n202), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n258), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  AND2_X1   g0075(.A1(new_n263), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n276), .B1(KEYINPUT72), .B2(KEYINPUT9), .ZN(new_n277));
  NAND2_X1  g0077(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n277), .B(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT69), .B(G1698), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n280), .A2(G222), .B1(G223), .B2(G1698), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT3), .B(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n283), .B(new_n284), .C1(G77), .C2(new_n282), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n286));
  INV_X1    g0086(.A(G274), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n284), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n286), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n285), .B(new_n289), .C1(new_n215), .C2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G190), .ZN(new_n293));
  OR2_X1    g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT73), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n292), .A2(G200), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n294), .A2(new_n295), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  OR3_X1    g0099(.A1(new_n279), .A2(KEYINPUT10), .A3(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(KEYINPUT10), .B1(new_n279), .B2(new_n299), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G33), .A2(G97), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n280), .A2(G226), .B1(G232), .B2(G1698), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n266), .A2(KEYINPUT3), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT3), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G33), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n304), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n288), .B1(new_n310), .B2(new_n284), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(new_n219), .B2(new_n291), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n312), .B(KEYINPUT13), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n313), .A2(KEYINPUT75), .A3(G169), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT14), .ZN(new_n315));
  INV_X1    g0115(.A(new_n313), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G179), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT14), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n313), .A2(KEYINPUT75), .A3(new_n318), .A4(G169), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n315), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n254), .A2(G68), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT12), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  XOR2_X1   g0123(.A(new_n323), .B(KEYINPUT74), .Z(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(new_n322), .B2(new_n321), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n267), .A2(G77), .B1(G20), .B2(new_n218), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n270), .A2(G50), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n259), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  XOR2_X1   g0128(.A(new_n328), .B(KEYINPUT11), .Z(new_n329));
  INV_X1    g0129(.A(new_n261), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G68), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n325), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  XOR2_X1   g0132(.A(new_n332), .B(KEYINPUT76), .Z(new_n333));
  NAND2_X1  g0133(.A1(new_n320), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G200), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n316), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n332), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(new_n313), .B2(new_n293), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n280), .A2(G232), .B1(G238), .B2(G1698), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n282), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT71), .B(G107), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n342), .B(new_n284), .C1(new_n282), .C2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n291), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G244), .ZN(new_n347));
  AND3_X1   g0147(.A1(new_n345), .A2(new_n289), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G190), .ZN(new_n349));
  INV_X1    g0149(.A(G77), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n255), .A2(new_n350), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n264), .A2(new_n270), .B1(G20), .B2(G77), .ZN(new_n352));
  XOR2_X1   g0152(.A(KEYINPUT15), .B(G87), .Z(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n352), .B1(new_n268), .B2(new_n354), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n355), .A2(new_n258), .B1(G77), .B2(new_n330), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n345), .A2(new_n289), .A3(new_n347), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G200), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n349), .A2(new_n351), .A3(new_n356), .A4(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G179), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n348), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G169), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n356), .A2(new_n351), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n361), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n359), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n276), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n292), .A2(new_n362), .ZN(new_n368));
  OR2_X1    g0168(.A1(new_n292), .A2(G179), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n334), .A2(new_n340), .A3(new_n366), .A4(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT16), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT7), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(new_n282), .B2(G20), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n309), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n218), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AND2_X1   g0176(.A1(G58), .A2(G68), .ZN(new_n377));
  OAI21_X1  g0177(.A(G20), .B1(new_n377), .B2(new_n202), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT78), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n270), .A2(G159), .ZN(new_n381));
  OAI211_X1 g0181(.A(KEYINPUT78), .B(G20), .C1(new_n377), .C2(new_n202), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n372), .B1(new_n376), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT79), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI211_X1 g0186(.A(KEYINPUT79), .B(new_n372), .C1(new_n376), .C2(new_n383), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT77), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n266), .B2(KEYINPUT3), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n307), .A2(KEYINPUT77), .A3(G33), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(G20), .B1(new_n392), .B2(new_n306), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n218), .B1(new_n393), .B2(new_n373), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n390), .A2(new_n391), .B1(KEYINPUT3), .B2(new_n266), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT7), .B1(new_n395), .B2(G20), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n383), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n259), .B1(new_n397), .B2(KEYINPUT16), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n388), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT80), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n264), .A2(new_n260), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n402), .B(KEYINPUT81), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n403), .A2(new_n259), .A3(new_n254), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n265), .A2(new_n255), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT82), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT82), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n404), .A2(new_n408), .A3(new_n405), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n388), .A2(new_n398), .A3(KEYINPUT80), .ZN(new_n411));
  AND3_X1   g0211(.A1(new_n401), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n280), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n392), .A2(new_n306), .ZN(new_n414));
  INV_X1    g0214(.A(G87), .ZN(new_n415));
  OAI22_X1  g0215(.A1(new_n413), .A2(new_n414), .B1(new_n266), .B2(new_n415), .ZN(new_n416));
  OR2_X1    g0216(.A1(new_n416), .A2(KEYINPUT83), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(KEYINPUT83), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(new_n284), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n288), .B1(new_n346), .B2(G232), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(G200), .ZN(new_n422));
  XOR2_X1   g0222(.A(KEYINPUT84), .B(G190), .Z(new_n423));
  NAND3_X1  g0223(.A1(new_n419), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n412), .A2(KEYINPUT17), .A3(new_n422), .A4(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT17), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n401), .A2(new_n410), .A3(new_n424), .A4(new_n411), .ZN(new_n427));
  INV_X1    g0227(.A(new_n422), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n401), .A2(new_n410), .A3(new_n411), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n421), .A2(G169), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(new_n360), .B2(new_n421), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n430), .A2(new_n432), .A3(KEYINPUT18), .ZN(new_n433));
  AOI21_X1  g0233(.A(KEYINPUT18), .B1(new_n430), .B2(new_n432), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n425), .B(new_n429), .C1(new_n433), .C2(new_n434), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n303), .A2(new_n371), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n343), .A2(G20), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G33), .A2(G116), .ZN(new_n439));
  OR3_X1    g0239(.A1(new_n439), .A2(KEYINPUT94), .A3(G20), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT94), .B1(new_n439), .B2(G20), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n438), .A2(KEYINPUT23), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n395), .A2(KEYINPUT22), .A3(new_n207), .A4(G87), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT22), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n207), .A2(G87), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n309), .B2(new_n445), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n447));
  XNOR2_X1  g0247(.A(new_n447), .B(KEYINPUT95), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n442), .A2(new_n443), .A3(new_n446), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT96), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n450), .A2(KEYINPUT24), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n450), .A2(KEYINPUT24), .ZN(new_n452));
  OAI22_X1  g0252(.A1(new_n451), .A2(new_n452), .B1(KEYINPUT96), .B2(new_n449), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n258), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n255), .A2(new_n250), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT97), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT25), .ZN(new_n457));
  XOR2_X1   g0257(.A(KEYINPUT97), .B(KEYINPUT25), .Z(new_n458));
  OAI211_X1 g0258(.A(new_n259), .B(new_n254), .C1(G1), .C2(new_n266), .ZN(new_n459));
  OAI221_X1 g0259(.A(new_n457), .B1(new_n455), .B2(new_n458), .C1(new_n459), .C2(new_n250), .ZN(new_n460));
  XOR2_X1   g0260(.A(new_n460), .B(KEYINPUT98), .Z(new_n461));
  AND2_X1   g0261(.A1(new_n206), .A2(G45), .ZN(new_n462));
  AND2_X1   g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  NOR2_X1   g0263(.A1(KEYINPUT5), .A2(G41), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OR2_X1    g0265(.A1(new_n465), .A2(new_n287), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n280), .A2(G250), .B1(G257), .B2(G1698), .ZN(new_n468));
  INV_X1    g0268(.A(G294), .ZN(new_n469));
  OAI22_X1  g0269(.A1(new_n468), .A2(new_n414), .B1(new_n266), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n284), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n467), .B1(new_n471), .B2(KEYINPUT99), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n465), .A2(new_n290), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G264), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n472), .B(new_n474), .C1(KEYINPUT99), .C2(new_n471), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n471), .A2(new_n466), .A3(new_n474), .ZN(new_n476));
  OAI22_X1  g0276(.A1(new_n475), .A2(G190), .B1(G200), .B2(new_n476), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n454), .A2(new_n461), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n475), .A2(G169), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n476), .A2(G179), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n454), .A2(new_n461), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G250), .A2(G1698), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n280), .A2(G244), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT4), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n486), .A2(new_n282), .B1(G33), .B2(G283), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n485), .B1(new_n414), .B2(new_n484), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n290), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n473), .A2(G257), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NOR3_X1   g0291(.A1(new_n489), .A2(new_n467), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(KEYINPUT86), .B1(new_n492), .B2(new_n335), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n254), .A2(G97), .ZN(new_n494));
  INV_X1    g0294(.A(new_n459), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n494), .B1(new_n495), .B2(G97), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT6), .ZN(new_n497));
  INV_X1    g0297(.A(G97), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(new_n250), .ZN(new_n499));
  NOR2_X1   g0299(.A1(G97), .A2(G107), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n497), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n250), .A2(KEYINPUT6), .A3(G97), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(new_n207), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n343), .B1(new_n374), .B2(new_n375), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n270), .A2(G77), .ZN(new_n506));
  XNOR2_X1  g0306(.A(new_n506), .B(KEYINPUT85), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n504), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n496), .B1(new_n508), .B2(new_n259), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n509), .B1(new_n492), .B2(G190), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n487), .A2(new_n488), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n466), .B(new_n490), .C1(new_n511), .C2(new_n290), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT86), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n512), .A2(new_n513), .A3(G200), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n493), .A2(new_n510), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n512), .A2(new_n362), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n492), .A2(new_n360), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n516), .A2(new_n517), .A3(new_n509), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n395), .A2(G264), .A3(G1698), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT93), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n309), .A2(G303), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT93), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n395), .A2(new_n523), .A3(G264), .A4(G1698), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n395), .A2(G257), .A3(new_n280), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n521), .A2(new_n522), .A3(new_n524), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n284), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n473), .A2(G270), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n527), .A2(new_n466), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n495), .A2(G116), .ZN(new_n530));
  AOI21_X1  g0330(.A(G20), .B1(new_n266), .B2(G97), .ZN(new_n531));
  INV_X1    g0331(.A(G283), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n531), .B1(new_n266), .B2(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n533), .B(new_n258), .C1(new_n207), .C2(G116), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT20), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n534), .A2(new_n535), .ZN(new_n537));
  OAI221_X1 g0337(.A(new_n530), .B1(G116), .B2(new_n254), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n529), .A2(G169), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT21), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n529), .A2(G200), .ZN(new_n542));
  INV_X1    g0342(.A(new_n538), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n527), .A2(new_n423), .A3(new_n466), .A4(new_n528), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n529), .A2(new_n360), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n538), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n529), .A2(KEYINPUT21), .A3(G169), .A4(new_n538), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n541), .A2(new_n545), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n519), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n495), .A2(G87), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n280), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n439), .B1(new_n552), .B2(new_n414), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n284), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n462), .A2(G250), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n555), .A2(new_n284), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n462), .A2(new_n287), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n293), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(G200), .B2(new_n559), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT19), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT87), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT87), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(KEYINPUT19), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n207), .B1(new_n566), .B2(new_n304), .ZN(new_n567));
  NOR2_X1   g0367(.A1(G87), .A2(G97), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT88), .B1(new_n343), .B2(new_n568), .ZN(new_n569));
  AND2_X1   g0369(.A1(KEYINPUT71), .A2(G107), .ZN(new_n570));
  NOR2_X1   g0370(.A1(KEYINPUT71), .A2(G107), .ZN(new_n571));
  OAI211_X1 g0371(.A(KEYINPUT88), .B(new_n568), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n567), .B1(new_n569), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n566), .B1(new_n268), .B2(new_n498), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n395), .A2(new_n207), .A3(G68), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT89), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT89), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n574), .A2(new_n579), .A3(new_n575), .A4(new_n576), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n258), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n354), .A2(new_n255), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n581), .A2(KEYINPUT90), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(KEYINPUT90), .B1(new_n581), .B2(new_n582), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n551), .B(new_n561), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT92), .ZN(new_n586));
  XNOR2_X1  g0386(.A(new_n353), .B(KEYINPUT91), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n587), .A2(new_n459), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n581), .A2(new_n582), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT90), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n581), .A2(KEYINPUT90), .A3(new_n582), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n588), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n559), .A2(new_n360), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(G169), .B2(new_n559), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n585), .B(new_n586), .C1(new_n593), .C2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n588), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n583), .B2(new_n584), .ZN(new_n599));
  INV_X1    g0399(.A(new_n595), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n586), .B1(new_n601), .B2(new_n585), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n482), .B(new_n550), .C1(new_n597), .C2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n437), .A2(new_n603), .ZN(G372));
  INV_X1    g0404(.A(new_n370), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n303), .A2(KEYINPUT102), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n300), .A2(KEYINPUT102), .A3(new_n301), .ZN(new_n607));
  OR2_X1    g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OR2_X1    g0408(.A1(new_n433), .A2(new_n434), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n425), .A2(new_n429), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n365), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n340), .A2(new_n612), .B1(new_n320), .B2(new_n333), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n609), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n605), .B1(new_n608), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n518), .ZN(new_n616));
  XOR2_X1   g0416(.A(KEYINPUT101), .B(KEYINPUT26), .Z(new_n617));
  OAI211_X1 g0417(.A(new_n616), .B(new_n617), .C1(new_n597), .C2(new_n602), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT26), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n585), .B1(new_n593), .B2(new_n595), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n619), .B1(new_n620), .B2(new_n518), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n541), .A2(new_n547), .A3(new_n548), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n481), .A2(new_n623), .ZN(new_n624));
  OR2_X1    g0424(.A1(new_n624), .A2(KEYINPUT100), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n620), .A2(new_n478), .A3(new_n519), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n624), .A2(KEYINPUT100), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n622), .A2(new_n628), .A3(new_n601), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n615), .B1(new_n437), .B2(new_n630), .ZN(G369));
  INV_X1    g0431(.A(new_n482), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n633));
  XNOR2_X1  g0433(.A(new_n633), .B(KEYINPUT103), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT27), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(new_n637), .A3(G213), .ZN(new_n638));
  INV_X1    g0438(.A(G343), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n641), .B1(new_n454), .B2(new_n461), .ZN(new_n642));
  INV_X1    g0442(.A(new_n481), .ZN(new_n643));
  OAI22_X1  g0443(.A1(new_n632), .A2(new_n642), .B1(new_n643), .B2(new_n641), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n543), .A2(new_n641), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n623), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n549), .B2(new_n645), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n647), .A2(G330), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n481), .A2(new_n641), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n623), .A2(new_n641), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n482), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n649), .A2(new_n650), .A3(new_n653), .ZN(G399));
  OR3_X1    g0454(.A1(new_n569), .A2(new_n573), .A3(G116), .ZN(new_n655));
  INV_X1    g0455(.A(new_n232), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n656), .A2(G41), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n655), .A2(new_n657), .A3(new_n206), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n658), .B1(new_n228), .B2(new_n657), .ZN(new_n659));
  XOR2_X1   g0459(.A(new_n659), .B(KEYINPUT28), .Z(new_n660));
  NOR3_X1   g0460(.A1(new_n620), .A2(new_n619), .A3(new_n518), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n620), .A2(KEYINPUT92), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n518), .B1(new_n663), .B2(new_n596), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n662), .B1(new_n664), .B2(new_n617), .ZN(new_n665));
  INV_X1    g0465(.A(new_n601), .ZN(new_n666));
  INV_X1    g0466(.A(new_n624), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n666), .B1(new_n626), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n640), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT29), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n666), .B1(new_n618), .B2(new_n621), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n640), .B1(new_n671), .B2(new_n628), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n670), .B1(new_n672), .B2(KEYINPUT29), .ZN(new_n673));
  INV_X1    g0473(.A(new_n559), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n512), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n675), .A2(new_n471), .A3(new_n546), .A4(new_n474), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT30), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n529), .A2(new_n674), .ZN(new_n680));
  OR4_X1    g0480(.A1(G179), .A2(new_n680), .A3(new_n476), .A4(new_n492), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n678), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n640), .ZN(new_n683));
  OAI211_X1 g0483(.A(KEYINPUT31), .B(new_n683), .C1(new_n603), .C2(new_n640), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n683), .A2(KEYINPUT31), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G330), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n673), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n660), .B1(new_n688), .B2(G1), .ZN(G364));
  NAND2_X1  g0489(.A1(new_n207), .A2(G13), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT104), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G45), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G1), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(new_n657), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n648), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(G330), .B2(new_n647), .ZN(new_n696));
  NOR2_X1   g0496(.A1(G13), .A2(G33), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(G20), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n647), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n230), .B1(G20), .B2(new_n362), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(KEYINPUT105), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(KEYINPUT105), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n207), .A2(G190), .ZN(new_n706));
  NOR2_X1   g0506(.A1(G179), .A2(G200), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n709), .A2(G329), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n207), .A2(new_n360), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n423), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G200), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n335), .ZN(new_n714));
  AOI22_X1  g0514(.A1(G322), .A2(new_n713), .B1(new_n714), .B2(G326), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n207), .B1(new_n707), .B2(G190), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n715), .B(new_n309), .C1(new_n469), .C2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n706), .A2(G179), .A3(G200), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  XNOR2_X1  g0519(.A(KEYINPUT33), .B(G317), .ZN(new_n720));
  AOI211_X1 g0520(.A(new_n710), .B(new_n717), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n711), .A2(new_n293), .A3(new_n335), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G311), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n335), .A2(G179), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n706), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n721), .B(new_n724), .C1(new_n532), .C2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n725), .A2(G20), .A3(G190), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n727), .B1(G303), .B2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n716), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n719), .A2(G68), .B1(new_n731), .B2(G97), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT32), .ZN(new_n733));
  XNOR2_X1  g0533(.A(KEYINPUT106), .B(G159), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n708), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n732), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n729), .A2(G87), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n282), .ZN(new_n739));
  XOR2_X1   g0539(.A(new_n739), .B(KEYINPUT107), .Z(new_n740));
  AOI211_X1 g0540(.A(new_n737), .B(new_n740), .C1(G58), .C2(new_n713), .ZN(new_n741));
  INV_X1    g0541(.A(new_n726), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G107), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n736), .A2(new_n733), .B1(G77), .B2(new_n723), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n741), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n745), .B1(G50), .B2(new_n714), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n705), .B1(new_n730), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n656), .A2(new_n309), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G355), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n248), .A2(G45), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n656), .A2(new_n395), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(new_n229), .B2(G45), .ZN(new_n752));
  OAI221_X1 g0552(.A(new_n749), .B1(G116), .B2(new_n232), .C1(new_n750), .C2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n705), .A2(new_n699), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n701), .A2(new_n747), .A3(new_n755), .A4(new_n694), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n696), .A2(new_n756), .ZN(G396));
  NAND4_X1  g0557(.A1(new_n361), .A2(new_n364), .A3(new_n363), .A4(new_n640), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT109), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n640), .A2(new_n364), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n366), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(KEYINPUT108), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT108), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n366), .A2(new_n763), .A3(new_n760), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n759), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n672), .B(new_n766), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n767), .A2(new_n687), .ZN(new_n768));
  INV_X1    g0568(.A(new_n694), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n767), .A2(new_n687), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n766), .A2(new_n698), .ZN(new_n772));
  INV_X1    g0572(.A(new_n705), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n713), .A2(G143), .B1(G150), .B2(new_n719), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(new_n735), .B2(new_n722), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(G137), .B2(new_n714), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT34), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n726), .A2(new_n218), .ZN(new_n778));
  INV_X1    g0578(.A(G132), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n395), .B1(new_n779), .B2(new_n708), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n777), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n781), .B1(new_n214), .B2(new_n728), .C1(new_n247), .C2(new_n716), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n722), .A2(new_n220), .B1(new_n728), .B2(new_n250), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n282), .B(new_n783), .C1(G283), .C2(new_n719), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n709), .A2(G311), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n714), .A2(G303), .B1(G97), .B2(new_n731), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n726), .A2(new_n415), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(new_n713), .B2(G294), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n784), .A2(new_n785), .A3(new_n786), .A4(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n773), .B1(new_n782), .B2(new_n789), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n772), .A2(new_n790), .A3(new_n769), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n705), .A2(new_n697), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n791), .B1(G77), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n771), .A2(new_n794), .ZN(G384));
  INV_X1    g0595(.A(KEYINPUT40), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n333), .A2(new_n640), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n334), .A2(new_n340), .A3(new_n797), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n333), .B(new_n640), .C1(new_n320), .C2(new_n339), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n765), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AND3_X1   g0600(.A1(new_n684), .A2(new_n685), .A3(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n638), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n435), .A2(new_n430), .A3(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n412), .A2(new_n422), .A3(new_n424), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n430), .B1(new_n432), .B2(new_n802), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(KEYINPUT37), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT37), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n804), .A2(new_n808), .A3(new_n805), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n803), .A2(new_n810), .ZN(new_n811));
  XOR2_X1   g0611(.A(KEYINPUT111), .B(KEYINPUT38), .Z(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n397), .A2(KEYINPUT16), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n406), .B1(new_n814), .B2(new_n398), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n435), .A2(new_n802), .A3(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n432), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n815), .B1(new_n818), .B2(new_n638), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n427), .A2(new_n428), .ZN(new_n820));
  OAI21_X1  g0620(.A(KEYINPUT37), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n809), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n817), .A2(KEYINPUT38), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n813), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n796), .B1(new_n801), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n823), .ZN(new_n826));
  AOI21_X1  g0626(.A(KEYINPUT38), .B1(new_n817), .B2(new_n822), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n684), .A2(new_n796), .A3(new_n685), .A4(new_n800), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n436), .B(new_n686), .C1(new_n825), .C2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G330), .ZN(new_n832));
  INV_X1    g0632(.A(new_n812), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(new_n803), .B2(new_n810), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n826), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n684), .A2(new_n800), .A3(new_n685), .ZN(new_n836));
  OAI21_X1  g0636(.A(KEYINPUT40), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n817), .A2(new_n822), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT38), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n823), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n801), .A2(new_n796), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n832), .B1(new_n837), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n686), .A2(new_n436), .A3(G330), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n831), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT112), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n670), .B(new_n436), .C1(KEYINPUT29), .C2(new_n672), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n615), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n847), .B(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n798), .A2(new_n799), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n640), .B(new_n765), .C1(new_n671), .C2(new_n628), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n365), .A2(new_n640), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n841), .B(new_n851), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  OR2_X1    g0654(.A1(new_n609), .A2(new_n802), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT39), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n826), .B2(new_n834), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n840), .A2(KEYINPUT39), .A3(new_n823), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n334), .A2(new_n640), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT110), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n859), .B(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n857), .A2(new_n858), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n854), .A2(new_n855), .A3(new_n862), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n850), .B(new_n863), .Z(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n206), .B2(new_n691), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT35), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n207), .B(new_n230), .C1(new_n503), .C2(new_n866), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n867), .B(G116), .C1(new_n866), .C2(new_n503), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT36), .ZN(new_n869));
  INV_X1    g0669(.A(G13), .ZN(new_n870));
  NOR3_X1   g0670(.A1(new_n229), .A2(new_n350), .A3(new_n377), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n201), .A2(new_n218), .ZN(new_n872));
  OAI211_X1 g0672(.A(G1), .B(new_n870), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n865), .A2(new_n869), .A3(new_n873), .ZN(G367));
  NAND2_X1  g0674(.A1(new_n616), .A2(new_n640), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n509), .A2(new_n640), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n515), .A2(new_n518), .A3(new_n876), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n653), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n879), .B(KEYINPUT42), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n518), .B1(new_n643), .B2(new_n877), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n641), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n591), .A2(new_n592), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n641), .B1(new_n883), .B2(new_n551), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n666), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n620), .B2(new_n884), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n880), .A2(new_n882), .B1(KEYINPUT43), .B2(new_n886), .ZN(new_n887));
  OR2_X1    g0687(.A1(new_n886), .A2(KEYINPUT43), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n887), .B(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n649), .A2(new_n878), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n889), .B(new_n890), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n657), .B(KEYINPUT41), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n653), .A2(new_n650), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n878), .ZN(new_n895));
  XOR2_X1   g0695(.A(new_n895), .B(KEYINPUT44), .Z(new_n896));
  NOR2_X1   g0696(.A1(new_n894), .A2(new_n878), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(KEYINPUT45), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n896), .A2(new_n649), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n649), .B1(new_n896), .B2(new_n898), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n653), .B1(new_n644), .B2(new_n652), .ZN(new_n902));
  INV_X1    g0702(.A(new_n648), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n904), .A2(new_n649), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n673), .A2(new_n687), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT113), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT113), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n673), .A2(new_n908), .A3(new_n687), .A4(new_n905), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n901), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n893), .B1(new_n910), .B2(new_n688), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n891), .B1(new_n911), .B2(new_n693), .ZN(new_n912));
  INV_X1    g0712(.A(new_n713), .ZN(new_n913));
  INV_X1    g0713(.A(G303), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n913), .A2(new_n914), .B1(new_n532), .B2(new_n722), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT46), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n728), .B2(new_n220), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n915), .B1(KEYINPUT114), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(KEYINPUT114), .B2(new_n917), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n716), .A2(new_n343), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n728), .A2(new_n916), .A3(new_n220), .ZN(new_n921));
  NOR4_X1   g0721(.A1(new_n919), .A2(new_n395), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n714), .A2(G311), .B1(G317), .B2(new_n709), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI221_X1 g0724(.A(new_n924), .B1(new_n498), .B2(new_n726), .C1(new_n469), .C2(new_n718), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n719), .A2(new_n734), .ZN(new_n926));
  INV_X1    g0726(.A(new_n714), .ZN(new_n927));
  INV_X1    g0727(.A(G143), .ZN(new_n928));
  OAI221_X1 g0728(.A(new_n926), .B1(new_n247), .B2(new_n728), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(G137), .B2(new_n709), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n731), .A2(G68), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n723), .A2(new_n201), .B1(new_n742), .B2(G77), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n282), .B1(new_n913), .B2(new_n269), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n925), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT47), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n705), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n886), .A2(new_n700), .ZN(new_n938));
  INV_X1    g0738(.A(new_n751), .ZN(new_n939));
  OAI221_X1 g0739(.A(new_n754), .B1(new_n232), .B2(new_n354), .C1(new_n243), .C2(new_n939), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n937), .A2(new_n694), .A3(new_n938), .A4(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n912), .A2(new_n941), .ZN(G387));
  NOR2_X1   g0742(.A1(new_n644), .A2(new_n700), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n728), .A2(new_n350), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n587), .A2(new_n716), .ZN(new_n945));
  AOI211_X1 g0745(.A(new_n944), .B(new_n945), .C1(G159), .C2(new_n714), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n414), .B1(G150), .B2(new_n709), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n713), .A2(G50), .B1(G97), .B2(new_n742), .ZN(new_n948));
  AOI22_X1  g0748(.A1(G68), .A2(new_n723), .B1(new_n719), .B2(new_n264), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT115), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n946), .A2(new_n947), .A3(new_n948), .A4(new_n950), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n713), .A2(G317), .B1(G303), .B2(new_n723), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n714), .A2(G322), .B1(G311), .B2(new_n719), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(KEYINPUT116), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n953), .A2(KEYINPUT116), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n952), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT48), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n958), .B1(new_n532), .B2(new_n716), .C1(new_n469), .C2(new_n728), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT49), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n709), .A2(G326), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n742), .A2(G116), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n961), .A2(new_n414), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n959), .A2(new_n960), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n951), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n705), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n694), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n939), .B1(new_n240), .B2(G45), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n655), .B2(new_n748), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n264), .A2(new_n214), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT50), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n218), .A2(new_n350), .ZN(new_n973));
  NOR4_X1   g0773(.A1(new_n972), .A2(new_n655), .A3(G45), .A4(new_n973), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n970), .A2(new_n974), .B1(G107), .B2(new_n232), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n943), .B(new_n968), .C1(new_n754), .C2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(new_n693), .B2(new_n905), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n907), .A2(new_n909), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n688), .B2(new_n905), .ZN(new_n979));
  INV_X1    g0779(.A(new_n657), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n977), .B1(new_n979), .B2(new_n980), .ZN(G393));
  NAND2_X1  g0781(.A1(new_n878), .A2(new_n699), .ZN(new_n982));
  AOI22_X1  g0782(.A1(G311), .A2(new_n713), .B1(new_n714), .B2(G317), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT52), .Z(new_n984));
  NAND2_X1  g0784(.A1(new_n709), .A2(G322), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n984), .B(new_n985), .C1(new_n914), .C2(new_n718), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n716), .A2(new_n220), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n743), .B1(new_n532), .B2(new_n728), .C1(new_n469), .C2(new_n722), .ZN(new_n988));
  NOR4_X1   g0788(.A1(new_n986), .A2(new_n282), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  AOI22_X1  g0789(.A1(G150), .A2(new_n714), .B1(new_n713), .B2(G159), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT51), .Z(new_n991));
  NOR2_X1   g0791(.A1(new_n716), .A2(new_n350), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(new_n201), .B2(new_n719), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n991), .B(new_n993), .C1(new_n265), .C2(new_n722), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n728), .A2(new_n218), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n395), .B1(new_n928), .B2(new_n708), .ZN(new_n996));
  NOR4_X1   g0796(.A1(new_n994), .A2(new_n787), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n705), .B1(new_n989), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n252), .A2(new_n751), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n999), .B(new_n754), .C1(new_n498), .C2(new_n232), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n982), .A2(new_n694), .A3(new_n998), .A4(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n901), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n978), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1004), .A2(new_n657), .A3(new_n910), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT117), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1004), .A2(KEYINPUT117), .A3(new_n657), .A4(new_n910), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1002), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n901), .A2(new_n693), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(G390));
  NAND4_X1  g0811(.A1(new_n684), .A2(new_n685), .A3(G330), .A4(new_n766), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n851), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n1015), .A2(new_n1016), .B1(new_n852), .B2(new_n853), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1016), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n853), .B1(new_n669), .B2(new_n766), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1018), .A2(new_n1019), .A3(new_n1014), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n615), .A2(new_n848), .A3(new_n844), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n616), .B1(new_n597), .B2(new_n602), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n617), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n661), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n626), .A2(new_n667), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n601), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n641), .B(new_n766), .C1(new_n1027), .C2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n853), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1013), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n859), .B(KEYINPUT110), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n826), .B2(new_n834), .ZN(new_n1034));
  OAI21_X1  g0834(.A(KEYINPUT118), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT118), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n861), .B1(new_n823), .B2(new_n813), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1036), .B(new_n1037), .C1(new_n1019), .C2(new_n1013), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n857), .A2(new_n858), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n629), .A2(new_n641), .A3(new_n766), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1013), .B1(new_n1041), .B2(new_n1031), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1040), .B1(new_n1042), .B2(new_n861), .ZN(new_n1043));
  AND3_X1   g0843(.A1(new_n1039), .A2(new_n1043), .A3(new_n1018), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1018), .B1(new_n1039), .B2(new_n1043), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1024), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n851), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1036), .B1(new_n1048), .B2(new_n1037), .ZN(new_n1049));
  NOR3_X1   g0849(.A1(new_n1032), .A2(KEYINPUT118), .A3(new_n1034), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1043), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n1016), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1039), .A2(new_n1043), .A3(new_n1018), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1022), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  AND3_X1   g0855(.A1(new_n1046), .A2(new_n1055), .A3(new_n657), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1052), .A2(new_n693), .A3(new_n1053), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n698), .B1(new_n857), .B2(new_n858), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n793), .A2(new_n264), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n309), .B1(new_n913), .B2(new_n220), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n719), .A2(new_n344), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n498), .B2(new_n722), .C1(new_n927), .C2(new_n532), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1063), .A2(KEYINPUT120), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(KEYINPUT120), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n992), .B(new_n1060), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1066), .B(new_n738), .C1(new_n469), .C2(new_n708), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1067), .A2(new_n778), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(KEYINPUT54), .B(G143), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n722), .A2(new_n1069), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n282), .B1(new_n273), .B2(new_n726), .C1(new_n913), .C2(new_n779), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(G128), .C2(new_n714), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n719), .A2(G137), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G125), .A2(new_n709), .B1(new_n731), .B2(G159), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n728), .A2(new_n269), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .A4(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n773), .B1(new_n1068), .B2(new_n1078), .ZN(new_n1079));
  NOR4_X1   g0879(.A1(new_n1058), .A2(new_n769), .A3(new_n1059), .A4(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1057), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(KEYINPUT121), .B1(new_n1056), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1046), .A2(new_n1055), .A3(new_n657), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1080), .B1(new_n1085), .B2(new_n693), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT121), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1084), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1083), .A2(new_n1088), .ZN(G378));
  OAI21_X1  g0889(.A(new_n370), .B1(new_n606), .B2(new_n607), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n367), .A2(new_n802), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT55), .Z(new_n1092));
  NAND2_X1  g0892(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(KEYINPUT125), .B(KEYINPUT56), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1092), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n370), .B(new_n1095), .C1(new_n606), .C2(new_n607), .ZN(new_n1096));
  AND3_X1   g0896(.A1(new_n1093), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1094), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(G330), .B1(new_n825), .B2(new_n830), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n862), .A2(new_n855), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1100), .B1(new_n854), .B2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n863), .A2(new_n843), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1099), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1101), .A2(new_n1100), .A3(new_n854), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n863), .A2(new_n843), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1106), .A2(new_n697), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n931), .B1(new_n927), .B2(new_n220), .ZN(new_n1111));
  XOR2_X1   g0911(.A(new_n1111), .B(KEYINPUT122), .Z(new_n1112));
  AOI211_X1 g0912(.A(new_n944), .B(new_n1112), .C1(G97), .C2(new_n719), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n726), .A2(new_n247), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n395), .A2(G41), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n587), .B2(new_n722), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1114), .B(new_n1116), .C1(G283), .C2(new_n709), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1113), .B(new_n1117), .C1(new_n250), .C2(new_n913), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT58), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n718), .A2(new_n779), .ZN(new_n1121));
  INV_X1    g0921(.A(G128), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n913), .A2(new_n1122), .B1(new_n728), .B2(new_n1069), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT123), .Z(new_n1124));
  AOI211_X1 g0924(.A(new_n1121), .B(new_n1124), .C1(G137), .C2(new_n723), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n269), .B2(new_n716), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(G125), .B2(new_n714), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n1128));
  XOR2_X1   g0928(.A(new_n1127), .B(new_n1128), .Z(new_n1129));
  AOI211_X1 g0929(.A(G33), .B(G41), .C1(new_n709), .C2(G124), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n726), .B2(new_n735), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1119), .B1(new_n1115), .B2(new_n1120), .C1(new_n1129), .C2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n705), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1110), .A2(new_n694), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n792), .A2(new_n273), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1109), .A2(new_n693), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1055), .A2(new_n1023), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1137), .A2(KEYINPUT57), .A3(new_n1109), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n657), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1055), .A2(new_n1023), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1140), .A2(KEYINPUT57), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1136), .B1(new_n1139), .B2(new_n1141), .ZN(G375));
  NOR2_X1   g0942(.A1(new_n708), .A2(new_n914), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n945), .B1(new_n344), .B2(new_n723), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n282), .B1(new_n714), .B2(G294), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n713), .A2(G283), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G116), .A2(new_n719), .B1(new_n742), .B2(G77), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1143), .B(new_n1148), .C1(G97), .C2(new_n729), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n714), .A2(G132), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n713), .A2(G137), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n723), .A2(G150), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1114), .B1(G159), .B2(new_n729), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n716), .A2(new_n214), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n708), .A2(new_n1122), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n395), .B1(new_n718), .B2(new_n1069), .ZN(new_n1157));
  NOR4_X1   g0957(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n705), .B1(new_n1149), .B2(new_n1158), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n694), .B(new_n1159), .C1(new_n851), .C2(new_n698), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n218), .B2(new_n792), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n1021), .B2(new_n693), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1022), .A2(new_n1017), .A3(new_n1020), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n892), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1162), .B1(new_n1164), .B2(new_n1054), .ZN(G381));
  NAND4_X1  g0965(.A1(new_n1009), .A2(new_n912), .A3(new_n941), .A4(new_n1010), .ZN(new_n1166));
  OR2_X1    g0966(.A1(G393), .A2(G396), .ZN(new_n1167));
  NOR4_X1   g0967(.A1(new_n1166), .A2(G384), .A3(G381), .A4(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n693), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1171), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n980), .B1(new_n1140), .B2(KEYINPUT57), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT57), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1022), .B1(new_n1085), .B2(new_n1054), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1176), .B1(new_n1177), .B2(new_n1172), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1174), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1168), .A2(new_n1170), .A3(new_n1179), .ZN(G407));
  NOR2_X1   g0980(.A1(new_n1168), .A2(new_n639), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1179), .A2(new_n1170), .ZN(new_n1182));
  OAI21_X1  g0982(.A(G213), .B1(new_n1181), .B2(new_n1182), .ZN(G409));
  INV_X1    g0983(.A(G213), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1184), .A2(G343), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(G2897), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT60), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n980), .B1(new_n1163), .B2(new_n1187), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1022), .A2(new_n1017), .A3(new_n1020), .A4(KEYINPUT60), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1188), .A2(new_n1024), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n1162), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1191), .A2(new_n771), .A3(new_n794), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT126), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1190), .A2(G384), .A3(new_n1162), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1193), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1186), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1198));
  OAI211_X1 g0998(.A(G2897), .B(new_n1185), .C1(new_n1198), .C2(KEYINPUT126), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1140), .A2(new_n892), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1169), .B1(new_n1200), .B2(new_n1136), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n1179), .B2(G378), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1197), .B(new_n1199), .C1(new_n1202), .C2(new_n1185), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(KEYINPUT63), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n1202), .A2(new_n1185), .A3(new_n1198), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1084), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1087), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  AND2_X1   g1010(.A1(new_n1200), .A2(new_n1136), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(G375), .A2(new_n1210), .B1(new_n1169), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1185), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1212), .A2(KEYINPUT63), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(G390), .A2(G387), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(G393), .B(G396), .ZN(new_n1217));
  AND3_X1   g1017(.A1(new_n1216), .A2(new_n1166), .A3(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1217), .B1(new_n1216), .B2(new_n1166), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT61), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1215), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1207), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1220), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT62), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1203), .B1(new_n1205), .B2(new_n1225), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1212), .A2(new_n1225), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n1221), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1224), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1223), .A2(new_n1229), .ZN(G405));
  INV_X1    g1030(.A(KEYINPUT127), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1198), .A2(new_n1231), .ZN(new_n1232));
  OR3_X1    g1032(.A1(new_n1218), .A2(new_n1219), .A3(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(G375), .A2(new_n1170), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1179), .A2(G378), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1234), .A2(new_n1235), .B1(new_n1231), .B2(new_n1198), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1232), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n1233), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1236), .B1(new_n1233), .B2(new_n1237), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(G402));
endmodule


