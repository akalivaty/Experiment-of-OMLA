//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1225, new_n1226,
    new_n1227, new_n1228;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  XOR2_X1   g029(.A(G325), .B(KEYINPUT65), .Z(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G125), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g042(.A(G2105), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n470), .B1(G2104), .B2(new_n471), .ZN(new_n472));
  NOR3_X1   g047(.A1(new_n462), .A2(KEYINPUT66), .A3(G2105), .ZN(new_n473));
  OAI21_X1  g048(.A(G101), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(G137), .A3(new_n471), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n469), .A2(new_n477), .ZN(G160));
  AOI21_X1  g053(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n471), .B1(new_n463), .B2(new_n464), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  AND2_X1   g061(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n487));
  NOR2_X1   g062(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n488));
  OAI211_X1 g063(.A(G138), .B(new_n471), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n475), .A2(new_n491), .A3(G138), .A4(new_n471), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT67), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n471), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n498), .A2(new_n500), .A3(KEYINPUT67), .A4(G2104), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n481), .A2(G126), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n493), .A2(new_n504), .ZN(G164));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(KEYINPUT68), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT68), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(KEYINPUT5), .A3(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G62), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n518), .B1(new_n508), .B2(new_n510), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n519), .A2(KEYINPUT69), .ZN(new_n520));
  NAND2_X1  g095(.A1(G75), .A2(G543), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n521), .B1(new_n519), .B2(KEYINPUT69), .ZN(new_n522));
  OAI21_X1  g097(.A(G651), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT70), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n517), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI211_X1 g100(.A(KEYINPUT70), .B(G651), .C1(new_n520), .C2(new_n522), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(G166));
  AND2_X1   g102(.A1(new_n512), .A2(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n529), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n511), .A2(new_n512), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n534), .A2(G89), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n533), .A2(new_n535), .ZN(G168));
  AOI22_X1  g111(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  INV_X1    g112(.A(G651), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n513), .A2(new_n540), .B1(new_n515), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(G171));
  XOR2_X1   g118(.A(KEYINPUT71), .B(G81), .Z(new_n544));
  NAND2_X1  g119(.A1(new_n534), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n528), .A2(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n538), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  XOR2_X1   g130(.A(KEYINPUT72), .B(KEYINPUT9), .Z(new_n556));
  NAND3_X1  g131(.A1(new_n528), .A2(G53), .A3(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n558));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n515), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n511), .A2(G91), .A3(new_n512), .ZN(new_n561));
  AND3_X1   g136(.A1(new_n557), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n563), .B1(new_n508), .B2(new_n510), .ZN(new_n564));
  AND2_X1   g139(.A1(G78), .A2(G543), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT73), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g143(.A(KEYINPUT73), .B(G651), .C1(new_n564), .C2(new_n565), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n562), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(G168), .ZN(G286));
  NAND2_X1  g148(.A1(new_n525), .A2(new_n526), .ZN(G303));
  OAI21_X1  g149(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n512), .A2(G49), .A3(G543), .ZN(new_n576));
  INV_X1    g151(.A(G87), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n575), .B(new_n576), .C1(new_n577), .C2(new_n513), .ZN(G288));
  INV_X1    g153(.A(G86), .ZN(new_n579));
  INV_X1    g154(.A(G48), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n513), .A2(new_n579), .B1(new_n515), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n582), .B1(new_n508), .B2(new_n510), .ZN(new_n583));
  AND2_X1   g158(.A1(G73), .A2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT74), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g162(.A(KEYINPUT74), .B(G651), .C1(new_n583), .C2(new_n584), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n581), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G305));
  AOI22_X1  g165(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n538), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n528), .A2(G47), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n511), .A2(G85), .A3(new_n512), .ZN(new_n595));
  AND3_X1   g170(.A1(new_n594), .A2(KEYINPUT75), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(KEYINPUT75), .B1(new_n594), .B2(new_n595), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n593), .B1(new_n596), .B2(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT76), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(new_n534), .B2(G92), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  NOR3_X1   g178(.A1(new_n513), .A2(KEYINPUT76), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n600), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT77), .Z(new_n607));
  NAND2_X1  g182(.A1(new_n511), .A2(G66), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n538), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(G54), .B2(new_n528), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n534), .A2(new_n601), .A3(G92), .ZN(new_n611));
  OAI21_X1  g186(.A(KEYINPUT76), .B1(new_n513), .B2(new_n603), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n611), .A2(KEYINPUT10), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n605), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n599), .B1(new_n615), .B2(G868), .ZN(G284));
  OAI21_X1  g191(.A(new_n599), .B1(new_n615), .B2(G868), .ZN(G321));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  NOR2_X1   g193(.A1(G286), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(G299), .B(KEYINPUT78), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(new_n618), .ZN(G297));
  AOI21_X1  g196(.A(new_n619), .B1(new_n620), .B2(new_n618), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n615), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n615), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g203(.A1(new_n472), .A2(new_n473), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(new_n475), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT12), .Z(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT13), .Z(new_n632));
  INV_X1    g207(.A(G2100), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  INV_X1    g211(.A(G111), .ZN(new_n637));
  AOI22_X1  g212(.A1(new_n636), .A2(KEYINPUT79), .B1(new_n637), .B2(G2105), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(KEYINPUT79), .B2(new_n636), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n479), .A2(G135), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n481), .A2(G123), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2096), .Z(new_n643));
  NAND3_X1  g218(.A1(new_n634), .A2(new_n635), .A3(new_n643), .ZN(G156));
  INV_X1    g219(.A(KEYINPUT14), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2427), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2430), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n649), .B1(new_n648), .B2(new_n647), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n650), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(new_n658), .A3(G14), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT80), .Z(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G401));
  XOR2_X1   g236(.A(KEYINPUT81), .B(KEYINPUT18), .Z(new_n662));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g240(.A1(new_n665), .A2(KEYINPUT17), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n663), .A2(new_n664), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n662), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2072), .B(G2078), .Z(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n665), .B2(new_n662), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n668), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2096), .B(G2100), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT20), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n676), .A2(new_n677), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n675), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(new_n675), .B2(new_n681), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1991), .B(G1996), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT82), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n686), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n689), .B(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(G229));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G21), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G168), .B2(new_n694), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G1966), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT93), .B(KEYINPUT31), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G11), .ZN(new_n699));
  INV_X1    g274(.A(G28), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n700), .A2(KEYINPUT30), .ZN(new_n701));
  AOI21_X1  g276(.A(G29), .B1(new_n700), .B2(KEYINPUT30), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n699), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n697), .B(new_n703), .C1(new_n704), .C2(new_n642), .ZN(new_n705));
  NOR2_X1   g280(.A1(G171), .A2(new_n694), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G5), .B2(new_n694), .ZN(new_n707));
  INV_X1    g282(.A(G1961), .ZN(new_n708));
  OAI22_X1  g283(.A1(new_n707), .A2(new_n708), .B1(new_n696), .B2(G1966), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT94), .ZN(new_n710));
  OR3_X1    g285(.A1(new_n705), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(G162), .A2(G29), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G29), .B2(G35), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT29), .B(G2090), .Z(new_n714));
  AND2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n704), .A2(G33), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n475), .A2(G127), .ZN(new_n717));
  NAND2_X1  g292(.A1(G115), .A2(G2104), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(G2105), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT25), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n723), .A2(new_n724), .B1(new_n479), .B2(G139), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n720), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n716), .B1(new_n726), .B2(G29), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(G2072), .Z(new_n728));
  INV_X1    g303(.A(G2084), .ZN(new_n729));
  NAND2_X1  g304(.A1(G160), .A2(G29), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT24), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n731), .A2(G34), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n704), .B1(new_n731), .B2(G34), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n730), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AOI211_X1 g309(.A(new_n715), .B(new_n728), .C1(new_n729), .C2(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n734), .A2(new_n729), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n704), .A2(G32), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT92), .B(KEYINPUT26), .Z(new_n738));
  NAND3_X1  g313(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n481), .A2(G129), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n629), .A2(G105), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n479), .A2(G141), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n740), .A2(new_n741), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n737), .B1(new_n744), .B2(G29), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT27), .B(G1996), .ZN(new_n746));
  OAI22_X1  g321(.A1(new_n713), .A2(new_n714), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AOI211_X1 g322(.A(new_n736), .B(new_n747), .C1(new_n745), .C2(new_n746), .ZN(new_n748));
  NOR2_X1   g323(.A1(G27), .A2(G29), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G164), .B2(G29), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n707), .A2(new_n708), .B1(new_n750), .B2(G2078), .ZN(new_n751));
  AND4_X1   g326(.A1(new_n711), .A2(new_n735), .A3(new_n748), .A4(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n710), .B1(new_n705), .B2(new_n709), .ZN(new_n753));
  NOR2_X1   g328(.A1(G4), .A2(G16), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n615), .B2(G16), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT90), .B(G1348), .Z(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT89), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n755), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n704), .A2(G26), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT28), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n479), .A2(G140), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n481), .A2(G128), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n471), .A2(G116), .ZN(new_n763));
  OAI21_X1  g338(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n761), .B(new_n762), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT91), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n760), .B1(new_n769), .B2(G29), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2067), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT95), .B(G1956), .Z(new_n772));
  NAND2_X1  g347(.A1(G299), .A2(G16), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n694), .A2(G20), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT23), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n771), .B1(new_n772), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(G16), .A2(G19), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n550), .B2(G16), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(G1341), .Z(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G2078), .B2(new_n750), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n776), .A2(new_n772), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n777), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n752), .A2(new_n753), .A3(new_n758), .A4(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(G290), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(G16), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G16), .B2(G24), .ZN(new_n788));
  INV_X1    g363(.A(G1986), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OR2_X1    g365(.A1(G95), .A2(G2105), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n791), .B(G2104), .C1(G107), .C2(new_n471), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT83), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n479), .A2(G131), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n481), .A2(G119), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n796), .A2(new_n704), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G25), .B2(G29), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT35), .B(G1991), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT84), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n800), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n797), .B(new_n802), .C1(G25), .C2(G29), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n787), .B(G1986), .C1(G16), .C2(G24), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n790), .A2(new_n804), .A3(KEYINPUT88), .A4(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n525), .A2(G16), .A3(new_n526), .ZN(new_n807));
  OR2_X1    g382(.A1(G16), .A2(G22), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(G1971), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n807), .A2(G1971), .A3(new_n808), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n694), .A2(G23), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G288), .B2(G16), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT33), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI211_X1 g391(.A(KEYINPUT33), .B(new_n813), .C1(G288), .C2(G16), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n816), .A2(new_n818), .A3(G1976), .ZN(new_n819));
  INV_X1    g394(.A(G1976), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n814), .A2(new_n815), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(new_n817), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n811), .A2(new_n812), .A3(new_n819), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n694), .A2(G6), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n589), .B2(new_n694), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(KEYINPUT85), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT85), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n827), .B(new_n824), .C1(new_n589), .C2(new_n694), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT32), .B(G1981), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT86), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n831), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n826), .A2(new_n833), .A3(new_n828), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n823), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT34), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n806), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n812), .A2(new_n819), .A3(new_n822), .ZN(new_n838));
  AOI21_X1  g413(.A(G1971), .B1(new_n807), .B2(new_n808), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n832), .A2(new_n834), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(KEYINPUT87), .B1(new_n842), .B2(KEYINPUT34), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT87), .ZN(new_n844));
  AOI211_X1 g419(.A(new_n844), .B(new_n836), .C1(new_n840), .C2(new_n841), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n837), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(KEYINPUT36), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT36), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n837), .B(new_n848), .C1(new_n843), .C2(new_n845), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n785), .B1(new_n847), .B2(new_n849), .ZN(G311));
  NAND2_X1  g425(.A1(new_n847), .A2(new_n849), .ZN(new_n851));
  INV_X1    g426(.A(new_n785), .ZN(new_n852));
  AOI21_X1  g427(.A(KEYINPUT96), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT96), .ZN(new_n854));
  AOI211_X1 g429(.A(new_n854), .B(new_n785), .C1(new_n847), .C2(new_n849), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n853), .A2(new_n855), .ZN(G150));
  INV_X1    g431(.A(new_n549), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n857), .A2(KEYINPUT98), .A3(new_n546), .A4(new_n545), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT98), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n859), .B1(new_n547), .B2(new_n549), .ZN(new_n860));
  AOI22_X1  g435(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n861), .A2(new_n538), .ZN(new_n862));
  INV_X1    g437(.A(G93), .ZN(new_n863));
  XOR2_X1   g438(.A(KEYINPUT97), .B(G55), .Z(new_n864));
  OAI22_X1  g439(.A1(new_n513), .A2(new_n863), .B1(new_n515), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n858), .A2(new_n860), .A3(new_n866), .ZN(new_n867));
  OAI221_X1 g442(.A(new_n859), .B1(new_n862), .B2(new_n865), .C1(new_n547), .C2(new_n549), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT38), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n614), .A2(new_n623), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n872), .A2(KEYINPUT39), .ZN(new_n873));
  INV_X1    g448(.A(G860), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(KEYINPUT39), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n866), .A2(new_n874), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT37), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(G145));
  XOR2_X1   g454(.A(KEYINPUT101), .B(G37), .Z(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n631), .B(new_n796), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n481), .A2(G130), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n471), .A2(G118), .ZN(new_n884));
  OAI21_X1  g459(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n475), .A2(new_n471), .ZN(new_n887));
  INV_X1    g462(.A(G142), .ZN(new_n888));
  OR3_X1    g463(.A1(new_n887), .A2(KEYINPUT99), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT99), .B1(new_n887), .B2(new_n888), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n886), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n882), .B(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n726), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n767), .A2(G164), .A3(new_n768), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(G164), .B1(new_n767), .B2(new_n768), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n893), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NOR3_X1   g473(.A1(new_n895), .A2(new_n893), .A3(new_n896), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n744), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n899), .ZN(new_n901));
  INV_X1    g476(.A(new_n744), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n902), .A3(new_n897), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n892), .A2(new_n900), .A3(new_n903), .A4(KEYINPUT102), .ZN(new_n904));
  XNOR2_X1  g479(.A(G160), .B(G162), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(new_n642), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n892), .A2(new_n900), .A3(new_n903), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT100), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n900), .A2(new_n903), .ZN(new_n913));
  INV_X1    g488(.A(new_n892), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n913), .A2(new_n914), .A3(new_n912), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n881), .B1(new_n911), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n917), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n910), .B1(new_n920), .B2(new_n915), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n906), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n919), .A2(KEYINPUT40), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT40), .B1(new_n919), .B2(new_n922), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(G395));
  OAI21_X1  g500(.A(new_n618), .B1(new_n862), .B2(new_n865), .ZN(new_n926));
  INV_X1    g501(.A(G288), .ZN(new_n927));
  XNOR2_X1  g502(.A(G290), .B(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(G303), .A2(new_n589), .ZN(new_n929));
  AOI21_X1  g504(.A(G305), .B1(new_n526), .B2(new_n525), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(G290), .B(G288), .ZN(new_n932));
  NAND2_X1  g507(.A1(G166), .A2(G305), .ZN(new_n933));
  INV_X1    g508(.A(new_n930), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT42), .B1(new_n931), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT103), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n931), .A2(new_n935), .A3(KEYINPUT103), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n936), .B1(new_n942), .B2(KEYINPUT42), .ZN(new_n943));
  OR2_X1    g518(.A1(new_n614), .A2(G299), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n614), .A2(G299), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT41), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n944), .A2(KEYINPUT41), .A3(new_n945), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n946), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n625), .B(new_n869), .ZN(new_n952));
  MUX2_X1   g527(.A(new_n950), .B(new_n951), .S(new_n952), .Z(new_n953));
  XNOR2_X1  g528(.A(new_n943), .B(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n926), .B1(new_n954), .B2(new_n618), .ZN(G295));
  OAI21_X1  g530(.A(new_n926), .B1(new_n954), .B2(new_n618), .ZN(G331));
  OAI21_X1  g531(.A(KEYINPUT104), .B1(new_n533), .B2(new_n535), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n530), .A2(new_n532), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n534), .A2(G89), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n958), .A2(new_n959), .A3(new_n960), .A4(new_n529), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n957), .A2(G301), .A3(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(G168), .A2(G171), .A3(new_n960), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n869), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n867), .A2(new_n962), .A3(new_n868), .A4(new_n963), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n948), .A2(new_n967), .A3(new_n949), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n951), .A2(new_n966), .A3(new_n965), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n931), .A2(new_n935), .A3(KEYINPUT103), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT103), .B1(new_n931), .B2(new_n935), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G37), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n940), .A2(new_n941), .A3(new_n968), .A4(new_n969), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n970), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n971), .A2(new_n972), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT43), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n881), .B1(new_n942), .B2(new_n970), .ZN(new_n980));
  AOI22_X1  g555(.A1(new_n976), .A2(KEYINPUT43), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT105), .B1(new_n981), .B2(KEYINPUT44), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT105), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT44), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n979), .A2(new_n980), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n986));
  AOI21_X1  g561(.A(G37), .B1(new_n942), .B2(new_n970), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n986), .B1(new_n987), .B2(new_n975), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n983), .B(new_n984), .C1(new_n985), .C2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n984), .B1(new_n979), .B2(new_n987), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n973), .A2(new_n880), .A3(new_n975), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n990), .A2(new_n992), .A3(KEYINPUT106), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT106), .B1(new_n990), .B2(new_n992), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n982), .B(new_n989), .C1(new_n993), .C2(new_n994), .ZN(G397));
  XNOR2_X1  g570(.A(new_n769), .B(G2067), .ZN(new_n996));
  INV_X1    g571(.A(G1384), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(new_n493), .B2(new_n504), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT45), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n468), .A2(G40), .A3(new_n474), .A4(new_n476), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1002), .B(KEYINPUT107), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n996), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n996), .A2(new_n1003), .A3(KEYINPUT108), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1003), .A2(new_n744), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1002), .ZN(new_n1009));
  INV_X1    g584(.A(G1996), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n744), .A2(new_n1010), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n1006), .A2(new_n1007), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n799), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n796), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n796), .A2(new_n1015), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1003), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g594(.A(G290), .B(G1986), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1019), .B1(new_n1009), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G1981), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n589), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n589), .A2(new_n1022), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT113), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1025), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(new_n1028), .A3(new_n1023), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT49), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1026), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n998), .A2(new_n1000), .ZN(new_n1032));
  XOR2_X1   g607(.A(KEYINPUT111), .B(G8), .Z(new_n1033));
  NOR2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT114), .B1(new_n1035), .B2(KEYINPUT49), .ZN(new_n1036));
  AND4_X1   g611(.A1(KEYINPUT114), .A2(new_n1027), .A3(KEYINPUT49), .A4(new_n1023), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1031), .B(new_n1034), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1034), .B1(new_n820), .B2(G288), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1039), .B1(KEYINPUT112), .B2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1040), .A2(KEYINPUT112), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1034), .B(new_n1042), .C1(new_n820), .C2(G288), .ZN(new_n1043));
  NAND3_X1  g618(.A1(G288), .A2(new_n1040), .A3(new_n820), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1041), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n1038), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT116), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1038), .A2(new_n1045), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n490), .A2(new_n492), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n497), .A2(new_n501), .B1(new_n481), .B2(G126), .ZN(new_n1052));
  AOI21_X1  g627(.A(G1384), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT50), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1001), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1056), .B(KEYINPUT115), .C1(G164), .C2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G2090), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n1061));
  NOR2_X1   g636(.A1(G164), .A2(new_n1058), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1061), .B1(new_n1055), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1059), .A2(new_n1060), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1000), .B1(new_n1053), .B2(KEYINPUT45), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n998), .A2(new_n999), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n810), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1033), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G8), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1070), .B1(new_n525), .B2(new_n526), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT110), .ZN(new_n1072));
  OR3_X1    g647(.A1(new_n1071), .A2(new_n1072), .A3(KEYINPUT55), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(KEYINPUT55), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1072), .B1(new_n1071), .B2(KEYINPUT55), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  OR2_X1    g651(.A1(new_n1069), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT109), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1078), .B1(new_n1079), .B2(new_n1057), .ZN(new_n1080));
  AOI211_X1 g655(.A(KEYINPUT109), .B(new_n1058), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1082), .A2(new_n1055), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n1060), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1070), .B1(new_n1084), .B2(new_n1068), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1076), .A2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1047), .A2(new_n1050), .A3(new_n1077), .A4(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT109), .B1(G164), .B2(new_n1058), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1079), .A2(new_n1078), .A3(new_n1057), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1090), .A2(new_n729), .A3(new_n1056), .ZN(new_n1091));
  INV_X1    g666(.A(G1966), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1067), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1033), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(G168), .A2(new_n1033), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1097), .A2(KEYINPUT51), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1082), .A2(G2084), .A3(new_n1055), .ZN(new_n1100));
  AOI21_X1  g675(.A(G1966), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1101));
  OAI211_X1 g676(.A(G286), .B(new_n1095), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT51), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1097), .B1(new_n1094), .B2(G8), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1099), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(G2078), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1065), .A2(new_n1066), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT121), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1065), .A2(new_n1066), .A3(new_n1109), .A4(new_n1106), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1108), .A2(KEYINPUT53), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1107), .A2(KEYINPUT122), .A3(new_n1112), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1090), .A2(new_n1056), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n708), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1111), .A2(new_n1115), .A3(new_n1116), .A4(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(G171), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1114), .A2(new_n1113), .B1(new_n1117), .B2(new_n708), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1121), .A2(G301), .A3(new_n1116), .A4(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1120), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1105), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1115), .A2(new_n1118), .A3(new_n1116), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1128), .A2(G301), .A3(new_n1111), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1115), .A2(new_n1118), .A3(new_n1116), .ZN(new_n1131));
  OAI21_X1  g706(.A(G171), .B1(new_n1131), .B2(new_n1122), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1129), .A2(new_n1130), .A3(new_n1132), .A4(KEYINPUT54), .ZN(new_n1133));
  INV_X1    g708(.A(G1956), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n1055), .B2(new_n1062), .ZN(new_n1135));
  XOR2_X1   g710(.A(KEYINPUT56), .B(G2072), .Z(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(KEYINPUT119), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1065), .A2(new_n1066), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT118), .ZN(new_n1139));
  NAND3_X1  g714(.A1(G299), .A2(new_n1139), .A3(KEYINPUT57), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(KEYINPUT57), .ZN(new_n1141));
  OR2_X1    g716(.A1(new_n1139), .A2(KEYINPUT57), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n562), .A2(new_n570), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1135), .A2(new_n1138), .A3(new_n1140), .A4(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n756), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1145), .B1(new_n1090), .B2(new_n1056), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n998), .A2(G2067), .A3(new_n1000), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n614), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n1135), .A2(new_n1138), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1144), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT60), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1153), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1154));
  OAI211_X1 g729(.A(KEYINPUT60), .B(new_n1149), .C1(new_n1083), .C2(new_n1145), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1154), .A2(new_n615), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1157), .B1(new_n1160), .B2(new_n1151), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1151), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1162), .A2(KEYINPUT61), .A3(new_n1144), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1156), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g739(.A(KEYINPUT58), .B(G1341), .ZN(new_n1165));
  OAI22_X1  g740(.A1(new_n1067), .A2(G1996), .B1(new_n1032), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(new_n550), .ZN(new_n1167));
  NAND2_X1  g742(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1166), .A2(KEYINPUT120), .A3(KEYINPUT59), .A4(new_n550), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1169), .B(new_n1170), .C1(new_n615), .C2(new_n1155), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1152), .B1(new_n1164), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(G301), .B1(new_n1128), .B2(new_n1123), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1111), .A2(G301), .ZN(new_n1174));
  OAI21_X1  g749(.A(KEYINPUT54), .B1(new_n1131), .B2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(KEYINPUT123), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1127), .A2(new_n1133), .A3(new_n1172), .A4(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1120), .B1(new_n1105), .B2(new_n1178), .ZN(new_n1179));
  OAI211_X1 g754(.A(new_n1099), .B(KEYINPUT62), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT63), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1096), .A2(G286), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n1179), .A2(new_n1180), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1087), .B1(new_n1177), .B2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1048), .A2(new_n1086), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1038), .A2(new_n820), .A3(new_n927), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(new_n1023), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1185), .B1(new_n1034), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1086), .A2(new_n1182), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1076), .A2(new_n1085), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT117), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1046), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  OAI21_X1  g768(.A(KEYINPUT117), .B1(new_n1048), .B2(new_n1190), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1189), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1188), .B1(new_n1195), .B2(new_n1181), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1021), .B1(new_n1184), .B2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1009), .A2(new_n786), .A3(new_n789), .ZN(new_n1198));
  XNOR2_X1  g773(.A(new_n1198), .B(KEYINPUT48), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1199), .B1(new_n1019), .B2(KEYINPUT127), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT127), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1201), .B1(new_n1014), .B2(new_n1018), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1003), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n769), .A2(G2067), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1204), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1205));
  OAI22_X1  g780(.A1(new_n1200), .A2(new_n1202), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1004), .A2(new_n1008), .ZN(new_n1207));
  OR2_X1    g782(.A1(new_n1207), .A2(KEYINPUT125), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1207), .A2(KEYINPUT125), .ZN(new_n1209));
  NOR2_X1   g784(.A1(KEYINPUT124), .A2(KEYINPUT46), .ZN(new_n1210));
  NOR2_X1   g785(.A1(new_n1011), .A2(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g786(.A(KEYINPUT124), .B(KEYINPUT46), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1211), .B1(new_n1011), .B2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1208), .A2(new_n1209), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1214), .A2(KEYINPUT126), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT126), .ZN(new_n1216));
  NAND4_X1  g791(.A1(new_n1208), .A2(new_n1216), .A3(new_n1209), .A4(new_n1213), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1218), .A2(KEYINPUT47), .ZN(new_n1219));
  INV_X1    g794(.A(KEYINPUT47), .ZN(new_n1220));
  NAND3_X1  g795(.A1(new_n1215), .A2(new_n1220), .A3(new_n1217), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n1206), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1197), .A2(new_n1222), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g798(.A1(G227), .A2(new_n458), .ZN(new_n1225));
  NOR3_X1   g799(.A1(G229), .A2(G401), .A3(new_n1225), .ZN(new_n1226));
  NAND2_X1  g800(.A1(new_n919), .A2(new_n922), .ZN(new_n1227));
  INV_X1    g801(.A(new_n981), .ZN(new_n1228));
  AND3_X1   g802(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .ZN(G308));
  NAND3_X1  g803(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .ZN(G225));
endmodule


