//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 0 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(G137), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT67), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G137), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT11), .A2(G134), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT68), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT68), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n189), .A2(new_n191), .A3(new_n192), .A4(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G131), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT11), .ZN(new_n199));
  INV_X1    g013(.A(G134), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(G137), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  OAI211_X1 g017(.A(KEYINPUT66), .B(new_n199), .C1(new_n200), .C2(G137), .ZN(new_n204));
  AOI22_X1  g018(.A1(new_n203), .A2(new_n204), .B1(new_n200), .B2(G137), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n197), .A2(new_n198), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT65), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n208), .A2(new_n210), .A3(G143), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  INV_X1    g027(.A(G128), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(KEYINPUT1), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n211), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n214), .B1(new_n211), .B2(KEYINPUT1), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n212), .A2(G146), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n208), .A2(new_n210), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n218), .B1(new_n219), .B2(new_n212), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n216), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT67), .B(G137), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(G134), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n200), .A2(G137), .ZN(new_n224));
  OAI21_X1  g038(.A(G131), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n206), .A2(new_n221), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT71), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AND2_X1   g042(.A1(KEYINPUT0), .A2(G128), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n211), .A2(new_n213), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n230), .B1(new_n220), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n197), .A2(new_n198), .A3(new_n205), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n198), .B1(new_n197), .B2(new_n205), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n206), .A2(new_n221), .A3(KEYINPUT71), .A4(new_n225), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n228), .A2(new_n238), .A3(KEYINPUT30), .A4(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n195), .B1(new_n222), .B2(new_n192), .ZN(new_n242));
  AND4_X1   g056(.A1(new_n195), .A2(new_n189), .A3(new_n191), .A4(new_n192), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n203), .A2(new_n204), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n200), .A2(G137), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(G131), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n234), .B1(new_n248), .B2(new_n206), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n206), .A2(new_n221), .A3(new_n225), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n241), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G116), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(G119), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT70), .B(G116), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n253), .B1(new_n254), .B2(G119), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT2), .ZN(new_n257));
  INV_X1    g071(.A(G113), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT69), .B1(KEYINPUT2), .B2(G113), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(KEYINPUT2), .A2(G113), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n255), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n255), .B1(new_n261), .B2(new_n262), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n240), .A2(new_n251), .A3(new_n266), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n228), .A2(new_n238), .A3(new_n265), .A4(new_n239), .ZN(new_n268));
  INV_X1    g082(.A(G237), .ZN(new_n269));
  INV_X1    g083(.A(G953), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n270), .A3(G210), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n271), .B(KEYINPUT27), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT26), .B(G101), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n272), .B(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT31), .B1(new_n267), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n238), .A2(new_n265), .A3(new_n226), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT28), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n265), .B1(new_n238), .B2(new_n226), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n279), .B(new_n281), .C1(new_n278), .C2(new_n268), .ZN(new_n282));
  INV_X1    g096(.A(new_n274), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n276), .A2(new_n284), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n268), .A2(new_n274), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n240), .A2(new_n251), .A3(new_n266), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT31), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n286), .A2(new_n287), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n286), .A2(new_n289), .A3(new_n288), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT72), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n285), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(G472), .A2(G902), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n187), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n228), .A2(new_n238), .A3(new_n239), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n266), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n268), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT28), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT73), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n277), .A2(new_n301), .A3(new_n278), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n301), .B1(new_n277), .B2(new_n278), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT29), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n283), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n300), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT74), .ZN(new_n308));
  OR2_X1    g122(.A1(new_n268), .A2(new_n278), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n280), .B1(new_n278), .B2(new_n277), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n283), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n288), .A2(new_n268), .A3(new_n283), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n305), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G902), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT74), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n300), .A2(new_n304), .A3(new_n315), .A4(new_n306), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n308), .A2(new_n313), .A3(new_n314), .A4(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G472), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n292), .A2(new_n290), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n286), .A2(new_n288), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n320), .A2(KEYINPUT31), .B1(new_n282), .B2(new_n283), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(KEYINPUT32), .A3(new_n294), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n296), .A2(new_n318), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n296), .A2(new_n318), .A3(KEYINPUT75), .A4(new_n323), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G217), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n329), .B1(G234), .B2(new_n314), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n214), .B(G119), .C1(KEYINPUT77), .C2(KEYINPUT23), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT23), .ZN(new_n332));
  INV_X1    g146(.A(G119), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n332), .B1(new_n333), .B2(G128), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n335), .B1(new_n333), .B2(G128), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n331), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT78), .B1(new_n337), .B2(G110), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT23), .B1(new_n214), .B2(G119), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n339), .B(new_n335), .C1(new_n333), .C2(G128), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n341));
  INV_X1    g155(.A(G110), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n340), .A2(new_n341), .A3(new_n342), .A4(new_n331), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT24), .B(G110), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n344), .B(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(G119), .B(G128), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n338), .B(new_n343), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT16), .ZN(new_n349));
  INV_X1    g163(.A(G140), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n350), .A3(G125), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(G125), .ZN(new_n352));
  INV_X1    g166(.A(G125), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G140), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n351), .B1(new_n355), .B2(new_n349), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n356), .A2(new_n207), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n219), .A2(new_n355), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n348), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n346), .A2(new_n347), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n337), .A2(G110), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n356), .A2(new_n207), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n361), .B(new_n362), .C1(new_n363), .C2(new_n357), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT80), .B1(new_n360), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n270), .A2(G221), .A3(G234), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n366), .B(KEYINPUT79), .ZN(new_n367));
  XNOR2_X1  g181(.A(KEYINPUT22), .B(G137), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n367), .B(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n360), .A2(new_n364), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT80), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n360), .A2(new_n364), .A3(KEYINPUT80), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n370), .B1(new_n375), .B2(new_n369), .ZN(new_n376));
  AOI21_X1  g190(.A(KEYINPUT25), .B1(new_n376), .B2(new_n314), .ZN(new_n377));
  INV_X1    g191(.A(new_n369), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n378), .B1(new_n373), .B2(new_n374), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT25), .ZN(new_n380));
  NOR4_X1   g194(.A1(new_n379), .A2(new_n370), .A3(new_n380), .A4(G902), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n330), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n330), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n314), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n385), .B(KEYINPUT81), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n376), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(KEYINPUT9), .B(G234), .ZN(new_n389));
  OAI21_X1  g203(.A(G221), .B1(new_n389), .B2(G902), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(G110), .B(G140), .ZN(new_n392));
  INV_X1    g206(.A(G227), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n393), .A2(G953), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n392), .B(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G104), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT82), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G104), .ZN(new_n399));
  INV_X1    g213(.A(G107), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n397), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n401), .B(G101), .C1(new_n396), .C2(new_n400), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n397), .B(new_n399), .C1(KEYINPUT3), .C2(G107), .ZN(new_n403));
  AND2_X1   g217(.A1(KEYINPUT3), .A2(G107), .ZN(new_n404));
  NOR2_X1   g218(.A1(KEYINPUT3), .A2(G107), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n404), .B1(G104), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G101), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n403), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n402), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT10), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n221), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n407), .B1(new_n403), .B2(new_n406), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT83), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n414), .B1(new_n413), .B2(new_n415), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n408), .A2(KEYINPUT4), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n235), .B1(new_n413), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n412), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n211), .A2(new_n213), .A3(new_n215), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT1), .B1(new_n212), .B2(G146), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n211), .A2(new_n213), .B1(G128), .B2(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT84), .B1(new_n425), .B2(new_n409), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n402), .A2(new_n408), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n211), .A2(new_n213), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n423), .A2(G128), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n216), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT84), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n427), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(KEYINPUT10), .B1(new_n426), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n236), .A2(new_n237), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n421), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  NOR3_X1   g250(.A1(new_n425), .A2(new_n409), .A3(KEYINPUT84), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n431), .B1(new_n427), .B2(new_n430), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n410), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n408), .A2(KEYINPUT4), .ZN(new_n440));
  INV_X1    g254(.A(new_n413), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n234), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n403), .A2(new_n406), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(new_n415), .A3(G101), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(KEYINPUT83), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n442), .A2(new_n447), .B1(new_n221), .B2(new_n411), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n434), .B1(new_n439), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n395), .B1(new_n436), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT12), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n437), .A2(new_n438), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n427), .A2(new_n221), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n451), .B(new_n435), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n439), .A2(new_n448), .A3(new_n434), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n453), .B1(new_n432), .B2(new_n426), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT12), .B1(new_n456), .B2(new_n434), .ZN(new_n457));
  INV_X1    g271(.A(new_n395), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n454), .A2(new_n455), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  AOI211_X1 g273(.A(G469), .B(G902), .C1(new_n450), .C2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G469), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(new_n314), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n395), .ZN(new_n465));
  INV_X1    g279(.A(new_n449), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n455), .A3(new_n458), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n467), .A3(G469), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n391), .B1(new_n463), .B2(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT90), .B(KEYINPUT20), .ZN(new_n470));
  XNOR2_X1  g284(.A(G113), .B(G122), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(new_n396), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n269), .A2(new_n270), .A3(G214), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n212), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n269), .A2(new_n270), .A3(G143), .A4(G214), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(KEYINPUT18), .A2(G131), .ZN(new_n477));
  XOR2_X1   g291(.A(new_n476), .B(new_n477), .Z(new_n478));
  XNOR2_X1  g292(.A(new_n355), .B(KEYINPUT91), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n358), .B1(new_n479), .B2(G146), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n356), .B(new_n207), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n476), .A2(KEYINPUT17), .A3(G131), .ZN(new_n484));
  OR2_X1    g298(.A1(new_n484), .A2(KEYINPUT92), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(KEYINPUT92), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT93), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n476), .B(G131), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n491), .A2(KEYINPUT17), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(new_n487), .B2(new_n488), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n472), .B(new_n482), .C1(new_n490), .C2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n479), .A2(KEYINPUT19), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n496), .B1(KEYINPUT19), .B2(new_n355), .ZN(new_n497));
  OAI221_X1 g311(.A(new_n491), .B1(new_n207), .B2(new_n356), .C1(new_n497), .C2(new_n219), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n482), .ZN(new_n499));
  INV_X1    g313(.A(new_n472), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(G475), .A2(G902), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n470), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n503), .ZN(new_n505));
  AOI211_X1 g319(.A(KEYINPUT20), .B(new_n505), .C1(new_n495), .C2(new_n501), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n482), .B1(new_n490), .B2(new_n494), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n500), .ZN(new_n508));
  AOI21_X1  g322(.A(G902), .B1(new_n508), .B2(new_n495), .ZN(new_n509));
  INV_X1    g323(.A(G475), .ZN(new_n510));
  OAI22_X1  g324(.A1(new_n504), .A2(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(G128), .B(G143), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(G134), .ZN(new_n514));
  AOI211_X1 g328(.A(KEYINPUT13), .B(new_n200), .C1(new_n214), .C2(G143), .ZN(new_n515));
  OR2_X1    g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n515), .ZN(new_n517));
  AND2_X1   g331(.A1(KEYINPUT94), .A2(G122), .ZN(new_n518));
  NOR2_X1   g332(.A1(KEYINPUT94), .A2(G122), .ZN(new_n519));
  OAI21_X1  g333(.A(G116), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT95), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT95), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n522), .B(G116), .C1(new_n518), .C2(new_n519), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n254), .A2(G122), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n400), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n400), .B1(new_n524), .B2(new_n525), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n516), .B(new_n517), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n525), .A2(KEYINPUT14), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n521), .A2(new_n523), .B1(new_n525), .B2(KEYINPUT14), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n530), .B1(new_n531), .B2(KEYINPUT97), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n525), .A2(KEYINPUT14), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n524), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT97), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n400), .B1(new_n532), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT96), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n526), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n524), .A2(KEYINPUT96), .A3(new_n400), .A4(new_n525), .ZN(new_n540));
  INV_X1    g354(.A(new_n514), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n529), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n389), .A2(new_n329), .A3(G953), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n529), .B(new_n544), .C1(new_n537), .C2(new_n542), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(KEYINPUT98), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT98), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n543), .A2(new_n549), .A3(new_n545), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n548), .A2(new_n314), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G478), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(KEYINPUT15), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n553), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n548), .A2(new_n314), .A3(new_n550), .A4(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n554), .A2(KEYINPUT99), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n554), .A2(new_n556), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT99), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n270), .A2(G952), .ZN(new_n561));
  INV_X1    g375(.A(G234), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n561), .B1(new_n562), .B2(new_n269), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  AOI211_X1 g378(.A(new_n314), .B(new_n270), .C1(G234), .C2(G237), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT21), .B(G898), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n512), .A2(new_n557), .A3(new_n560), .A4(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(G210), .B1(G237), .B2(G902), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n252), .A2(KEYINPUT70), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT70), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(G116), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(new_n574), .A3(G119), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n575), .B(KEYINPUT5), .C1(new_n252), .C2(G119), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT5), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n258), .B1(new_n253), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT85), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n255), .A2(new_n261), .A3(new_n262), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n576), .A2(KEYINPUT85), .A3(new_n578), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n581), .A2(new_n582), .A3(new_n427), .A4(new_n583), .ZN(new_n584));
  OAI22_X1  g398(.A1(new_n263), .A2(new_n264), .B1(new_n419), .B2(new_n413), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n584), .B1(new_n418), .B2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(G110), .B(G122), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n584), .B(new_n587), .C1(new_n418), .C2(new_n585), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(KEYINPUT6), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n234), .A2(G125), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n353), .B(new_n216), .C1(new_n217), .C2(new_n220), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT86), .B(G224), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n270), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(KEYINPUT87), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n594), .B(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT6), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n586), .A2(new_n599), .A3(new_n588), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n591), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n596), .A2(KEYINPUT7), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n594), .B(new_n603), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n579), .A2(KEYINPUT88), .A3(new_n582), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT88), .B1(new_n579), .B2(new_n582), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n427), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n581), .A2(new_n582), .A3(new_n409), .A4(new_n583), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n587), .B(KEYINPUT8), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n604), .A2(new_n610), .A3(new_n590), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n314), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n571), .B1(new_n601), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n612), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n591), .A2(new_n598), .A3(new_n600), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n614), .A2(new_n615), .A3(new_n570), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n613), .A2(KEYINPUT89), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(G214), .B1(G237), .B2(G902), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n601), .A2(new_n612), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT89), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n619), .A2(new_n620), .A3(new_n570), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n617), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n569), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n328), .A2(new_n388), .A3(new_n469), .A4(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G101), .ZN(G3));
  OAI21_X1  g439(.A(G472), .B1(new_n293), .B2(G902), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n626), .B1(new_n295), .B2(new_n293), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n469), .A2(new_n388), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n613), .A2(KEYINPUT100), .A3(new_n616), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT100), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n619), .A2(new_n631), .A3(new_n570), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n630), .A2(new_n618), .A3(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT33), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n548), .A2(new_n635), .A3(new_n550), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n546), .A2(KEYINPUT33), .A3(new_n547), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n636), .A2(G478), .A3(new_n314), .A4(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n551), .A2(new_n552), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n511), .A2(new_n640), .A3(new_n568), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n634), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n629), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT34), .B(G104), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G6));
  NAND2_X1  g459(.A1(new_n502), .A2(new_n503), .ZN(new_n646));
  INV_X1    g460(.A(new_n470), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n502), .A2(new_n470), .A3(new_n503), .ZN(new_n649));
  INV_X1    g463(.A(new_n495), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n485), .A2(new_n486), .ZN(new_n651));
  INV_X1    g465(.A(new_n483), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(KEYINPUT93), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n654), .A2(new_n489), .A3(new_n493), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n472), .B1(new_n655), .B2(new_n482), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n314), .B1(new_n650), .B2(new_n656), .ZN(new_n657));
  AOI22_X1  g471(.A1(new_n648), .A2(new_n649), .B1(new_n657), .B2(G475), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n554), .A2(KEYINPUT99), .A3(new_n556), .ZN(new_n659));
  AOI21_X1  g473(.A(KEYINPUT99), .B1(new_n554), .B2(new_n556), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n658), .B(new_n568), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(KEYINPUT101), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n560), .A2(new_n557), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT101), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n663), .A2(new_n664), .A3(new_n568), .A4(new_n658), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n662), .A2(new_n665), .A3(new_n633), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n629), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT35), .B(G107), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G9));
  NOR2_X1   g483(.A1(new_n369), .A2(KEYINPUT36), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n371), .B(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n386), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n382), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n450), .A2(new_n459), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n674), .A2(new_n461), .A3(new_n314), .ZN(new_n675));
  INV_X1    g489(.A(new_n462), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n675), .A2(new_n676), .A3(new_n468), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n673), .A2(new_n677), .A3(new_n390), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n627), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n623), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT37), .B(G110), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G12));
  INV_X1    g496(.A(new_n565), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n563), .B1(new_n683), .B2(G900), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT102), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n663), .A2(new_n658), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n687), .B1(new_n326), .B2(new_n327), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n634), .A2(new_n678), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G128), .ZN(G30));
  XOR2_X1   g505(.A(new_n685), .B(KEYINPUT39), .Z(new_n692));
  NAND2_X1  g506(.A1(new_n469), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT40), .ZN(new_n694));
  OR2_X1    g508(.A1(new_n694), .A2(KEYINPUT104), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(KEYINPUT104), .ZN(new_n696));
  AOI21_X1  g510(.A(KEYINPUT32), .B1(new_n322), .B2(new_n294), .ZN(new_n697));
  AOI211_X1 g511(.A(new_n187), .B(new_n295), .C1(new_n319), .C2(new_n321), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n288), .A2(new_n268), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n274), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n314), .B1(new_n299), .B2(new_n274), .ZN(new_n703));
  OAI21_X1  g517(.A(G472), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n512), .B1(new_n557), .B2(new_n560), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n617), .A2(new_n621), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n618), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n713), .A2(new_n714), .A3(new_n673), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n695), .A2(new_n696), .A3(new_n709), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G143), .ZN(G45));
  NAND3_X1  g531(.A1(new_n511), .A2(new_n640), .A3(new_n686), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n634), .A2(new_n678), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n328), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(KEYINPUT105), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT105), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n328), .A2(new_n722), .A3(new_n719), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G146), .ZN(G48));
  INV_X1    g539(.A(new_n388), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n461), .B1(new_n674), .B2(new_n314), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n727), .A2(new_n460), .A3(new_n391), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT75), .B1(new_n699), .B2(new_n318), .ZN(new_n731));
  INV_X1    g545(.A(new_n327), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n642), .B(new_n730), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT106), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n328), .A2(KEYINPUT106), .A3(new_n642), .A4(new_n730), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XOR2_X1   g551(.A(KEYINPUT41), .B(G113), .Z(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT107), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n737), .B(new_n739), .ZN(G15));
  NAND3_X1  g554(.A1(new_n666), .A2(new_n328), .A3(new_n730), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G116), .ZN(G18));
  NAND4_X1  g556(.A1(new_n728), .A2(new_n618), .A3(new_n632), .A4(new_n630), .ZN(new_n743));
  INV_X1    g557(.A(new_n673), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n743), .A2(new_n569), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n328), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G119), .ZN(G21));
  NOR4_X1   g561(.A1(new_n727), .A2(new_n460), .A3(new_n391), .A4(new_n567), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n633), .A2(new_n663), .A3(new_n748), .A4(new_n511), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n300), .A2(new_n304), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n276), .B1(new_n750), .B2(new_n274), .ZN(new_n751));
  INV_X1    g565(.A(new_n319), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n294), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n626), .A2(new_n388), .A3(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  XOR2_X1   g569(.A(new_n755), .B(G122), .Z(G24));
  AND3_X1   g570(.A1(new_n511), .A2(new_n640), .A3(new_n686), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n757), .A2(new_n626), .A3(new_n673), .A4(new_n753), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n743), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(new_n353), .ZN(G27));
  OR2_X1    g574(.A1(new_n323), .A2(KEYINPUT109), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n323), .A2(KEYINPUT109), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n761), .A2(new_n296), .A3(new_n318), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n465), .A2(new_n467), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT108), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n465), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n765), .A2(G469), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n391), .B1(new_n768), .B2(new_n463), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n714), .B1(new_n617), .B2(new_n621), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(new_n770), .A3(new_n388), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n763), .A2(new_n772), .A3(KEYINPUT42), .A4(new_n757), .ZN(new_n773));
  AOI211_X1 g587(.A(new_n718), .B(new_n771), .C1(new_n326), .C2(new_n327), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n773), .B1(new_n774), .B2(KEYINPUT42), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G131), .ZN(G33));
  AOI211_X1 g590(.A(new_n687), .B(new_n771), .C1(new_n326), .C2(new_n327), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(new_n200), .ZN(G36));
  AND3_X1   g592(.A1(new_n765), .A2(KEYINPUT45), .A3(new_n767), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n780));
  AOI211_X1 g594(.A(new_n461), .B(new_n779), .C1(new_n780), .C2(new_n764), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(new_n462), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n782), .A2(KEYINPUT46), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n675), .B1(new_n782), .B2(KEYINPUT46), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n390), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n692), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n770), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n512), .A2(new_n640), .ZN(new_n789));
  XOR2_X1   g603(.A(new_n789), .B(KEYINPUT43), .Z(new_n790));
  AND3_X1   g604(.A1(new_n790), .A2(new_n627), .A3(new_n673), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n788), .B1(new_n791), .B2(KEYINPUT44), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n787), .B(new_n792), .C1(KEYINPUT44), .C2(new_n791), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G137), .ZN(G39));
  XNOR2_X1  g608(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n785), .B(new_n795), .ZN(new_n796));
  NOR4_X1   g610(.A1(new_n328), .A2(new_n388), .A3(new_n718), .A4(new_n788), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT111), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G140), .ZN(G42));
  NOR2_X1   g614(.A1(new_n727), .A2(new_n460), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n802), .A2(KEYINPUT49), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n388), .A2(new_n390), .A3(new_n618), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n802), .A2(KEYINPUT49), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n803), .A2(new_n804), .A3(new_n805), .A4(new_n789), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n706), .A3(new_n713), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n754), .A2(new_n563), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n790), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n770), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n801), .A2(new_n391), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n810), .B1(new_n796), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n712), .A2(new_n618), .A3(new_n729), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n809), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT50), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n809), .A2(KEYINPUT50), .A3(new_n814), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n770), .A2(new_n728), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n820), .A2(KEYINPUT121), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(KEYINPUT121), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n821), .A2(new_n822), .A3(new_n563), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(new_n388), .A3(new_n706), .ZN(new_n824));
  OR3_X1    g638(.A1(new_n824), .A2(new_n511), .A3(new_n640), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n626), .A2(new_n753), .A3(new_n673), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n823), .A2(new_n790), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n819), .B(new_n825), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  OR3_X1    g642(.A1(new_n812), .A2(new_n813), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n813), .B1(new_n812), .B2(new_n828), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n763), .A2(new_n388), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT48), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n809), .A2(new_n633), .A3(new_n728), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n511), .A2(new_n640), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n834), .B(new_n561), .C1(new_n835), .C2(new_n824), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n829), .A2(new_n830), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT122), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n759), .B1(new_n688), .B2(new_n689), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n673), .A2(new_n685), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n769), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n769), .A2(KEYINPUT115), .A3(new_n842), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n709), .A2(new_n847), .A3(new_n633), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n328), .A2(new_n722), .A3(new_n719), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n722), .B1(new_n328), .B2(new_n719), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n841), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT52), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n724), .A2(KEYINPUT52), .A3(new_n841), .A4(new_n848), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n755), .B1(new_n328), .B2(new_n745), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n856), .A2(new_n741), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(new_n737), .A3(new_n775), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n512), .A2(new_n558), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n860), .A2(new_n622), .A3(new_n567), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n629), .A2(new_n861), .B1(new_n679), .B2(new_n623), .ZN(new_n862));
  OR3_X1    g676(.A1(new_n641), .A2(new_n622), .A3(KEYINPUT112), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT112), .B1(new_n641), .B2(new_n622), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n629), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n624), .A2(new_n862), .A3(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n673), .A2(new_n390), .A3(new_n677), .ZN(new_n867));
  INV_X1    g681(.A(new_n558), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT113), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n658), .A2(new_n868), .A3(new_n869), .A4(new_n686), .ZN(new_n870));
  AOI211_X1 g684(.A(new_n647), .B(new_n505), .C1(new_n495), .C2(new_n501), .ZN(new_n871));
  OAI22_X1  g685(.A1(new_n504), .A2(new_n871), .B1(new_n509), .B2(new_n510), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n554), .A2(new_n556), .A3(new_n686), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT113), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AND4_X1   g688(.A1(new_n867), .A2(new_n870), .A3(new_n770), .A4(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n875), .B1(new_n731), .B2(new_n732), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n769), .A2(new_n770), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n758), .A2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT114), .B1(new_n880), .B2(new_n777), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n878), .B1(new_n328), .B2(new_n875), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT114), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n688), .A2(new_n772), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n866), .B1(new_n881), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g700(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n855), .A2(new_n859), .A3(new_n886), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT117), .ZN(new_n890));
  INV_X1    g704(.A(new_n866), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n880), .A2(KEYINPUT114), .A3(new_n777), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n883), .B1(new_n882), .B2(new_n884), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n894), .A2(new_n858), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT117), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n895), .A2(new_n896), .A3(new_n855), .A4(new_n888), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n855), .A2(new_n859), .A3(new_n886), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT53), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n890), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT54), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(KEYINPUT118), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n888), .B1(new_n895), .B2(new_n855), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n858), .A2(KEYINPUT119), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT119), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n857), .A2(new_n737), .A3(new_n775), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  OAI211_X1 g723(.A(KEYINPUT53), .B(new_n891), .C1(new_n892), .C2(new_n893), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n910), .B1(new_n853), .B2(new_n854), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n909), .A2(new_n911), .A3(KEYINPUT120), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT120), .ZN(new_n913));
  AOI211_X1 g727(.A(new_n899), .B(new_n866), .C1(new_n881), .C2(new_n885), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n855), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n913), .B1(new_n915), .B2(new_n908), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n904), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT54), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT118), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n901), .A2(new_n920), .A3(KEYINPUT54), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n903), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n838), .A2(new_n839), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n840), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(G952), .A2(G953), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n807), .B1(new_n924), .B2(new_n925), .ZN(G75));
  NOR2_X1   g740(.A1(new_n270), .A2(G952), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n917), .A2(new_n314), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT56), .B1(new_n929), .B2(G210), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n591), .A2(new_n600), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT123), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT55), .Z(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(new_n598), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n928), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(new_n930), .B2(new_n934), .ZN(G51));
  INV_X1    g750(.A(new_n904), .ZN(new_n937));
  AOI21_X1  g751(.A(KEYINPUT120), .B1(new_n909), .B2(new_n911), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n915), .A2(new_n908), .A3(new_n913), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(KEYINPUT54), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n919), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n462), .B(KEYINPUT57), .Z(new_n944));
  OAI21_X1  g758(.A(new_n674), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n929), .A2(new_n781), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n927), .B1(new_n945), .B2(new_n946), .ZN(G54));
  AND2_X1   g761(.A1(KEYINPUT58), .A2(G475), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n929), .A2(new_n502), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n502), .B1(new_n929), .B2(new_n948), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n949), .A2(new_n950), .A3(new_n927), .ZN(G60));
  INV_X1    g765(.A(KEYINPUT124), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n636), .A2(new_n637), .ZN(new_n953));
  NAND2_X1  g767(.A1(G478), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT59), .Z(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n953), .B1(new_n922), .B2(new_n956), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n953), .A2(new_n956), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n917), .A2(new_n918), .ZN(new_n959));
  AOI211_X1 g773(.A(KEYINPUT54), .B(new_n904), .C1(new_n912), .C2(new_n916), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n928), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n952), .B1(new_n957), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n927), .B1(new_n942), .B2(new_n958), .ZN(new_n964));
  AOI22_X1  g778(.A1(KEYINPUT117), .A2(new_n889), .B1(new_n898), .B2(new_n899), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n918), .B1(new_n965), .B2(new_n897), .ZN(new_n966));
  AOI22_X1  g780(.A1(new_n966), .A2(new_n920), .B1(new_n917), .B2(new_n918), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n955), .B1(new_n967), .B2(new_n903), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n964), .B(KEYINPUT124), .C1(new_n968), .C2(new_n953), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n963), .A2(new_n969), .ZN(G63));
  NAND2_X1  g784(.A1(G217), .A2(G902), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT60), .Z(new_n972));
  NAND3_X1  g786(.A1(new_n940), .A2(new_n671), .A3(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n940), .A2(new_n972), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n928), .B(new_n973), .C1(new_n974), .C2(new_n376), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT61), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(G66));
  INV_X1    g791(.A(new_n566), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n270), .B1(new_n978), .B2(new_n595), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n891), .A2(new_n857), .A3(new_n737), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n979), .B1(new_n980), .B2(new_n270), .ZN(new_n981));
  INV_X1    g795(.A(G898), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n932), .B1(new_n982), .B2(G953), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n981), .B(new_n983), .ZN(G69));
  NAND2_X1  g798(.A1(new_n240), .A2(new_n251), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n497), .B(KEYINPUT125), .Z(new_n986));
  XNOR2_X1  g800(.A(new_n985), .B(new_n986), .ZN(new_n987));
  OAI211_X1 g801(.A(G900), .B(G953), .C1(new_n987), .C2(G227), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n988), .B1(G227), .B2(new_n987), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n724), .A2(new_n841), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n793), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT127), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n831), .A2(new_n634), .A3(new_n708), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n777), .B1(new_n787), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n799), .A2(new_n775), .A3(new_n994), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(G953), .B1(new_n996), .B2(new_n987), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n990), .A2(new_n716), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n998), .A2(KEYINPUT62), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT126), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n998), .A2(KEYINPUT62), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n860), .A2(new_n835), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n693), .A2(new_n788), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n328), .A2(new_n388), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n799), .A2(new_n1001), .A3(new_n793), .A4(new_n1004), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1000), .A2(new_n1005), .ZN(new_n1006));
  OR2_X1    g820(.A1(new_n1006), .A2(new_n987), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n989), .B1(new_n997), .B2(new_n1007), .ZN(G72));
  AOI22_X1  g822(.A1(new_n996), .A2(new_n312), .B1(new_n1006), .B2(new_n702), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1009), .A2(new_n980), .ZN(new_n1010));
  NAND2_X1  g824(.A1(G472), .A2(G902), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT63), .Z(new_n1012));
  NOR2_X1   g826(.A1(new_n702), .A2(new_n312), .ZN(new_n1013));
  AND3_X1   g827(.A1(new_n901), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n928), .B1(new_n1013), .B2(new_n1012), .ZN(new_n1015));
  NOR3_X1   g829(.A1(new_n1010), .A2(new_n1014), .A3(new_n1015), .ZN(G57));
endmodule


