//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n549,
    new_n551, new_n552, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT65), .Z(G319));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n459), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n459), .A2(new_n461), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n462), .A2(new_n468), .ZN(G160));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G136), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n472), .A2(new_n461), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  MUX2_X1   g051(.A(G100), .B(G112), .S(G2105), .Z(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2104), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n474), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  NAND2_X1  g055(.A1(new_n461), .A2(G102), .ZN(new_n481));
  NAND2_X1  g056(.A1(G114), .A2(G2105), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n463), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AND2_X1   g058(.A1(G126), .A2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n484), .B1(new_n470), .B2(new_n471), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT66), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT66), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(new_n484), .C1(new_n470), .C2(new_n471), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n483), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  OAI211_X1 g064(.A(G138), .B(new_n461), .C1(new_n470), .C2(new_n471), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n459), .A2(new_n492), .A3(G138), .A4(new_n461), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  INV_X1    g071(.A(KEYINPUT67), .ZN(new_n497));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(KEYINPUT5), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(KEYINPUT67), .A3(G543), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n499), .A2(new_n501), .B1(KEYINPUT5), .B2(new_n498), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n502), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(new_n504), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n505), .A2(new_n512), .ZN(G166));
  NAND3_X1  g088(.A1(new_n502), .A2(G63), .A3(G651), .ZN(new_n514));
  XOR2_X1   g089(.A(new_n514), .B(KEYINPUT68), .Z(new_n515));
  NAND2_X1  g090(.A1(new_n499), .A2(new_n501), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n498), .A2(KEYINPUT5), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n516), .A2(new_n517), .A3(new_n510), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G89), .ZN(new_n520));
  XOR2_X1   g095(.A(KEYINPUT71), .B(KEYINPUT7), .Z(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n521), .B(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT69), .ZN(new_n524));
  INV_X1    g099(.A(new_n509), .ZN(new_n525));
  NOR2_X1   g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n508), .A2(KEYINPUT69), .A3(new_n509), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n498), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  XOR2_X1   g105(.A(KEYINPUT70), .B(G51), .Z(new_n531));
  OAI211_X1 g106(.A(new_n520), .B(new_n523), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n515), .A2(new_n532), .ZN(G168));
  NAND2_X1  g108(.A1(new_n529), .A2(G52), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n535), .B2(new_n518), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n502), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n504), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n536), .A2(new_n538), .ZN(G171));
  AOI22_X1  g114(.A1(new_n502), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT72), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g117(.A(G651), .B1(new_n540), .B2(new_n541), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n519), .A2(G81), .B1(new_n529), .B2(G43), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(G188));
  NAND2_X1  g128(.A1(new_n529), .A2(G53), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT9), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n518), .A2(KEYINPUT73), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT73), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n502), .A2(new_n557), .A3(new_n510), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n556), .A2(G91), .A3(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n502), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n560), .A2(new_n504), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n555), .A2(new_n559), .A3(new_n561), .ZN(G299));
  INV_X1    g137(.A(G171), .ZN(G301));
  INV_X1    g138(.A(G168), .ZN(G286));
  INV_X1    g139(.A(G166), .ZN(G303));
  NAND2_X1  g140(.A1(new_n516), .A2(new_n517), .ZN(new_n566));
  INV_X1    g141(.A(G74), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n568), .A2(G651), .B1(new_n529), .B2(G49), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n556), .A2(G87), .A3(new_n558), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(G288));
  NAND3_X1  g146(.A1(new_n510), .A2(G48), .A3(G543), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(G73), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G61), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n566), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n573), .B1(new_n576), .B2(G651), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n556), .A2(G86), .A3(new_n558), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT74), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n579), .A2(new_n580), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n582), .A2(new_n583), .ZN(G305));
  AOI22_X1  g159(.A1(new_n519), .A2(G85), .B1(new_n529), .B2(G47), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n504), .B2(new_n586), .ZN(G290));
  INV_X1    g162(.A(G868), .ZN(new_n588));
  NOR2_X1   g163(.A1(G301), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n556), .A2(G92), .A3(new_n558), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n566), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(new_n529), .B2(G54), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n589), .B1(new_n597), .B2(new_n588), .ZN(G284));
  AOI21_X1  g173(.A(new_n589), .B1(new_n597), .B2(new_n588), .ZN(G321));
  MUX2_X1   g174(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g175(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g176(.A(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n597), .B1(new_n602), .B2(G860), .ZN(G148));
  NAND2_X1  g178(.A1(new_n592), .A2(new_n596), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(G559), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G868), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G868), .B2(new_n546), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT75), .ZN(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g184(.A1(new_n473), .A2(G2104), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT12), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(KEYINPUT13), .Z(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G2100), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT76), .Z(new_n614));
  NOR2_X1   g189(.A1(new_n612), .A2(G2100), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT77), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n473), .A2(G135), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n475), .A2(G123), .ZN(new_n618));
  AND2_X1   g193(.A1(G111), .A2(G2105), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(G99), .B2(new_n461), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n617), .B(new_n618), .C1(new_n463), .C2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(G2096), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n614), .A2(new_n616), .A3(new_n623), .ZN(G156));
  INV_X1    g199(.A(KEYINPUT14), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT15), .B(G2435), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2438), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2427), .ZN(new_n628));
  INV_X1    g203(.A(G2430), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n625), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(new_n629), .B2(new_n628), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G1341), .B(G1348), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n631), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n631), .A2(new_n637), .ZN(new_n639));
  AND3_X1   g214(.A1(new_n638), .A2(G14), .A3(new_n639), .ZN(G401));
  XOR2_X1   g215(.A(G2072), .B(G2078), .Z(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  XNOR2_X1  g218(.A(G2067), .B(G2678), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT78), .B(KEYINPUT18), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n642), .A2(KEYINPUT17), .A3(new_n643), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n643), .B1(new_n642), .B2(KEYINPUT17), .ZN(new_n649));
  INV_X1    g224(.A(new_n644), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n643), .A2(new_n644), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n642), .B1(new_n652), .B2(KEYINPUT17), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n647), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(new_n622), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2100), .ZN(G227));
  XNOR2_X1  g231(.A(G1956), .B(G2474), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT80), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1961), .B(G1966), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G1971), .B(G1976), .Z(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT79), .B(KEYINPUT19), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT20), .Z(new_n666));
  OR2_X1    g241(.A1(new_n658), .A2(new_n660), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n667), .A2(new_n661), .A3(new_n664), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n666), .B(new_n668), .C1(new_n664), .C2(new_n667), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1991), .B(G1996), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1981), .B(G1986), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n671), .B(new_n674), .ZN(G229));
  OR2_X1    g250(.A1(G6), .A2(G16), .ZN(new_n676));
  INV_X1    g251(.A(G16), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n676), .B1(G305), .B2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT83), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n679), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT32), .B(G1981), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(G16), .A2(G22), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(G166), .B2(G16), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT85), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT84), .B(G1971), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n677), .A2(G23), .ZN(new_n691));
  INV_X1    g266(.A(G288), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(new_n677), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT33), .B(G1976), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n685), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT82), .B(KEYINPUT34), .Z(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n685), .A2(new_n696), .A3(new_n698), .ZN(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(KEYINPUT81), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(KEYINPUT81), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n705), .A2(G25), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n473), .A2(G131), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n475), .A2(G119), .ZN(new_n708));
  MUX2_X1   g283(.A(G95), .B(G107), .S(G2105), .Z(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G2104), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n707), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n706), .B1(new_n712), .B2(new_n705), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT35), .B(G1991), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(KEYINPUT86), .A2(KEYINPUT36), .ZN(new_n716));
  INV_X1    g291(.A(G1986), .ZN(new_n717));
  OR2_X1    g292(.A1(G16), .A2(G24), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G290), .B2(new_n677), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n715), .B(new_n716), .C1(new_n717), .C2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n717), .B2(new_n719), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n700), .A2(new_n701), .A3(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(KEYINPUT86), .A2(KEYINPUT36), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(KEYINPUT95), .B1(G29), .B2(G32), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT93), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G129), .B2(new_n475), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n473), .A2(G141), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT94), .B(KEYINPUT26), .ZN(new_n730));
  NAND3_X1  g305(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n728), .A2(new_n729), .A3(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(new_n702), .ZN(new_n734));
  MUX2_X1   g309(.A(new_n725), .B(KEYINPUT95), .S(new_n734), .Z(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT27), .B(G1996), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(G29), .A2(G33), .ZN(new_n738));
  AOI21_X1  g313(.A(KEYINPUT25), .B1(new_n464), .B2(G103), .ZN(new_n739));
  AND3_X1   g314(.A1(new_n464), .A2(KEYINPUT25), .A3(G103), .ZN(new_n740));
  INV_X1    g315(.A(G139), .ZN(new_n741));
  OAI22_X1  g316(.A1(new_n739), .A2(new_n740), .B1(new_n466), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n459), .A2(G127), .ZN(new_n743));
  NAND2_X1  g318(.A1(G115), .A2(G2104), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n461), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n738), .B1(new_n746), .B2(G29), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT92), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G2072), .ZN(new_n749));
  NOR2_X1   g324(.A1(G168), .A2(new_n677), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n677), .B2(G21), .ZN(new_n751));
  INV_X1    g326(.A(G1966), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n705), .A2(G27), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G164), .B2(new_n705), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G2078), .ZN(new_n756));
  NOR4_X1   g331(.A1(new_n737), .A2(new_n749), .A3(new_n753), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n751), .A2(new_n752), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT96), .ZN(new_n759));
  INV_X1    g334(.A(new_n705), .ZN(new_n760));
  NOR2_X1   g335(.A1(KEYINPUT24), .A2(G34), .ZN(new_n761));
  AND2_X1   g336(.A1(KEYINPUT24), .A2(G34), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G160), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(new_n702), .ZN(new_n765));
  INV_X1    g340(.A(G2084), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n621), .A2(new_n760), .ZN(new_n769));
  OR2_X1    g344(.A1(KEYINPUT30), .A2(G28), .ZN(new_n770));
  NAND2_X1  g345(.A1(KEYINPUT30), .A2(G28), .ZN(new_n771));
  AOI21_X1  g346(.A(G29), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT31), .B(G11), .Z(new_n773));
  NOR3_X1   g348(.A1(new_n769), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n767), .A2(new_n768), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n677), .A2(G5), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G171), .B2(new_n677), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n777), .A2(G1961), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(G1961), .ZN(new_n779));
  NOR3_X1   g354(.A1(new_n775), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  AND3_X1   g355(.A1(new_n757), .A2(new_n759), .A3(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT97), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n677), .A2(G20), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT23), .Z(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G299), .B2(G16), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1956), .ZN(new_n788));
  NOR2_X1   g363(.A1(G4), .A2(G16), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT87), .Z(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n604), .B2(new_n677), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT88), .B(G1348), .Z(new_n792));
  OAI21_X1  g367(.A(new_n788), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n791), .B2(new_n792), .ZN(new_n794));
  NOR2_X1   g369(.A1(G16), .A2(G19), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n547), .B2(G16), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(G1341), .Z(new_n797));
  NAND2_X1  g372(.A1(new_n760), .A2(G26), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT28), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n473), .A2(G140), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT89), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n475), .A2(G128), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT90), .ZN(new_n803));
  MUX2_X1   g378(.A(G104), .B(G116), .S(G2105), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(G2104), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT91), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n801), .A2(new_n803), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n799), .B1(new_n807), .B2(G29), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G2067), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n705), .A2(G35), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G162), .B2(new_n705), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT29), .ZN(new_n812));
  INV_X1    g387(.A(G2090), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n794), .A2(new_n797), .A3(new_n809), .A4(new_n814), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n783), .A2(new_n784), .A3(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n723), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n700), .A2(new_n701), .A3(new_n721), .A4(new_n817), .ZN(new_n818));
  AND3_X1   g393(.A1(new_n724), .A2(new_n816), .A3(new_n818), .ZN(G311));
  NAND3_X1  g394(.A1(new_n724), .A2(new_n816), .A3(new_n818), .ZN(G150));
  AOI22_X1  g395(.A1(new_n502), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(KEYINPUT98), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(KEYINPUT98), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n822), .A2(G651), .A3(new_n823), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n519), .A2(G93), .B1(new_n529), .B2(G55), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(G860), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT37), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n546), .A2(new_n826), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n544), .A2(new_n824), .A3(new_n545), .A4(new_n825), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT38), .Z(new_n832));
  NOR2_X1   g407(.A1(new_n604), .A2(new_n602), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n835), .A2(KEYINPUT39), .ZN(new_n836));
  INV_X1    g411(.A(G860), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n835), .B2(KEYINPUT39), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n828), .B1(new_n836), .B2(new_n838), .ZN(G145));
  XNOR2_X1  g414(.A(new_n611), .B(new_n711), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n473), .A2(G142), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT100), .Z(new_n842));
  NAND2_X1  g417(.A1(new_n475), .A2(G130), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT101), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n844), .A2(new_n461), .A3(G118), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n844), .B1(new_n461), .B2(G118), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n846), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n842), .B(new_n843), .C1(new_n845), .C2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n840), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT102), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n807), .B(new_n495), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n733), .B(new_n746), .Z(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(G160), .B(KEYINPUT99), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n621), .B(new_n479), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n857), .B1(new_n853), .B2(new_n849), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(KEYINPUT103), .B(G37), .Z(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n850), .B(new_n853), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n861), .B1(new_n857), .B2(new_n862), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT40), .Z(G395));
  NAND3_X1  g439(.A1(new_n824), .A2(new_n588), .A3(new_n825), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n831), .B(new_n605), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n597), .A2(G299), .ZN(new_n868));
  NAND3_X1  g443(.A1(G299), .A2(new_n592), .A3(new_n596), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(KEYINPUT104), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT104), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n597), .A2(new_n871), .A3(G299), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n868), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT41), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n870), .ZN(new_n876));
  INV_X1    g451(.A(new_n868), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n876), .A2(new_n874), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n867), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n876), .A2(new_n877), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n867), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n882), .A2(KEYINPUT42), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(KEYINPUT42), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(G303), .B1(new_n582), .B2(new_n583), .ZN(new_n886));
  INV_X1    g461(.A(new_n583), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n887), .A2(G166), .A3(new_n581), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n692), .B(G290), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n890), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n892), .A2(new_n886), .A3(new_n888), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n894), .A2(KEYINPUT105), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n885), .A2(new_n895), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n883), .B(new_n884), .C1(KEYINPUT105), .C2(new_n894), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n866), .B1(new_n898), .B2(G868), .ZN(G295));
  AOI21_X1  g474(.A(new_n866), .B1(new_n898), .B2(G868), .ZN(G331));
  NAND2_X1  g475(.A1(G286), .A2(G301), .ZN(new_n901));
  NAND2_X1  g476(.A1(G168), .A2(G171), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n903), .A2(new_n831), .ZN(new_n904));
  AOI22_X1  g479(.A1(new_n901), .A2(new_n902), .B1(new_n829), .B2(new_n830), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n880), .A2(KEYINPUT41), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n873), .A2(new_n874), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(new_n873), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n894), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n904), .A2(new_n905), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n875), .B2(new_n878), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT106), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n892), .A2(new_n886), .A3(new_n888), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n892), .B1(new_n886), .B2(new_n888), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n891), .A2(KEYINPUT106), .A3(new_n893), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n914), .A2(new_n910), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n912), .A2(new_n921), .A3(new_n860), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT43), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n925));
  INV_X1    g500(.A(G37), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n912), .A2(new_n921), .A3(KEYINPUT43), .A4(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n912), .A2(new_n921), .A3(new_n923), .A4(new_n926), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n929), .A2(KEYINPUT44), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT107), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AND4_X1   g507(.A1(KEYINPUT107), .A2(new_n931), .A3(KEYINPUT44), .A4(new_n929), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n928), .B1(new_n932), .B2(new_n933), .ZN(G397));
  INV_X1    g509(.A(G1384), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n495), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT45), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(G160), .A2(G40), .ZN(new_n939));
  OR3_X1    g514(.A1(new_n938), .A2(KEYINPUT108), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT108), .B1(new_n938), .B2(new_n939), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n807), .B(G2067), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT109), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n942), .A2(KEYINPUT109), .A3(new_n943), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n733), .B(G1996), .ZN(new_n946));
  AOI211_X1 g521(.A(new_n944), .B(new_n945), .C1(new_n942), .C2(new_n946), .ZN(new_n947));
  XOR2_X1   g522(.A(new_n711), .B(new_n714), .Z(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT110), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n942), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n942), .ZN(new_n952));
  OR2_X1    g527(.A1(G290), .A2(G1986), .ZN(new_n953));
  NAND2_X1  g528(.A1(G290), .A2(G1986), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n936), .A2(KEYINPUT111), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT50), .ZN(new_n958));
  AOI21_X1  g533(.A(G1384), .B1(new_n489), .B2(new_n494), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n957), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n960), .B1(new_n495), .B2(new_n935), .ZN(new_n965));
  AOI211_X1 g540(.A(KEYINPUT111), .B(G1384), .C1(new_n489), .C2(new_n494), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n967), .A2(KEYINPUT112), .A3(new_n958), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n964), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n959), .A2(new_n970), .A3(new_n958), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n970), .B1(new_n959), .B2(new_n958), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n939), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n969), .A2(new_n813), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n959), .A2(KEYINPUT45), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n938), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n939), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G1971), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n975), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(G303), .A2(G8), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT55), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n982), .A2(G8), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n957), .A2(new_n978), .A3(new_n961), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(G8), .ZN(new_n988));
  INV_X1    g563(.A(G1981), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n577), .A2(new_n989), .A3(new_n578), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n502), .A2(G86), .A3(new_n510), .ZN(new_n991));
  AOI22_X1  g566(.A1(new_n502), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n572), .B(new_n991), .C1(new_n992), .C2(new_n504), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(G1981), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT49), .B1(new_n990), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n988), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n990), .A2(KEYINPUT49), .A3(new_n994), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT115), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT115), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n990), .A2(new_n994), .A3(new_n999), .A4(KEYINPUT49), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n692), .A2(G1976), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n987), .A2(new_n1002), .A3(G8), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n996), .A2(new_n1001), .B1(new_n1003), .B2(KEYINPUT52), .ZN(new_n1004));
  INV_X1    g579(.A(G1976), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT52), .B1(G288), .B2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n987), .A2(new_n1002), .A3(new_n1006), .A4(G8), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT114), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G8), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1010), .B1(new_n967), .B2(new_n978), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1011), .A2(KEYINPUT114), .A3(new_n1002), .A4(new_n1006), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1004), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n986), .A2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n988), .B(KEYINPUT116), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n998), .A2(new_n1000), .ZN(new_n1017));
  INV_X1    g592(.A(new_n995), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1011), .A2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1005), .B(new_n692), .C1(new_n1017), .C2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1016), .B1(new_n1020), .B2(new_n990), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1015), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT120), .ZN(new_n1023));
  AOI21_X1  g598(.A(G1348), .B1(new_n969), .B2(new_n974), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n987), .A2(G2067), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1023), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1025), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT113), .B1(new_n936), .B2(KEYINPUT50), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n978), .B1(new_n1028), .B2(new_n971), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1029), .B1(new_n964), .B2(new_n968), .ZN(new_n1030));
  OAI211_X1 g605(.A(KEYINPUT120), .B(new_n1027), .C1(new_n1030), .C2(G1348), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1026), .A2(new_n597), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G1956), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n959), .A2(KEYINPUT50), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1034), .B1(new_n967), .B2(KEYINPUT50), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1033), .B1(new_n1035), .B2(new_n939), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT56), .B(G2072), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n977), .A2(new_n978), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n1040));
  NAND2_X1  g615(.A1(G299), .A2(new_n1040), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n555), .A2(KEYINPUT57), .A3(new_n559), .A4(new_n561), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1039), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1036), .A2(new_n1038), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT119), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT119), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1036), .A2(new_n1047), .A3(new_n1038), .A4(new_n1044), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1032), .A2(new_n1043), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT60), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1026), .A2(new_n1050), .A3(new_n1031), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1026), .A2(new_n1031), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n604), .B1(new_n1052), .B2(KEYINPUT60), .ZN(new_n1053));
  AOI211_X1 g628(.A(new_n1050), .B(new_n597), .C1(new_n1026), .C2(new_n1031), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1051), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1043), .A2(KEYINPUT61), .A3(new_n1045), .ZN(new_n1056));
  XOR2_X1   g631(.A(KEYINPUT58), .B(G1341), .Z(new_n1057));
  NAND2_X1  g632(.A1(new_n987), .A2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(new_n979), .B2(G1996), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT59), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT121), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1059), .A2(new_n547), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1061), .B1(new_n1059), .B2(new_n547), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1060), .A2(KEYINPUT121), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1056), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT61), .B1(new_n1067), .B2(new_n1043), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1049), .B1(new_n1055), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT112), .B1(new_n967), .B2(new_n958), .ZN(new_n1071));
  NOR4_X1   g646(.A1(new_n965), .A2(new_n966), .A3(new_n963), .A4(KEYINPUT50), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n974), .B(new_n766), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n939), .B1(KEYINPUT45), .B2(new_n959), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1074), .B1(new_n967), .B2(KEYINPUT45), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n752), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1010), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(G286), .A2(G8), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT122), .ZN(new_n1079));
  XNOR2_X1  g654(.A(new_n1078), .B(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT123), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT51), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g658(.A(KEYINPUT123), .B(KEYINPUT51), .C1(new_n1077), .C2(new_n1080), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1030), .A2(new_n766), .B1(new_n752), .B2(new_n1075), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1078), .B(KEYINPUT122), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n1090));
  AND2_X1   g665(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1003), .A2(KEYINPUT52), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1092), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1090), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1035), .A2(new_n939), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1095), .A2(new_n813), .B1(new_n980), .B2(new_n979), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n984), .B1(new_n1096), .B2(new_n1010), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1004), .A2(KEYINPUT117), .A3(new_n1013), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1094), .A2(new_n986), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n1030), .A2(G1961), .ZN(new_n1101));
  XOR2_X1   g676(.A(KEYINPUT124), .B(KEYINPUT53), .Z(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n979), .B2(G2078), .ZN(new_n1103));
  INV_X1    g678(.A(G2078), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT53), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1101), .B(new_n1103), .C1(new_n1075), .C2(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(G171), .B(KEYINPUT54), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n462), .ZN(new_n1109));
  XOR2_X1   g684(.A(new_n468), .B(KEYINPUT125), .Z(new_n1110));
  INV_X1    g685(.A(KEYINPUT126), .ZN(new_n1111));
  OAI211_X1 g686(.A(KEYINPUT53), .B(G40), .C1(new_n1111), .C2(G2078), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(new_n1111), .B2(G2078), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n977), .A2(new_n1109), .A3(new_n1110), .A4(new_n1113), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1103), .A2(new_n1114), .A3(new_n1107), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1106), .A2(new_n1108), .B1(new_n1101), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1089), .A2(new_n1100), .A3(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1022), .B1(new_n1070), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT118), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n986), .A2(new_n1097), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1077), .A2(G168), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1120), .A2(new_n1094), .A3(new_n1098), .A4(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT63), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1119), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1119), .B(new_n1124), .C1(new_n1099), .C2(new_n1121), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n982), .A2(G8), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1121), .B1(new_n984), .B2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1014), .A2(new_n1124), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(new_n986), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1126), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1087), .B1(new_n1086), .B2(new_n1010), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT51), .B1(new_n1133), .B2(KEYINPUT123), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1084), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1132), .B(new_n1088), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1106), .A2(G171), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1099), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1132), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1140));
  OAI22_X1  g715(.A1(new_n1125), .A2(new_n1131), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n956), .B1(new_n1118), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n947), .A2(new_n712), .A3(new_n714), .ZN(new_n1143));
  OR2_X1    g718(.A1(new_n807), .A2(G2067), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n952), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(G1996), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n942), .A2(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(KEYINPUT46), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n942), .B1(new_n943), .B2(new_n733), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  XOR2_X1   g725(.A(new_n1150), .B(KEYINPUT47), .Z(new_n1151));
  INV_X1    g726(.A(new_n951), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n952), .A2(new_n953), .ZN(new_n1153));
  XNOR2_X1  g728(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  AOI211_X1 g730(.A(new_n1145), .B(new_n1151), .C1(new_n1152), .C2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1142), .A2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g732(.A1(G401), .A2(G227), .A3(new_n457), .ZN(new_n1159));
  NOR3_X1   g733(.A1(new_n863), .A2(G229), .A3(new_n1159), .ZN(new_n1160));
  AND3_X1   g734(.A1(new_n1160), .A2(new_n924), .A3(new_n927), .ZN(G308));
  NAND3_X1  g735(.A1(new_n1160), .A2(new_n924), .A3(new_n927), .ZN(G225));
endmodule


