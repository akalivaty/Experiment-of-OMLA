

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593;

  XOR2_X2 U324 ( .A(n368), .B(n367), .Z(n419) );
  XNOR2_X1 U325 ( .A(n455), .B(n379), .ZN(n380) );
  XNOR2_X1 U326 ( .A(n392), .B(KEYINPUT109), .ZN(n393) );
  XNOR2_X1 U327 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U328 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U329 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U330 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U331 ( .A(n450), .B(KEYINPUT121), .ZN(n451) );
  XNOR2_X1 U332 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U333 ( .A(n490), .B(KEYINPUT37), .ZN(n491) );
  XNOR2_X1 U334 ( .A(n342), .B(n341), .ZN(n348) );
  XNOR2_X1 U335 ( .A(n492), .B(n491), .ZN(n514) );
  XNOR2_X1 U336 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U337 ( .A(n409), .B(n408), .Z(n583) );
  XNOR2_X1 U338 ( .A(G183GAT), .B(KEYINPUT124), .ZN(n473) );
  XNOR2_X1 U339 ( .A(n495), .B(G106GAT), .ZN(n496) );
  XNOR2_X1 U340 ( .A(n474), .B(n473), .ZN(G1350GAT) );
  XOR2_X1 U341 ( .A(G183GAT), .B(KEYINPUT17), .Z(n293) );
  XNOR2_X1 U342 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n292) );
  XNOR2_X1 U343 ( .A(n293), .B(n292), .ZN(n435) );
  XOR2_X1 U344 ( .A(G120GAT), .B(G71GAT), .Z(n334) );
  XOR2_X1 U345 ( .A(n435), .B(n334), .Z(n295) );
  XNOR2_X1 U346 ( .A(G99GAT), .B(G134GAT), .ZN(n294) );
  XNOR2_X1 U347 ( .A(n295), .B(n294), .ZN(n301) );
  XOR2_X1 U348 ( .A(G127GAT), .B(KEYINPUT0), .Z(n297) );
  XNOR2_X1 U349 ( .A(G113GAT), .B(KEYINPUT80), .ZN(n296) );
  XNOR2_X1 U350 ( .A(n297), .B(n296), .ZN(n316) );
  XOR2_X1 U351 ( .A(n316), .B(KEYINPUT82), .Z(n299) );
  NAND2_X1 U352 ( .A1(G227GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U353 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U354 ( .A(n301), .B(n300), .Z(n309) );
  XOR2_X1 U355 ( .A(KEYINPUT83), .B(KEYINPUT20), .Z(n303) );
  XNOR2_X1 U356 ( .A(G43GAT), .B(G190GAT), .ZN(n302) );
  XNOR2_X1 U357 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U358 ( .A(G176GAT), .B(KEYINPUT81), .Z(n305) );
  XNOR2_X1 U359 ( .A(G169GAT), .B(G15GAT), .ZN(n304) );
  XNOR2_X1 U360 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U362 ( .A(n309), .B(n308), .Z(n541) );
  INV_X1 U363 ( .A(n541), .ZN(n546) );
  XOR2_X1 U364 ( .A(KEYINPUT93), .B(KEYINPUT1), .Z(n311) );
  XNOR2_X1 U365 ( .A(G120GAT), .B(G148GAT), .ZN(n310) );
  XNOR2_X1 U366 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U367 ( .A(G85GAT), .B(G155GAT), .Z(n313) );
  XNOR2_X1 U368 ( .A(G29GAT), .B(G162GAT), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U370 ( .A(n315), .B(n314), .ZN(n333) );
  XOR2_X1 U371 ( .A(KEYINPUT77), .B(G134GAT), .Z(n378) );
  XOR2_X1 U372 ( .A(n378), .B(n316), .Z(n318) );
  NAND2_X1 U373 ( .A1(G225GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U374 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U375 ( .A(n319), .B(KEYINPUT92), .Z(n323) );
  XOR2_X1 U376 ( .A(KEYINPUT86), .B(KEYINPUT3), .Z(n321) );
  XNOR2_X1 U377 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n320) );
  XNOR2_X1 U378 ( .A(n321), .B(n320), .ZN(n458) );
  XNOR2_X1 U379 ( .A(n458), .B(KEYINPUT6), .ZN(n322) );
  XNOR2_X1 U380 ( .A(n323), .B(n322), .ZN(n331) );
  XOR2_X1 U381 ( .A(KEYINPUT4), .B(KEYINPUT88), .Z(n325) );
  XNOR2_X1 U382 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n324) );
  XNOR2_X1 U383 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U384 ( .A(G57GAT), .B(KEYINPUT91), .Z(n327) );
  XNOR2_X1 U385 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n326) );
  XNOR2_X1 U386 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U387 ( .A(n329), .B(n328), .Z(n330) );
  XNOR2_X1 U388 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U389 ( .A(n333), .B(n332), .ZN(n536) );
  XOR2_X1 U390 ( .A(G57GAT), .B(KEYINPUT13), .Z(n355) );
  XNOR2_X1 U391 ( .A(n334), .B(n355), .ZN(n350) );
  XOR2_X1 U392 ( .A(G78GAT), .B(G148GAT), .Z(n336) );
  XNOR2_X1 U393 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n335) );
  XNOR2_X1 U394 ( .A(n336), .B(n335), .ZN(n456) );
  XOR2_X1 U395 ( .A(G64GAT), .B(G92GAT), .Z(n338) );
  XNOR2_X1 U396 ( .A(G176GAT), .B(G204GAT), .ZN(n337) );
  XNOR2_X1 U397 ( .A(n338), .B(n337), .ZN(n432) );
  XNOR2_X1 U398 ( .A(n456), .B(n432), .ZN(n342) );
  XOR2_X1 U399 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n340) );
  XNOR2_X1 U400 ( .A(KEYINPUT73), .B(KEYINPUT31), .ZN(n339) );
  XNOR2_X1 U401 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U402 ( .A(G99GAT), .B(G85GAT), .ZN(n343) );
  XNOR2_X1 U403 ( .A(n343), .B(KEYINPUT72), .ZN(n384) );
  INV_X1 U404 ( .A(KEYINPUT70), .ZN(n344) );
  XNOR2_X1 U405 ( .A(n384), .B(n344), .ZN(n346) );
  NAND2_X1 U406 ( .A1(G230GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U407 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U408 ( .A(n350), .B(n349), .ZN(n586) );
  XOR2_X1 U409 ( .A(G64GAT), .B(G183GAT), .Z(n352) );
  XNOR2_X1 U410 ( .A(G127GAT), .B(G71GAT), .ZN(n351) );
  XNOR2_X1 U411 ( .A(n352), .B(n351), .ZN(n368) );
  XOR2_X1 U412 ( .A(KEYINPUT15), .B(KEYINPUT78), .Z(n354) );
  XNOR2_X1 U413 ( .A(G8GAT), .B(KEYINPUT12), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n354), .B(n353), .ZN(n359) );
  XOR2_X1 U415 ( .A(n355), .B(G78GAT), .Z(n357) );
  XOR2_X1 U416 ( .A(G22GAT), .B(G155GAT), .Z(n454) );
  XNOR2_X1 U417 ( .A(G211GAT), .B(n454), .ZN(n356) );
  XNOR2_X1 U418 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U419 ( .A(n359), .B(n358), .Z(n361) );
  NAND2_X1 U420 ( .A1(G231GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U421 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U422 ( .A(n362), .B(KEYINPUT14), .Z(n366) );
  XOR2_X1 U423 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n364) );
  XNOR2_X1 U424 ( .A(G15GAT), .B(G1GAT), .ZN(n363) );
  XNOR2_X1 U425 ( .A(n364), .B(n363), .ZN(n396) );
  XNOR2_X1 U426 ( .A(n396), .B(KEYINPUT79), .ZN(n365) );
  XNOR2_X1 U427 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U428 ( .A(KEYINPUT67), .B(KEYINPUT7), .Z(n370) );
  XNOR2_X1 U429 ( .A(G43GAT), .B(G29GAT), .ZN(n369) );
  XNOR2_X1 U430 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U431 ( .A(KEYINPUT8), .B(n371), .Z(n408) );
  INV_X1 U432 ( .A(n408), .ZN(n391) );
  XOR2_X1 U433 ( .A(KEYINPUT65), .B(KEYINPUT74), .Z(n373) );
  XNOR2_X1 U434 ( .A(G218GAT), .B(KEYINPUT76), .ZN(n372) );
  XNOR2_X1 U435 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U436 ( .A(KEYINPUT10), .B(KEYINPUT75), .Z(n375) );
  XNOR2_X1 U437 ( .A(KEYINPUT11), .B(KEYINPUT9), .ZN(n374) );
  XNOR2_X1 U438 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U439 ( .A(n377), .B(n376), .Z(n383) );
  XOR2_X1 U440 ( .A(G36GAT), .B(G190GAT), .Z(n431) );
  XNOR2_X1 U441 ( .A(n378), .B(n431), .ZN(n381) );
  XOR2_X1 U442 ( .A(G50GAT), .B(G162GAT), .Z(n455) );
  AND2_X1 U443 ( .A1(G232GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U444 ( .A(n383), .B(n382), .ZN(n385) );
  XNOR2_X1 U445 ( .A(n385), .B(n384), .ZN(n387) );
  XOR2_X1 U446 ( .A(G106GAT), .B(G92GAT), .Z(n386) );
  NAND2_X1 U447 ( .A1(n387), .A2(n386), .ZN(n389) );
  OR2_X1 U448 ( .A1(n387), .A2(n386), .ZN(n388) );
  NAND2_X1 U449 ( .A1(n389), .A2(n388), .ZN(n390) );
  XOR2_X1 U450 ( .A(n391), .B(n390), .Z(n411) );
  XNOR2_X1 U451 ( .A(KEYINPUT36), .B(n411), .ZN(n590) );
  NAND2_X1 U452 ( .A1(n419), .A2(n590), .ZN(n394) );
  INV_X1 U453 ( .A(KEYINPUT45), .ZN(n392) );
  NOR2_X1 U454 ( .A1(n586), .A2(n395), .ZN(n410) );
  XOR2_X1 U455 ( .A(G169GAT), .B(G8GAT), .Z(n445) );
  XOR2_X1 U456 ( .A(n445), .B(n396), .Z(n398) );
  XNOR2_X1 U457 ( .A(G36GAT), .B(G50GAT), .ZN(n397) );
  XNOR2_X1 U458 ( .A(n398), .B(n397), .ZN(n402) );
  XOR2_X1 U459 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n400) );
  NAND2_X1 U460 ( .A1(G229GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U461 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U462 ( .A(n402), .B(n401), .Z(n407) );
  XOR2_X1 U463 ( .A(G113GAT), .B(G197GAT), .Z(n404) );
  XNOR2_X1 U464 ( .A(G141GAT), .B(G22GAT), .ZN(n403) );
  XNOR2_X1 U465 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U466 ( .A(n405), .B(KEYINPUT29), .ZN(n406) );
  XNOR2_X1 U467 ( .A(n407), .B(n406), .ZN(n409) );
  INV_X1 U468 ( .A(n583), .ZN(n501) );
  NAND2_X1 U469 ( .A1(n410), .A2(n501), .ZN(n424) );
  INV_X1 U470 ( .A(KEYINPUT64), .ZN(n412) );
  NAND2_X1 U471 ( .A1(n586), .A2(n412), .ZN(n415) );
  INV_X1 U472 ( .A(n586), .ZN(n413) );
  NAND2_X1 U473 ( .A1(n413), .A2(KEYINPUT64), .ZN(n414) );
  NAND2_X1 U474 ( .A1(n415), .A2(n414), .ZN(n416) );
  XNOR2_X2 U475 ( .A(n416), .B(KEYINPUT41), .ZN(n565) );
  NAND2_X1 U476 ( .A1(n583), .A2(n565), .ZN(n418) );
  XNOR2_X1 U477 ( .A(KEYINPUT108), .B(KEYINPUT46), .ZN(n417) );
  XNOR2_X1 U478 ( .A(n418), .B(n417), .ZN(n420) );
  INV_X1 U479 ( .A(n419), .ZN(n502) );
  NAND2_X1 U480 ( .A1(n420), .A2(n502), .ZN(n421) );
  NOR2_X1 U481 ( .A1(n411), .A2(n421), .ZN(n422) );
  XNOR2_X1 U482 ( .A(n422), .B(KEYINPUT47), .ZN(n423) );
  NAND2_X1 U483 ( .A1(n424), .A2(n423), .ZN(n426) );
  XNOR2_X1 U484 ( .A(KEYINPUT110), .B(KEYINPUT48), .ZN(n425) );
  XNOR2_X1 U485 ( .A(n426), .B(n425), .ZN(n543) );
  XNOR2_X1 U486 ( .A(G211GAT), .B(KEYINPUT84), .ZN(n427) );
  XNOR2_X1 U487 ( .A(n427), .B(KEYINPUT21), .ZN(n428) );
  XOR2_X1 U488 ( .A(n428), .B(KEYINPUT85), .Z(n430) );
  XNOR2_X1 U489 ( .A(G197GAT), .B(G218GAT), .ZN(n429) );
  XOR2_X1 U490 ( .A(n430), .B(n429), .Z(n466) );
  XNOR2_X1 U491 ( .A(n431), .B(n432), .ZN(n434) );
  AND2_X1 U492 ( .A1(G226GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U493 ( .A(n434), .B(n433), .ZN(n439) );
  XNOR2_X1 U494 ( .A(n435), .B(KEYINPUT96), .ZN(n437) );
  INV_X1 U495 ( .A(KEYINPUT94), .ZN(n436) );
  NAND2_X1 U496 ( .A1(n440), .A2(KEYINPUT95), .ZN(n444) );
  INV_X1 U497 ( .A(n440), .ZN(n442) );
  INV_X1 U498 ( .A(KEYINPUT95), .ZN(n441) );
  NAND2_X1 U499 ( .A1(n442), .A2(n441), .ZN(n443) );
  NAND2_X1 U500 ( .A1(n444), .A2(n443), .ZN(n447) );
  XOR2_X1 U501 ( .A(n445), .B(KEYINPUT78), .Z(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U503 ( .A(n466), .B(n448), .Z(n476) );
  XOR2_X1 U504 ( .A(KEYINPUT119), .B(n476), .Z(n449) );
  NAND2_X1 U505 ( .A1(n543), .A2(n449), .ZN(n452) );
  XOR2_X1 U506 ( .A(KEYINPUT54), .B(KEYINPUT120), .Z(n450) );
  NOR2_X1 U507 ( .A1(n536), .A2(n453), .ZN(n580) );
  XNOR2_X1 U508 ( .A(n455), .B(n454), .ZN(n457) );
  XNOR2_X1 U509 ( .A(n457), .B(n456), .ZN(n462) );
  XOR2_X1 U510 ( .A(n458), .B(KEYINPUT22), .Z(n460) );
  NAND2_X1 U511 ( .A1(G228GAT), .A2(G233GAT), .ZN(n459) );
  XNOR2_X1 U512 ( .A(n460), .B(n459), .ZN(n461) );
  XOR2_X1 U513 ( .A(n462), .B(n461), .Z(n468) );
  XOR2_X1 U514 ( .A(KEYINPUT87), .B(KEYINPUT23), .Z(n464) );
  XNOR2_X1 U515 ( .A(G204GAT), .B(KEYINPUT24), .ZN(n463) );
  XNOR2_X1 U516 ( .A(n464), .B(n463), .ZN(n465) );
  XOR2_X1 U517 ( .A(n466), .B(n465), .Z(n467) );
  XNOR2_X1 U518 ( .A(n468), .B(n467), .ZN(n479) );
  NAND2_X1 U519 ( .A1(n580), .A2(n479), .ZN(n470) );
  XOR2_X1 U520 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n469) );
  XNOR2_X1 U521 ( .A(n470), .B(n469), .ZN(n471) );
  NOR2_X2 U522 ( .A1(n546), .A2(n471), .ZN(n472) );
  XOR2_X2 U523 ( .A(KEYINPUT123), .B(n472), .Z(n575) );
  NAND2_X1 U524 ( .A1(n575), .A2(n419), .ZN(n474) );
  INV_X1 U525 ( .A(KEYINPUT105), .ZN(n494) );
  XOR2_X1 U526 ( .A(n479), .B(KEYINPUT28), .Z(n531) );
  XNOR2_X1 U527 ( .A(n476), .B(KEYINPUT27), .ZN(n481) );
  NAND2_X1 U528 ( .A1(n481), .A2(n536), .ZN(n561) );
  NOR2_X1 U529 ( .A1(n531), .A2(n561), .ZN(n544) );
  NAND2_X1 U530 ( .A1(n546), .A2(n544), .ZN(n475) );
  XNOR2_X1 U531 ( .A(n475), .B(KEYINPUT97), .ZN(n487) );
  NAND2_X1 U532 ( .A1(n541), .A2(n476), .ZN(n477) );
  NAND2_X1 U533 ( .A1(n479), .A2(n477), .ZN(n478) );
  XOR2_X1 U534 ( .A(KEYINPUT25), .B(n478), .Z(n483) );
  NOR2_X1 U535 ( .A1(n541), .A2(n479), .ZN(n480) );
  XNOR2_X1 U536 ( .A(n480), .B(KEYINPUT26), .ZN(n581) );
  NAND2_X1 U537 ( .A1(n481), .A2(n581), .ZN(n482) );
  NAND2_X1 U538 ( .A1(n483), .A2(n482), .ZN(n484) );
  XOR2_X1 U539 ( .A(KEYINPUT98), .B(n484), .Z(n485) );
  NOR2_X1 U540 ( .A1(n536), .A2(n485), .ZN(n486) );
  NOR2_X1 U541 ( .A1(n487), .A2(n486), .ZN(n488) );
  XNOR2_X1 U542 ( .A(n488), .B(KEYINPUT99), .ZN(n504) );
  AND2_X1 U543 ( .A1(n502), .A2(n504), .ZN(n489) );
  NAND2_X1 U544 ( .A1(n590), .A2(n489), .ZN(n492) );
  XNOR2_X1 U545 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n490) );
  NAND2_X1 U546 ( .A1(n565), .A2(n501), .ZN(n525) );
  NOR2_X1 U547 ( .A1(n514), .A2(n525), .ZN(n493) );
  XNOR2_X1 U548 ( .A(n494), .B(n493), .ZN(n540) );
  NAND2_X1 U549 ( .A1(n540), .A2(n531), .ZN(n497) );
  XOR2_X1 U550 ( .A(KEYINPUT107), .B(KEYINPUT44), .Z(n495) );
  XNOR2_X1 U551 ( .A(n497), .B(n496), .ZN(G1339GAT) );
  NAND2_X1 U552 ( .A1(n575), .A2(n565), .ZN(n500) );
  XOR2_X1 U553 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n498) );
  XNOR2_X1 U554 ( .A(n498), .B(G176GAT), .ZN(n499) );
  XNOR2_X1 U555 ( .A(n500), .B(n499), .ZN(G1349GAT) );
  OR2_X1 U556 ( .A1(n501), .A2(n586), .ZN(n515) );
  NOR2_X1 U557 ( .A1(n411), .A2(n502), .ZN(n503) );
  XNOR2_X1 U558 ( .A(n503), .B(KEYINPUT16), .ZN(n505) );
  NAND2_X1 U559 ( .A1(n505), .A2(n504), .ZN(n524) );
  NOR2_X1 U560 ( .A1(n515), .A2(n524), .ZN(n511) );
  NAND2_X1 U561 ( .A1(n536), .A2(n511), .ZN(n506) );
  XNOR2_X1 U562 ( .A(n506), .B(KEYINPUT34), .ZN(n507) );
  XNOR2_X1 U563 ( .A(G1GAT), .B(n507), .ZN(G1324GAT) );
  NAND2_X1 U564 ( .A1(n476), .A2(n511), .ZN(n508) );
  XNOR2_X1 U565 ( .A(n508), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U566 ( .A(G15GAT), .B(KEYINPUT35), .Z(n510) );
  NAND2_X1 U567 ( .A1(n511), .A2(n541), .ZN(n509) );
  XNOR2_X1 U568 ( .A(n510), .B(n509), .ZN(G1326GAT) );
  NAND2_X1 U569 ( .A1(n511), .A2(n531), .ZN(n512) );
  XNOR2_X1 U570 ( .A(n512), .B(KEYINPUT100), .ZN(n513) );
  XNOR2_X1 U571 ( .A(G22GAT), .B(n513), .ZN(G1327GAT) );
  XOR2_X1 U572 ( .A(G29GAT), .B(KEYINPUT39), .Z(n518) );
  NOR2_X1 U573 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U574 ( .A(n516), .B(KEYINPUT38), .ZN(n522) );
  NAND2_X1 U575 ( .A1(n522), .A2(n536), .ZN(n517) );
  XNOR2_X1 U576 ( .A(n518), .B(n517), .ZN(G1328GAT) );
  NAND2_X1 U577 ( .A1(n522), .A2(n476), .ZN(n519) );
  XNOR2_X1 U578 ( .A(n519), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U579 ( .A1(n522), .A2(n541), .ZN(n520) );
  XNOR2_X1 U580 ( .A(n520), .B(KEYINPUT40), .ZN(n521) );
  XNOR2_X1 U581 ( .A(G43GAT), .B(n521), .ZN(G1330GAT) );
  NAND2_X1 U582 ( .A1(n522), .A2(n531), .ZN(n523) );
  XNOR2_X1 U583 ( .A(n523), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT103), .B(KEYINPUT42), .Z(n527) );
  NOR2_X1 U585 ( .A1(n525), .A2(n524), .ZN(n532) );
  NAND2_X1 U586 ( .A1(n532), .A2(n536), .ZN(n526) );
  XNOR2_X1 U587 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U588 ( .A(G57GAT), .B(n528), .ZN(G1332GAT) );
  NAND2_X1 U589 ( .A1(n476), .A2(n532), .ZN(n529) );
  XNOR2_X1 U590 ( .A(n529), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U591 ( .A1(n541), .A2(n532), .ZN(n530) );
  XNOR2_X1 U592 ( .A(n530), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT43), .B(KEYINPUT104), .Z(n534) );
  NAND2_X1 U594 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U595 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U596 ( .A(G78GAT), .B(n535), .ZN(G1335GAT) );
  XNOR2_X1 U597 ( .A(G85GAT), .B(KEYINPUT106), .ZN(n538) );
  NAND2_X1 U598 ( .A1(n540), .A2(n536), .ZN(n537) );
  XNOR2_X1 U599 ( .A(n538), .B(n537), .ZN(G1336GAT) );
  NAND2_X1 U600 ( .A1(n476), .A2(n540), .ZN(n539) );
  XNOR2_X1 U601 ( .A(n539), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U602 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U603 ( .A(n542), .B(G99GAT), .ZN(G1338GAT) );
  BUF_X1 U604 ( .A(n543), .Z(n559) );
  NAND2_X1 U605 ( .A1(n544), .A2(n559), .ZN(n545) );
  NOR2_X1 U606 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U607 ( .A(KEYINPUT111), .B(n547), .Z(n555) );
  NAND2_X1 U608 ( .A1(n555), .A2(n583), .ZN(n548) );
  XNOR2_X1 U609 ( .A(n548), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT49), .B(KEYINPUT112), .Z(n550) );
  NAND2_X1 U611 ( .A1(n555), .A2(n565), .ZN(n549) );
  XNOR2_X1 U612 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U613 ( .A(G120GAT), .B(n551), .ZN(G1341GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT50), .B(KEYINPUT113), .Z(n553) );
  NAND2_X1 U615 ( .A1(n555), .A2(n419), .ZN(n552) );
  XNOR2_X1 U616 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U617 ( .A(G127GAT), .B(n554), .ZN(G1342GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n557) );
  NAND2_X1 U619 ( .A1(n555), .A2(n411), .ZN(n556) );
  XNOR2_X1 U620 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U621 ( .A(G134GAT), .B(n558), .ZN(G1343GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n563) );
  NAND2_X1 U623 ( .A1(n559), .A2(n581), .ZN(n560) );
  NOR2_X1 U624 ( .A1(n561), .A2(n560), .ZN(n572) );
  NAND2_X1 U625 ( .A1(n572), .A2(n583), .ZN(n562) );
  XNOR2_X1 U626 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U627 ( .A(G141GAT), .B(n564), .ZN(G1344GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT117), .B(KEYINPUT53), .Z(n567) );
  NAND2_X1 U629 ( .A1(n572), .A2(n565), .ZN(n566) );
  XNOR2_X1 U630 ( .A(n567), .B(n566), .ZN(n569) );
  XOR2_X1 U631 ( .A(G148GAT), .B(KEYINPUT52), .Z(n568) );
  XNOR2_X1 U632 ( .A(n569), .B(n568), .ZN(G1345GAT) );
  NAND2_X1 U633 ( .A1(n572), .A2(n419), .ZN(n570) );
  XNOR2_X1 U634 ( .A(n570), .B(KEYINPUT118), .ZN(n571) );
  XNOR2_X1 U635 ( .A(G155GAT), .B(n571), .ZN(G1346GAT) );
  NAND2_X1 U636 ( .A1(n411), .A2(n572), .ZN(n573) );
  XNOR2_X1 U637 ( .A(n573), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U638 ( .A1(n575), .A2(n583), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n411), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(KEYINPUT58), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n577), .B(G190GAT), .ZN(G1351GAT) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n578), .B(KEYINPUT60), .ZN(n579) );
  XOR2_X1 U645 ( .A(KEYINPUT59), .B(n579), .Z(n585) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(KEYINPUT125), .ZN(n591) );
  NAND2_X1 U648 ( .A1(n591), .A2(n583), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(G1352GAT) );
  XOR2_X1 U650 ( .A(G204GAT), .B(KEYINPUT61), .Z(n588) );
  NAND2_X1 U651 ( .A1(n591), .A2(n586), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(G1353GAT) );
  NAND2_X1 U653 ( .A1(n591), .A2(n419), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n589), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(n592), .B(KEYINPUT62), .ZN(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

