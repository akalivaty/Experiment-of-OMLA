//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n823, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n911, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT71), .B(G197gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT22), .ZN(new_n205));
  NAND2_X1  g004(.A1(G211gat), .A2(G218gat), .ZN(new_n206));
  AOI22_X1  g005(.A1(new_n204), .A2(G204gat), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n207), .B1(G204gat), .B2(new_n204), .ZN(new_n208));
  XOR2_X1   g007(.A(G211gat), .B(G218gat), .Z(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n209), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n207), .B(new_n211), .C1(G204gat), .C2(new_n204), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT29), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT3), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT76), .ZN(new_n216));
  XNOR2_X1  g015(.A(G155gat), .B(G162gat), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G141gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G148gat), .ZN(new_n220));
  INV_X1    g019(.A(G148gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G141gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n220), .A2(new_n222), .B1(KEYINPUT2), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT75), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n216), .B(new_n218), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n223), .A2(KEYINPUT2), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n221), .A2(G141gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n219), .A2(G148gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT76), .B1(new_n230), .B2(KEYINPUT75), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n217), .B1(new_n224), .B2(new_n216), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n226), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT78), .ZN(new_n234));
  XNOR2_X1  g033(.A(G141gat), .B(G148gat), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n223), .A2(KEYINPUT2), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT76), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n225), .B1(new_n238), .B2(new_n227), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n237), .B(new_n217), .C1(new_n239), .C2(KEYINPUT76), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT78), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(new_n241), .A3(new_n226), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n234), .A2(new_n242), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n215), .A2(new_n243), .ZN(new_n244));
  AOI211_X1 g043(.A(KEYINPUT77), .B(KEYINPUT3), .C1(new_n240), .C2(new_n226), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT77), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n246), .B1(new_n233), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n214), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n213), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT81), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n244), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n249), .A2(KEYINPUT81), .A3(new_n250), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n203), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n251), .B(new_n203), .C1(new_n233), .C2(new_n215), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(G22gat), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT82), .B(G22gat), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n249), .A2(KEYINPUT81), .A3(new_n250), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT81), .B1(new_n249), .B2(new_n250), .ZN(new_n262));
  NOR3_X1   g061(.A1(new_n261), .A2(new_n262), .A3(new_n244), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n256), .B(new_n260), .C1(new_n263), .C2(new_n203), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(G50gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(G78gat), .B(G106gat), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n266), .B(new_n267), .Z(new_n268));
  NAND3_X1  g067(.A1(new_n258), .A2(new_n264), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT83), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT83), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n258), .A2(new_n264), .A3(new_n271), .A4(new_n268), .ZN(new_n272));
  INV_X1    g071(.A(new_n268), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n253), .A2(new_n254), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(new_n202), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n260), .B1(new_n275), .B2(new_n256), .ZN(new_n276));
  NOR3_X1   g075(.A1(new_n255), .A2(new_n257), .A3(new_n259), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n273), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n270), .A2(new_n272), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT25), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT64), .B(G169gat), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT23), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n282), .A2(G176gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(G183gat), .A2(G190gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT24), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OR2_X1    g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT65), .ZN(new_n292));
  NOR2_X1   g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n292), .B1(new_n293), .B2(KEYINPUT23), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n282), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n280), .B1(new_n291), .B2(new_n297), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT66), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n290), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n280), .B1(new_n293), .B2(KEYINPUT23), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n287), .A2(new_n288), .A3(KEYINPUT66), .A4(new_n289), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n299), .A2(new_n301), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n298), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT27), .B(G183gat), .ZN(new_n306));
  INV_X1    g105(.A(G190gat), .ZN(new_n307));
  AND2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT28), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n308), .A2(new_n309), .B1(G183gat), .B2(G190gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n293), .B(KEYINPUT26), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n306), .A2(new_n307), .ZN(new_n312));
  AOI22_X1  g111(.A1(new_n296), .A2(new_n311), .B1(new_n312), .B2(KEYINPUT28), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n305), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(G226gat), .ZN(new_n316));
  INV_X1    g115(.A(G233gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n315), .A2(KEYINPUT72), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n318), .ZN(new_n320));
  AOI22_X1  g119(.A1(new_n298), .A2(new_n304), .B1(new_n310), .B2(new_n313), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n320), .B1(new_n321), .B2(KEYINPUT29), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT72), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n323), .B1(new_n321), .B2(new_n320), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n319), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n250), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT73), .B1(new_n315), .B2(new_n318), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n328));
  NOR3_X1   g127(.A1(new_n321), .A2(new_n328), .A3(new_n320), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n213), .B(new_n322), .C1(new_n327), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G64gat), .B(G92gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(KEYINPUT74), .ZN(new_n333));
  XNOR2_X1  g132(.A(G8gat), .B(G36gat), .ZN(new_n334));
  XOR2_X1   g133(.A(new_n333), .B(new_n334), .Z(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n326), .A2(new_n330), .A3(new_n335), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(KEYINPUT30), .A3(new_n338), .ZN(new_n339));
  AND3_X1   g138(.A1(new_n326), .A2(new_n330), .A3(new_n335), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n335), .B1(new_n326), .B2(new_n330), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT30), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(G134gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(G127gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT67), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT67), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n349), .A2(new_n346), .A3(G127gat), .ZN(new_n350));
  INV_X1    g149(.A(G127gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G134gat), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n348), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT1), .ZN(new_n354));
  INV_X1    g153(.A(G113gat), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n355), .A2(G120gat), .ZN(new_n356));
  INV_X1    g155(.A(G120gat), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n357), .A2(G113gat), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n354), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n353), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT68), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n361), .B1(new_n357), .B2(G113gat), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n355), .A2(KEYINPUT68), .A3(G120gat), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n362), .B(new_n363), .C1(new_n355), .C2(G120gat), .ZN(new_n364));
  AND3_X1   g163(.A1(new_n347), .A2(new_n352), .A3(new_n354), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n360), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n233), .B(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT5), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n367), .B1(new_n233), .B2(new_n247), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n233), .A2(new_n247), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT77), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n233), .A2(new_n246), .A3(new_n247), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n377), .A2(new_n370), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT4), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n359), .A2(new_n353), .B1(new_n364), .B2(new_n365), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n233), .A2(KEYINPUT79), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT79), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n233), .A2(new_n380), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n382), .B1(new_n383), .B2(KEYINPUT4), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n367), .A2(KEYINPUT69), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT69), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n234), .A2(new_n242), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n381), .B(new_n384), .C1(new_n388), .C2(new_n379), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n378), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n369), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n383), .A2(new_n379), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n385), .A2(new_n387), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n243), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n392), .B1(new_n394), .B2(new_n379), .ZN(new_n395));
  INV_X1    g194(.A(new_n377), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT5), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n372), .B1(new_n391), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G1gat), .B(G29gat), .ZN(new_n399));
  INV_X1    g198(.A(G85gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n399), .B(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(KEYINPUT0), .B(G57gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  XOR2_X1   g202(.A(new_n403), .B(KEYINPUT84), .Z(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT39), .ZN(new_n406));
  INV_X1    g205(.A(new_n369), .ZN(new_n407));
  INV_X1    g206(.A(new_n392), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n408), .B1(new_n388), .B2(KEYINPUT4), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n406), .B(new_n407), .C1(new_n409), .C2(new_n377), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n369), .B1(new_n395), .B2(new_n396), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n368), .A2(new_n369), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT39), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n410), .B(new_n404), .C1(new_n411), .C2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT40), .ZN(new_n415));
  AOI22_X1  g214(.A1(new_n398), .A2(new_n405), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n407), .B1(new_n409), .B2(new_n377), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n417), .A2(KEYINPUT39), .A3(new_n412), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n418), .A2(KEYINPUT40), .A3(new_n404), .A4(new_n410), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n345), .A2(new_n416), .A3(KEYINPUT85), .A4(new_n419), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n403), .B(new_n372), .C1(new_n391), .C2(new_n397), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT6), .ZN(new_n422));
  INV_X1    g221(.A(new_n397), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n407), .B1(new_n378), .B2(new_n389), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n423), .A2(new_n424), .B1(new_n368), .B2(new_n371), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n421), .B(new_n422), .C1(new_n425), .C2(new_n404), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n336), .B1(new_n331), .B2(KEYINPUT37), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT37), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n429), .B1(new_n325), .B2(new_n213), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n250), .B(new_n322), .C1(new_n327), .C2(new_n329), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT38), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n340), .B1(new_n428), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n403), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n398), .A2(KEYINPUT6), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n429), .B1(new_n326), .B2(new_n330), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT38), .B1(new_n427), .B2(new_n436), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n426), .A2(new_n433), .A3(new_n435), .A4(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT85), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n414), .A2(new_n415), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n440), .B(new_n419), .C1(new_n425), .C2(new_n404), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n439), .B1(new_n441), .B2(new_n344), .ZN(new_n442));
  AND4_X1   g241(.A1(new_n279), .A2(new_n420), .A3(new_n438), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n315), .A2(new_n393), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n321), .A2(new_n385), .A3(new_n387), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n444), .A2(new_n445), .A3(G227gat), .A4(G233gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT32), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT70), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n446), .A2(KEYINPUT70), .A3(KEYINPUT32), .ZN(new_n450));
  XNOR2_X1  g249(.A(G15gat), .B(G43gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(G71gat), .B(G99gat), .ZN(new_n452));
  XOR2_X1   g251(.A(new_n451), .B(new_n452), .Z(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT33), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n454), .B1(new_n446), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n449), .A2(new_n450), .A3(new_n456), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n446), .B(KEYINPUT32), .C1(new_n455), .C2(new_n454), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n445), .ZN(new_n460));
  NAND2_X1  g259(.A1(G227gat), .A2(G233gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AND2_X1   g261(.A1(new_n462), .A2(KEYINPUT34), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n462), .A2(KEYINPUT34), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n459), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n463), .A2(new_n464), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n457), .A2(new_n466), .A3(new_n458), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT36), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n465), .A2(KEYINPUT36), .A3(new_n467), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n398), .A2(new_n434), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n473), .A2(new_n422), .A3(new_n421), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n345), .B1(new_n474), .B2(new_n435), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n472), .B1(new_n279), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n443), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(KEYINPUT86), .B(KEYINPUT35), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n344), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n479), .B1(new_n435), .B2(new_n426), .ZN(new_n480));
  INV_X1    g279(.A(new_n468), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n480), .A2(new_n279), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n279), .A2(new_n475), .A3(new_n481), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT35), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n482), .B1(new_n484), .B2(KEYINPUT87), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT87), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n483), .A2(new_n486), .A3(KEYINPUT35), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n477), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(G57gat), .B(G64gat), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT94), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(G71gat), .A2(G78gat), .ZN(new_n492));
  INV_X1    g291(.A(G71gat), .ZN(new_n493));
  INV_X1    g292(.A(G78gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT9), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n492), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n489), .A2(new_n490), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n491), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n492), .B(new_n495), .C1(new_n489), .C2(new_n496), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT21), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G127gat), .B(G155gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  XOR2_X1   g304(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n506));
  XNOR2_X1  g305(.A(G183gat), .B(G211gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n505), .B(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G15gat), .B(G22gat), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT16), .ZN(new_n511));
  AOI21_X1  g310(.A(G1gat), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(KEYINPUT91), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(KEYINPUT92), .A2(G8gat), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n510), .B(KEYINPUT91), .C1(new_n511), .C2(G1gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(KEYINPUT92), .A2(G8gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n518), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n514), .A2(new_n520), .A3(new_n515), .A4(new_n516), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(new_n502), .B2(new_n501), .ZN(new_n523));
  NAND2_X1  g322(.A1(G231gat), .A2(G233gat), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n524), .B(KEYINPUT95), .Z(new_n525));
  XNOR2_X1  g324(.A(new_n523), .B(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n509), .B(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT7), .ZN(new_n528));
  INV_X1    g327(.A(G92gat), .ZN(new_n529));
  OAI211_X1 g328(.A(KEYINPUT96), .B(new_n528), .C1(new_n400), .C2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT96), .ZN(new_n531));
  OAI211_X1 g330(.A(G85gat), .B(G92gat), .C1(new_n531), .C2(KEYINPUT7), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n528), .A2(KEYINPUT96), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(KEYINPUT97), .B(G85gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n529), .ZN(new_n536));
  NAND2_X1  g335(.A1(G99gat), .A2(G106gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT8), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT98), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n535), .A2(new_n529), .B1(KEYINPUT8), .B2(new_n537), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT98), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n534), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G99gat), .B(G106gat), .Z(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G43gat), .B(G50gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT15), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  OR3_X1    g348(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(KEYINPUT89), .ZN(new_n553));
  NAND2_X1  g352(.A1(G29gat), .A2(G36gat), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT89), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n554), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n549), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n547), .A2(KEYINPUT15), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n554), .B(KEYINPUT90), .Z(new_n559));
  NAND4_X1  g358(.A1(new_n558), .A2(new_n559), .A3(new_n548), .A4(new_n552), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT17), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n557), .A2(KEYINPUT17), .A3(new_n560), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT99), .B1(new_n546), .B2(new_n565), .ZN(new_n566));
  AND3_X1   g365(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n567), .B1(new_n546), .B2(new_n561), .ZN(new_n568));
  INV_X1    g367(.A(new_n534), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n539), .A2(KEYINPUT98), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n541), .A2(new_n542), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(new_n545), .ZN(new_n573));
  INV_X1    g372(.A(new_n545), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n574), .B(new_n569), .C1(new_n570), .C2(new_n571), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT99), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n576), .A2(new_n577), .A3(new_n563), .A4(new_n564), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n566), .A2(new_n568), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G190gat), .B(G218gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT100), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT101), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n581), .A2(new_n582), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n585), .B(new_n586), .Z(new_n587));
  XOR2_X1   g386(.A(G134gat), .B(G162gat), .Z(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n579), .A2(new_n583), .A3(new_n589), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G230gat), .A2(G233gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT102), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n501), .B1(new_n575), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n576), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n573), .B(new_n575), .C1(new_n595), .C2(new_n501), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT10), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT10), .ZN(new_n600));
  NOR3_X1   g399(.A1(new_n576), .A2(new_n600), .A3(new_n501), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n594), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n594), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n597), .A2(new_n603), .A3(new_n598), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G176gat), .B(G204gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT103), .ZN(new_n607));
  XOR2_X1   g406(.A(G120gat), .B(G148gat), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n605), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n522), .A2(new_n557), .A3(new_n560), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n519), .A2(new_n561), .A3(new_n521), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n614), .A2(KEYINPUT93), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G229gat), .A2(G233gat), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n617), .B(KEYINPUT13), .Z(new_n618));
  INV_X1    g417(.A(KEYINPUT93), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n519), .A2(new_n561), .A3(new_n619), .A4(new_n521), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n616), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n522), .A2(new_n563), .A3(new_n564), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n622), .A2(new_n617), .A3(new_n615), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT18), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n622), .A2(KEYINPUT18), .A3(new_n617), .A4(new_n615), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n621), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G113gat), .B(G141gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(G197gat), .ZN(new_n629));
  XOR2_X1   g428(.A(KEYINPUT11), .B(G169gat), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  AND3_X1   g431(.A1(new_n627), .A2(KEYINPUT88), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n632), .B1(new_n627), .B2(KEYINPUT88), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n613), .A2(new_n635), .ZN(new_n636));
  NOR4_X1   g435(.A1(new_n488), .A2(new_n527), .A3(new_n593), .A4(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n474), .A2(new_n435), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G1gat), .ZN(G1324gat));
  INV_X1    g440(.A(KEYINPUT104), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n637), .A2(new_n345), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT16), .B(G8gat), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n645), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n643), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(KEYINPUT42), .B2(new_n645), .ZN(G1325gat));
  AOI21_X1  g446(.A(G15gat), .B1(new_n637), .B2(new_n481), .ZN(new_n648));
  INV_X1    g447(.A(new_n472), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n649), .A2(G15gat), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n648), .B1(new_n637), .B2(new_n650), .ZN(G1326gat));
  INV_X1    g450(.A(new_n279), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT43), .B(G22gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(G1327gat));
  NAND2_X1  g454(.A1(new_n484), .A2(KEYINPUT87), .ZN(new_n656));
  INV_X1    g455(.A(new_n482), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n656), .A2(new_n657), .A3(new_n487), .ZN(new_n658));
  INV_X1    g457(.A(new_n477), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n527), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n636), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n660), .A2(new_n593), .A3(new_n662), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n663), .A2(G29gat), .A3(new_n638), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n664), .B(KEYINPUT45), .Z(new_n665));
  INV_X1    g464(.A(KEYINPUT108), .ZN(new_n666));
  INV_X1    g465(.A(new_n593), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT44), .B1(new_n488), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT106), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n579), .A2(new_n583), .A3(new_n589), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n589), .B1(new_n579), .B2(new_n583), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n591), .A2(KEYINPUT106), .A3(new_n592), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(KEYINPUT44), .ZN(new_n675));
  INV_X1    g474(.A(new_n487), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n486), .B1(new_n483), .B2(KEYINPUT35), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n676), .A2(new_n677), .A3(new_n482), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n675), .B1(new_n678), .B2(new_n477), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n668), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n662), .B(KEYINPUT105), .Z(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(KEYINPUT107), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT107), .ZN(new_n684));
  AOI211_X1 g483(.A(new_n684), .B(new_n681), .C1(new_n668), .C2(new_n679), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n666), .B(new_n639), .C1(new_n683), .C2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(G29gat), .ZN(new_n687));
  INV_X1    g486(.A(new_n675), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n688), .B1(new_n658), .B2(new_n659), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n660), .A2(new_n593), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n689), .B1(new_n690), .B2(KEYINPUT44), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n684), .B1(new_n691), .B2(new_n681), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n680), .A2(KEYINPUT107), .A3(new_n682), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n666), .B1(new_n694), .B2(new_n639), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n665), .B1(new_n687), .B2(new_n695), .ZN(G1328gat));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n345), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(G36gat), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n663), .A2(G36gat), .A3(new_n344), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT46), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(G1329gat));
  NAND2_X1  g500(.A1(new_n680), .A2(new_n682), .ZN(new_n702));
  OAI21_X1  g501(.A(G43gat), .B1(new_n702), .B2(new_n472), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n663), .A2(G43gat), .A3(new_n468), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT47), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n649), .B1(new_n683), .B2(new_n685), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n704), .B1(new_n708), .B2(G43gat), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n707), .B1(new_n709), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g509(.A(G50gat), .B1(new_n702), .B2(new_n279), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n279), .A2(G50gat), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n711), .B(KEYINPUT48), .C1(new_n663), .C2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n663), .A2(new_n712), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n652), .B1(new_n683), .B2(new_n685), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n714), .B1(new_n715), .B2(G50gat), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n713), .B1(new_n716), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g516(.A(new_n635), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n593), .A2(new_n527), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n488), .A2(new_n613), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n639), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT109), .B(G57gat), .Z(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1332gat));
  INV_X1    g523(.A(new_n721), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(new_n344), .ZN(new_n726));
  NOR2_X1   g525(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n727));
  AND2_X1   g526(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n729), .B1(new_n726), .B2(new_n727), .ZN(G1333gat));
  OAI21_X1  g529(.A(new_n493), .B1(new_n725), .B2(new_n468), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n721), .A2(G71gat), .A3(new_n649), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g533(.A1(new_n721), .A2(new_n652), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g535(.A1(new_n635), .A2(new_n661), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n660), .A2(new_n593), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT51), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n639), .A2(new_n535), .A3(new_n612), .ZN(new_n742));
  INV_X1    g541(.A(new_n737), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n613), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n680), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n745), .A2(new_n638), .ZN(new_n746));
  OAI22_X1  g545(.A1(new_n741), .A2(new_n742), .B1(new_n746), .B2(new_n535), .ZN(G1336gat));
  NOR3_X1   g546(.A1(new_n613), .A2(G92gat), .A3(new_n344), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n740), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n745), .A2(new_n344), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n750), .B2(new_n529), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT52), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n749), .B(new_n753), .C1(new_n529), .C2(new_n750), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(G1337gat));
  NOR3_X1   g554(.A1(new_n613), .A2(new_n468), .A3(G99gat), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT110), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n680), .A2(new_n758), .A3(new_n649), .A4(new_n744), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G99gat), .ZN(new_n760));
  INV_X1    g559(.A(new_n744), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n761), .B1(new_n668), .B2(new_n679), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n758), .B1(new_n762), .B2(new_n649), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n757), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT111), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT111), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n757), .B(new_n766), .C1(new_n760), .C2(new_n763), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(G1338gat));
  NOR2_X1   g567(.A1(KEYINPUT112), .A2(KEYINPUT53), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(G106gat), .B1(new_n745), .B2(new_n279), .ZN(new_n771));
  NAND2_X1  g570(.A1(KEYINPUT112), .A2(KEYINPUT53), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n279), .A2(G106gat), .A3(new_n613), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n738), .A2(new_n739), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n738), .A2(new_n739), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AND4_X1   g575(.A1(new_n770), .A2(new_n771), .A3(new_n772), .A4(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n772), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n778), .B1(new_n740), .B2(new_n773), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n770), .B1(new_n779), .B2(new_n771), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n777), .A2(new_n780), .ZN(G1339gat));
  INV_X1    g580(.A(new_n674), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n597), .A2(new_n598), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n600), .ZN(new_n785));
  INV_X1    g584(.A(new_n601), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n785), .A2(new_n603), .A3(new_n786), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n787), .A2(KEYINPUT54), .A3(new_n602), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n789), .B(new_n594), .C1(new_n599), .C2(new_n601), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n609), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n783), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n790), .A2(new_n609), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n787), .A2(KEYINPUT54), .A3(new_n602), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n793), .A2(KEYINPUT55), .A3(new_n794), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n792), .A2(new_n635), .A3(new_n610), .A4(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n618), .B1(new_n616), .B2(new_n620), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n617), .B1(new_n622), .B2(new_n615), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n631), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n621), .A2(new_n625), .A3(new_n626), .A4(new_n632), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n612), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n782), .B1(new_n796), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n795), .A2(new_n610), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT55), .B1(new_n793), .B2(new_n794), .ZN(new_n806));
  NOR4_X1   g605(.A1(new_n805), .A2(new_n674), .A3(new_n806), .A4(new_n801), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n527), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n720), .A2(new_n612), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n638), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n811), .A2(new_n279), .A3(new_n481), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n812), .A2(new_n344), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(G113gat), .B1(new_n814), .B2(new_n718), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n635), .A2(new_n355), .ZN(new_n816));
  XOR2_X1   g615(.A(new_n816), .B(KEYINPUT113), .Z(new_n817));
  OAI21_X1  g616(.A(new_n815), .B1(new_n814), .B2(new_n817), .ZN(G1340gat));
  OAI21_X1  g617(.A(G120gat), .B1(new_n814), .B2(new_n613), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n612), .A2(new_n357), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(KEYINPUT114), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n814), .B2(new_n821), .ZN(G1341gat));
  NAND2_X1  g621(.A1(new_n813), .A2(new_n661), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(G127gat), .ZN(G1342gat));
  AOI21_X1  g623(.A(new_n346), .B1(new_n813), .B2(new_n593), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n344), .A2(new_n593), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT115), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n812), .A2(new_n346), .A3(new_n828), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(KEYINPUT116), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT56), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n825), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n831), .A2(KEYINPUT117), .A3(new_n832), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n835), .B1(new_n830), .B2(KEYINPUT56), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n833), .B1(new_n834), .B2(new_n836), .ZN(G1343gat));
  AND2_X1   g636(.A1(new_n811), .A2(KEYINPUT119), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n649), .A2(new_n279), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n839), .B1(new_n811), .B2(KEYINPUT119), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT121), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n718), .A2(G141gat), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n344), .A3(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n649), .A2(new_n638), .A3(new_n345), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n808), .A2(new_n810), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT57), .B1(new_n847), .B2(new_n652), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n279), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n593), .B1(new_n796), .B2(new_n803), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n527), .B1(new_n852), .B2(new_n807), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n851), .B1(new_n853), .B2(new_n810), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n846), .B1(new_n848), .B2(new_n854), .ZN(new_n855));
  OR3_X1    g654(.A1(new_n855), .A2(KEYINPUT122), .A3(new_n718), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT122), .B1(new_n855), .B2(new_n718), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n856), .A2(G141gat), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n844), .A2(new_n845), .A3(new_n858), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n841), .A2(new_n344), .A3(new_n843), .ZN(new_n860));
  OAI211_X1 g659(.A(KEYINPUT118), .B(new_n846), .C1(new_n848), .C2(new_n854), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n853), .A2(new_n810), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n850), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n279), .B1(new_n808), .B2(new_n810), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(KEYINPUT57), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT118), .B1(new_n866), .B2(new_n846), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n635), .B1(new_n862), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n860), .B1(new_n868), .B2(G141gat), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT120), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n869), .A2(new_n870), .A3(new_n845), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n841), .A2(new_n344), .A3(new_n843), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n855), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n718), .B1(new_n874), .B2(new_n861), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n872), .B1(new_n875), .B2(new_n219), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT120), .B1(new_n876), .B2(KEYINPUT58), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n859), .B1(new_n871), .B2(new_n877), .ZN(G1344gat));
  NAND4_X1  g677(.A1(new_n842), .A2(new_n221), .A3(new_n344), .A4(new_n612), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n805), .A2(new_n806), .A3(new_n801), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n796), .A2(new_n803), .ZN(new_n882));
  MUX2_X1   g681(.A(new_n881), .B(new_n882), .S(new_n667), .Z(new_n883));
  AOI21_X1  g682(.A(new_n809), .B1(new_n883), .B2(new_n527), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n849), .B1(new_n884), .B2(new_n279), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n885), .A2(KEYINPUT123), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(KEYINPUT123), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n865), .A2(KEYINPUT57), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n612), .A3(new_n846), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n880), .B1(new_n890), .B2(G148gat), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n874), .A2(new_n861), .ZN(new_n892));
  AOI211_X1 g691(.A(KEYINPUT59), .B(new_n221), .C1(new_n892), .C2(new_n612), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n879), .B1(new_n891), .B2(new_n893), .ZN(G1345gat));
  NAND3_X1  g693(.A1(new_n842), .A2(new_n344), .A3(new_n661), .ZN(new_n895));
  INV_X1    g694(.A(G155gat), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n527), .A2(new_n896), .ZN(new_n897));
  AOI22_X1  g696(.A1(new_n895), .A2(new_n896), .B1(new_n892), .B2(new_n897), .ZN(G1346gat));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n827), .A2(G162gat), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n842), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n899), .B1(new_n842), .B2(new_n900), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT125), .B1(new_n892), .B2(new_n782), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n892), .A2(KEYINPUT125), .A3(new_n782), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(G162gat), .ZN(new_n905));
  OAI22_X1  g704(.A1(new_n901), .A2(new_n902), .B1(new_n903), .B2(new_n905), .ZN(G1347gat));
  AOI21_X1  g705(.A(new_n639), .B1(new_n808), .B2(new_n810), .ZN(new_n907));
  AND4_X1   g706(.A1(new_n345), .A2(new_n907), .A3(new_n279), .A4(new_n481), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n635), .ZN(new_n909));
  MUX2_X1   g708(.A(new_n281), .B(G169gat), .S(new_n909), .Z(G1348gat));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n612), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g711(.A1(new_n908), .A2(new_n661), .ZN(new_n913));
  MUX2_X1   g712(.A(new_n306), .B(G183gat), .S(new_n913), .Z(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g714(.A(new_n307), .B1(new_n908), .B2(new_n593), .ZN(new_n916));
  XOR2_X1   g715(.A(new_n916), .B(KEYINPUT61), .Z(new_n917));
  NAND3_X1  g716(.A1(new_n908), .A2(new_n307), .A3(new_n782), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1351gat));
  INV_X1    g718(.A(KEYINPUT126), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n889), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n886), .A2(KEYINPUT126), .A3(new_n887), .A4(new_n888), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n649), .A2(new_n639), .A3(new_n344), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(G197gat), .B1(new_n924), .B2(new_n718), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n907), .A2(new_n345), .A3(new_n839), .ZN(new_n926));
  OR3_X1    g725(.A1(new_n926), .A2(G197gat), .A3(new_n718), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1352gat));
  XNOR2_X1  g727(.A(KEYINPUT127), .B(G204gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n929), .B1(new_n924), .B2(new_n613), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n926), .A2(new_n613), .A3(new_n929), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT62), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(G1353gat));
  OR3_X1    g732(.A1(new_n926), .A2(G211gat), .A3(new_n527), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n889), .A2(new_n661), .A3(new_n923), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n935), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n936));
  AOI21_X1  g735(.A(KEYINPUT63), .B1(new_n935), .B2(G211gat), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(G1354gat));
  INV_X1    g737(.A(G218gat), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n667), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n921), .A2(new_n922), .A3(new_n923), .A4(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n939), .B1(new_n926), .B2(new_n674), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(G1355gat));
endmodule


