//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 0 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n616, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT66), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT67), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT68), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(G567), .A2(new_n455), .B1(new_n452), .B2(G2106), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(G125), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n464), .A2(new_n469), .ZN(G160));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(new_n466), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n459), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n459), .A2(G112), .ZN(new_n476));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n472), .A2(new_n473), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(new_n459), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n478), .B1(G136), .B2(new_n481), .ZN(new_n482));
  XNOR2_X1  g057(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n482), .B(new_n483), .ZN(G162));
  NAND2_X1  g059(.A1(KEYINPUT4), .A2(G138), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n485), .B1(new_n472), .B2(new_n473), .ZN(new_n486));
  AND2_X1   g061(.A1(G102), .A2(G2104), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n459), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G126), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n489), .B1(new_n472), .B2(new_n473), .ZN(new_n490));
  AND2_X1   g065(.A1(G114), .A2(G2104), .ZN(new_n491));
  OAI21_X1  g066(.A(G2105), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI211_X1 g067(.A(G138), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n488), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  OR2_X1    g073(.A1(KEYINPUT6), .A2(G651), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT6), .A2(G651), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G50), .ZN(new_n502));
  INV_X1    g077(.A(G88), .ZN(new_n503));
  OR2_X1    g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n499), .A2(new_n500), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n502), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n509), .A2(new_n512), .ZN(G166));
  NAND2_X1  g088(.A1(new_n501), .A2(G51), .ZN(new_n514));
  XOR2_X1   g089(.A(KEYINPUT71), .B(G89), .Z(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n508), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n517));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT7), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n516), .A2(new_n520), .ZN(G286));
  INV_X1    g096(.A(G286), .ZN(G168));
  NAND2_X1  g097(.A1(new_n501), .A2(G52), .ZN(new_n523));
  INV_X1    g098(.A(G90), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n508), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n523), .B(KEYINPUT73), .C1(new_n524), .C2(new_n508), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT74), .ZN(new_n530));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  AND2_X1   g106(.A1(KEYINPUT5), .A2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(KEYINPUT5), .A2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(G64), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n531), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT72), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n536), .A2(new_n539), .A3(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AND3_X1   g116(.A1(new_n529), .A2(new_n530), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n530), .B1(new_n529), .B2(new_n541), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n542), .A2(new_n543), .ZN(G171));
  AOI22_X1  g119(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n511), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n504), .A2(new_n505), .B1(new_n499), .B2(new_n500), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n547), .A2(G81), .B1(new_n501), .B2(G43), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  INV_X1    g129(.A(G65), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n555), .B1(new_n504), .B2(new_n505), .ZN(new_n556));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g133(.A(G651), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n547), .A2(G91), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n561), .B1(new_n501), .B2(G53), .ZN(new_n562));
  AND2_X1   g137(.A1(KEYINPUT6), .A2(G651), .ZN(new_n563));
  NOR2_X1   g138(.A1(KEYINPUT6), .A2(G651), .ZN(new_n564));
  OAI211_X1 g139(.A(G53), .B(G543), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n565), .A2(KEYINPUT9), .ZN(new_n566));
  OAI211_X1 g141(.A(new_n559), .B(new_n560), .C1(new_n562), .C2(new_n566), .ZN(G299));
  NOR2_X1   g142(.A1(new_n542), .A2(new_n543), .ZN(G301));
  INV_X1    g143(.A(G166), .ZN(G303));
  NAND2_X1  g144(.A1(new_n547), .A2(G87), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n501), .A2(G49), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(KEYINPUT75), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n570), .A2(new_n575), .A3(new_n571), .A4(new_n572), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(G288));
  NAND2_X1  g153(.A1(new_n547), .A2(G86), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT78), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n501), .A2(new_n582), .A3(G48), .ZN(new_n583));
  OAI211_X1 g158(.A(G48), .B(G543), .C1(new_n563), .C2(new_n564), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(KEYINPUT78), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n547), .A2(KEYINPUT77), .A3(G86), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n581), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AND2_X1   g163(.A1(G73), .A2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(G61), .B1(new_n532), .B2(new_n533), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n589), .B1(new_n590), .B2(KEYINPUT76), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT76), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n506), .A2(new_n592), .A3(G61), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n511), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G305));
  AOI22_X1  g171(.A1(new_n547), .A2(G85), .B1(new_n501), .B2(G47), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n511), .B2(new_n598), .ZN(G290));
  INV_X1    g174(.A(KEYINPUT79), .ZN(new_n600));
  AND3_X1   g175(.A1(new_n506), .A2(new_n507), .A3(G92), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT10), .ZN(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n534), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n605), .A2(G651), .B1(G54), .B2(new_n501), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n600), .B1(new_n608), .B2(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  MUX2_X1   g185(.A(new_n600), .B(new_n609), .S(new_n610), .Z(G284));
  MUX2_X1   g186(.A(new_n600), .B(new_n609), .S(new_n610), .Z(G321));
  XOR2_X1   g187(.A(G299), .B(KEYINPUT80), .Z(new_n613));
  MUX2_X1   g188(.A(new_n613), .B(G286), .S(G868), .Z(G280));
  XNOR2_X1  g189(.A(G280), .B(KEYINPUT81), .ZN(G297));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n608), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n608), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n479), .A2(new_n467), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  INV_X1    g199(.A(G2100), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n474), .A2(G123), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n459), .A2(G111), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  INV_X1    g205(.A(G135), .ZN(new_n631));
  OAI221_X1 g206(.A(new_n628), .B1(new_n629), .B2(new_n630), .C1(new_n631), .C2(new_n480), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(G2096), .Z(new_n633));
  NAND3_X1  g208(.A1(new_n626), .A2(new_n627), .A3(new_n633), .ZN(G156));
  XOR2_X1   g209(.A(G1341), .B(G1348), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT83), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2451), .B(G2454), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n636), .B(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT14), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT82), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2427), .B(G2430), .Z(new_n644));
  AOI21_X1  g219(.A(new_n640), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n644), .B2(new_n643), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n639), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(G14), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n647), .A2(new_n648), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(G401));
  XNOR2_X1  g227(.A(G2072), .B(G2078), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT85), .B(KEYINPUT17), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT84), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n657), .ZN(new_n661));
  OAI211_X1 g236(.A(new_n658), .B(new_n660), .C1(new_n661), .C2(new_n653), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT86), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n659), .A2(new_n656), .A3(new_n653), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT18), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n661), .A2(new_n660), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n665), .B1(new_n666), .B2(new_n655), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2096), .B(G2100), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G227));
  XOR2_X1   g245(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(G1986), .ZN(new_n673));
  XOR2_X1   g248(.A(G1956), .B(G2474), .Z(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n676), .A2(KEYINPUT87), .ZN(new_n677));
  XOR2_X1   g252(.A(G1971), .B(G1976), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(KEYINPUT87), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n677), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT20), .ZN(new_n682));
  INV_X1    g257(.A(G1981), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n674), .A2(new_n675), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(new_n676), .ZN(new_n685));
  MUX2_X1   g260(.A(new_n685), .B(new_n684), .S(new_n679), .Z(new_n686));
  NAND3_X1  g261(.A1(new_n682), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n683), .B1(new_n682), .B2(new_n686), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n673), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n689), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n691), .A2(G1986), .A3(new_n687), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n672), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G1991), .B(G1996), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT89), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT88), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n690), .A2(new_n692), .A3(new_n672), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n694), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n697), .ZN(new_n700));
  INV_X1    g275(.A(new_n698), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(new_n693), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(G229));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G32), .ZN(new_n706));
  AOI22_X1  g281(.A1(new_n481), .A2(G141), .B1(G129), .B2(new_n474), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT95), .B(KEYINPUT26), .ZN(new_n708));
  AND3_X1   g283(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  AOI22_X1  g286(.A1(new_n710), .A2(new_n711), .B1(G105), .B2(new_n467), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n707), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n706), .B1(new_n714), .B2(new_n705), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT96), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT27), .B(G1996), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G16), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G20), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT23), .ZN(new_n722));
  INV_X1    g297(.A(G299), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(new_n720), .ZN(new_n724));
  INV_X1    g299(.A(G1956), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n705), .A2(G26), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT28), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n474), .A2(G128), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT92), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n481), .A2(G140), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n459), .A2(G116), .ZN(new_n732));
  OAI21_X1  g307(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n730), .B(new_n731), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n728), .B1(new_n734), .B2(G29), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G2067), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n719), .A2(new_n726), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(G4), .A2(G16), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n608), .B2(G16), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT90), .B(G1348), .Z(new_n740));
  NOR2_X1   g315(.A1(G27), .A2(G29), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G164), .B2(G29), .ZN(new_n742));
  OAI22_X1  g317(.A1(new_n739), .A2(new_n740), .B1(G2078), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G2078), .B2(new_n742), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n720), .A2(G19), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n549), .B2(new_n720), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT91), .B(G1341), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(G168), .A2(new_n720), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n720), .B2(G21), .ZN(new_n751));
  INV_X1    g326(.A(G1966), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n749), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  AND2_X1   g328(.A1(KEYINPUT24), .A2(G34), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n705), .B1(KEYINPUT24), .B2(G34), .ZN(new_n755));
  OAI22_X1  g330(.A1(G160), .A2(new_n705), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI22_X1  g331(.A1(new_n746), .A2(new_n748), .B1(G2084), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n739), .A2(new_n740), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT30), .B(G28), .ZN(new_n760));
  OR2_X1    g335(.A1(KEYINPUT31), .A2(G11), .ZN(new_n761));
  NAND2_X1  g336(.A1(KEYINPUT31), .A2(G11), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n760), .A2(new_n705), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n632), .B2(new_n705), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n751), .B2(new_n752), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n744), .A2(new_n758), .A3(new_n759), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n705), .A2(G35), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G162), .B2(new_n705), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  AOI211_X1 g345(.A(new_n737), .B(new_n766), .C1(G2090), .C2(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(G5), .A2(G16), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G171), .B2(G16), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT98), .Z(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(G1961), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(G1961), .ZN(new_n776));
  AND3_X1   g351(.A1(new_n771), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n595), .A2(G16), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G6), .B2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT32), .B(G1981), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n779), .A2(new_n781), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n720), .A2(G22), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G166), .B2(new_n720), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(G1971), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n720), .A2(G23), .ZN(new_n787));
  INV_X1    g362(.A(new_n573), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(new_n720), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT33), .B(G1976), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n782), .A2(new_n783), .A3(new_n786), .A4(new_n791), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(KEYINPUT34), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(KEYINPUT34), .ZN(new_n794));
  MUX2_X1   g369(.A(G24), .B(G290), .S(G16), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(new_n673), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n705), .A2(G25), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n481), .A2(G131), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n474), .A2(G119), .ZN(new_n799));
  OR2_X1    g374(.A1(G95), .A2(G2105), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n800), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n798), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n797), .B1(new_n803), .B2(new_n705), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT35), .B(G1991), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n793), .A2(new_n794), .A3(new_n796), .A4(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT36), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n770), .A2(G2090), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT100), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n705), .A2(G33), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT93), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT25), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT94), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n479), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n816), .A2(new_n459), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n814), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n815), .ZN(new_n819));
  INV_X1    g394(.A(G139), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n820), .B2(new_n480), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n811), .B1(new_n822), .B2(new_n705), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(G2072), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n756), .A2(G2084), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n824), .B(new_n825), .C1(new_n718), .C2(new_n716), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT97), .Z(new_n827));
  NAND4_X1  g402(.A1(new_n777), .A2(new_n808), .A3(new_n810), .A4(new_n827), .ZN(G150));
  INV_X1    g403(.A(G150), .ZN(G311));
  NAND2_X1  g404(.A1(new_n501), .A2(G55), .ZN(new_n830));
  INV_X1    g405(.A(G93), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n831), .B2(new_n508), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n833), .A2(new_n511), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(G860), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT37), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n607), .A2(new_n616), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n549), .B(new_n835), .Z(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n844), .A2(KEYINPUT39), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n836), .B1(new_n844), .B2(KEYINPUT39), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n838), .B1(new_n845), .B2(new_n846), .ZN(G145));
  NAND2_X1  g422(.A1(new_n822), .A2(new_n714), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n713), .B1(new_n818), .B2(new_n821), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n848), .A2(new_n802), .A3(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n734), .B(G164), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n802), .B1(new_n848), .B2(new_n849), .ZN(new_n854));
  OR3_X1    g429(.A1(new_n851), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n853), .B1(new_n851), .B2(new_n854), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n474), .A2(G130), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n459), .A2(G118), .ZN(new_n859));
  OAI21_X1  g434(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n860));
  INV_X1    g435(.A(G142), .ZN(new_n861));
  OAI221_X1 g436(.A(new_n858), .B1(new_n859), .B2(new_n860), .C1(new_n861), .C2(new_n480), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n623), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n857), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT102), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n855), .A2(new_n863), .A3(new_n856), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n632), .B(G160), .Z(new_n869));
  XNOR2_X1  g444(.A(G162), .B(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(G37), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n865), .A2(new_n866), .A3(new_n867), .A4(new_n870), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g451(.A(G166), .B(KEYINPUT103), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n877), .A2(new_n595), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n595), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(G290), .B(new_n573), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT42), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n886));
  INV_X1    g461(.A(new_n884), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n881), .B1(new_n878), .B2(new_n879), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n883), .A2(KEYINPUT104), .A3(new_n884), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n885), .B1(new_n891), .B2(KEYINPUT42), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n607), .B(new_n723), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT41), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n842), .B(new_n618), .ZN(new_n896));
  MUX2_X1   g471(.A(new_n893), .B(new_n895), .S(new_n896), .Z(new_n897));
  XOR2_X1   g472(.A(new_n892), .B(new_n897), .Z(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(G868), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n899), .B1(G868), .B2(new_n835), .ZN(G295));
  OAI21_X1  g475(.A(new_n899), .B1(G868), .B2(new_n835), .ZN(G331));
  INV_X1    g476(.A(new_n842), .ZN(new_n902));
  NAND2_X1  g477(.A1(G301), .A2(G286), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(G301), .A2(G286), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n902), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(G171), .A2(G168), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n907), .A2(new_n842), .A3(new_n903), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n895), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n906), .A2(new_n893), .A3(new_n908), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n910), .A2(new_n890), .A3(new_n889), .A4(new_n911), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n906), .A2(new_n893), .A3(new_n908), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n894), .B1(new_n906), .B2(new_n908), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n891), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n912), .A2(new_n915), .A3(new_n873), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n916), .A2(KEYINPUT106), .A3(KEYINPUT43), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n912), .A2(new_n915), .A3(new_n921), .A4(new_n873), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n919), .A2(KEYINPUT44), .A3(new_n920), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n917), .A2(new_n922), .ZN(new_n924));
  XOR2_X1   g499(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(G397));
  INV_X1    g502(.A(KEYINPUT49), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n582), .B1(new_n501), .B2(G48), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n584), .A2(KEYINPUT78), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n579), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT113), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n594), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI22_X1  g508(.A1(new_n583), .A2(new_n585), .B1(G86), .B2(new_n547), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT113), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n683), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n588), .A2(G1981), .A3(new_n594), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n928), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n591), .A2(new_n593), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(G651), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n940), .B1(new_n934), .B2(KEYINPUT113), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n931), .A2(new_n932), .ZN(new_n942));
  OAI21_X1  g517(.A(G1981), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n581), .A2(new_n587), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n944), .A2(new_n683), .A3(new_n940), .A4(new_n586), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n943), .A2(KEYINPUT49), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G40), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n464), .A2(new_n469), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G1384), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n496), .A3(new_n949), .ZN(new_n950));
  XOR2_X1   g525(.A(KEYINPUT111), .B(G8), .Z(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT112), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n950), .A2(new_n955), .A3(new_n952), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n938), .A2(new_n946), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n788), .A2(G1976), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n950), .A2(new_n955), .A3(new_n952), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n955), .B1(new_n950), .B2(new_n952), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT52), .ZN(new_n963));
  INV_X1    g538(.A(G1976), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT52), .B1(G288), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n957), .A2(new_n959), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n958), .A2(new_n963), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(G8), .B1(new_n509), .B2(new_n512), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT55), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n968), .B(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n496), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n948), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT50), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n974), .B1(new_n496), .B2(new_n949), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n973), .A2(G2090), .A3(new_n975), .ZN(new_n976));
  XOR2_X1   g551(.A(KEYINPUT109), .B(G1971), .Z(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n496), .A2(new_n949), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n465), .A2(new_n468), .ZN(new_n982));
  INV_X1    g557(.A(G125), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n983), .B1(new_n472), .B2(new_n473), .ZN(new_n984));
  INV_X1    g559(.A(new_n463), .ZN(new_n985));
  OAI21_X1  g560(.A(G2105), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n982), .A2(new_n986), .A3(G40), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n980), .A2(G1384), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n987), .B1(new_n496), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n978), .B1(new_n981), .B2(new_n989), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n970), .B(G8), .C1(new_n976), .C2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n496), .A2(new_n988), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n948), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT45), .B1(new_n496), .B2(new_n949), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n979), .A2(KEYINPUT50), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n987), .B1(new_n496), .B2(new_n971), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI22_X1  g575(.A1(new_n997), .A2(new_n978), .B1(new_n1000), .B2(G2090), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n1001), .A2(KEYINPUT110), .A3(G8), .A4(new_n970), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n967), .B1(new_n993), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n970), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1001), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1004), .B1(new_n1005), .B2(new_n951), .ZN(new_n1006));
  INV_X1    g581(.A(G1961), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(new_n973), .B2(new_n975), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1009), .A2(G2078), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n981), .A2(new_n989), .A3(new_n1010), .ZN(new_n1011));
  NOR3_X1   g586(.A1(new_n995), .A2(G2078), .A3(new_n996), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1008), .B(new_n1011), .C1(new_n1012), .C2(KEYINPUT53), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(G171), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1003), .A2(new_n1006), .A3(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n752), .B1(new_n995), .B2(new_n996), .ZN(new_n1017));
  INV_X1    g592(.A(G2084), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n998), .A2(new_n1018), .A3(new_n999), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n952), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n1022));
  NAND2_X1  g597(.A1(G286), .A2(new_n952), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G8), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT121), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n1023), .B(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT51), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1024), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1023), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n1031), .B(KEYINPUT120), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT62), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1030), .A2(new_n1032), .A3(KEYINPUT62), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1016), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n958), .A2(new_n963), .A3(new_n966), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n993), .A2(new_n1002), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1021), .A2(G286), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n1006), .A4(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT63), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n970), .B1(new_n1001), .B2(G8), .ZN(new_n1043));
  NOR4_X1   g618(.A1(new_n1043), .A2(new_n1042), .A3(new_n1021), .A4(G286), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n1041), .A2(new_n1042), .B1(new_n1003), .B2(new_n1044), .ZN(new_n1045));
  AOI211_X1 g620(.A(G1976), .B(G288), .C1(new_n938), .C2(new_n946), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n957), .B1(new_n1046), .B2(new_n937), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1047), .B1(new_n1039), .B2(new_n967), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n1037), .A2(new_n1045), .A3(new_n1048), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1038), .A2(new_n1039), .A3(new_n1006), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n981), .A2(new_n989), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1009), .B1(new_n1051), .B2(G2078), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT45), .B1(new_n979), .B2(KEYINPUT107), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT107), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n496), .A2(new_n1054), .A3(new_n949), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n462), .A2(new_n463), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT122), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n459), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1059), .B1(new_n1058), .B2(new_n1057), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1009), .A2(new_n947), .A3(G2078), .ZN(new_n1061));
  AND4_X1   g636(.A1(new_n982), .A2(new_n994), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1056), .A2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(G301), .A2(new_n1052), .A3(new_n1063), .A4(new_n1008), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1014), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1030), .A2(new_n1032), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1052), .A2(new_n1063), .A3(new_n1008), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(G171), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT123), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1068), .A2(KEYINPUT123), .A3(G171), .ZN(new_n1072));
  OR2_X1    g647(.A1(new_n1013), .A2(G171), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1071), .A2(KEYINPUT54), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1050), .A2(new_n1067), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT124), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1050), .A2(new_n1067), .A3(new_n1074), .A4(KEYINPUT124), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n725), .B1(new_n973), .B2(new_n975), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n557), .B1(new_n534), .B2(new_n555), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1082), .A2(G651), .B1(new_n547), .B2(G91), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n501), .A2(new_n561), .A3(G53), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n565), .A2(KEYINPUT9), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI211_X1 g661(.A(KEYINPUT114), .B(new_n1081), .C1(new_n1083), .C2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT114), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT57), .B1(G299), .B2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT56), .B(G2072), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n981), .A2(new_n989), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1080), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1080), .A2(KEYINPUT115), .A3(new_n1092), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT115), .B1(new_n1080), .B2(new_n1092), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n1095), .A2(new_n1096), .A3(new_n1090), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n950), .A2(G2067), .ZN(new_n1099));
  INV_X1    g674(.A(G1348), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1099), .B1(new_n1000), .B2(new_n1100), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n1101), .A2(new_n607), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1094), .B1(new_n1098), .B2(new_n1102), .ZN(new_n1103));
  XOR2_X1   g678(.A(KEYINPUT58), .B(G1341), .Z(new_n1104));
  NAND2_X1  g679(.A1(new_n950), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n1051), .B2(G1996), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n549), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT59), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1107), .B(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT117), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1093), .A2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1080), .A2(new_n1090), .A3(new_n1092), .A4(KEYINPUT117), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT61), .B1(new_n1097), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1090), .B1(new_n1080), .B2(new_n1092), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT61), .B1(new_n1115), .B2(KEYINPUT116), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1093), .A2(KEYINPUT116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1116), .B1(new_n1117), .B2(new_n1115), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1109), .B1(new_n1114), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1101), .A2(KEYINPUT60), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(KEYINPUT118), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1101), .A2(new_n1122), .A3(KEYINPUT60), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1121), .A2(new_n608), .A3(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1120), .A2(KEYINPUT118), .A3(new_n607), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1124), .B(new_n1125), .C1(KEYINPUT60), .C2(new_n1101), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1103), .B1(new_n1119), .B2(new_n1126), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1077), .B(new_n1078), .C1(new_n1079), .C2(new_n1127), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1127), .A2(new_n1079), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1049), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1056), .A2(new_n987), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n713), .A2(G1996), .ZN(new_n1133));
  OR3_X1    g708(.A1(new_n1132), .A2(KEYINPUT108), .A3(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(KEYINPUT108), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n734), .B(G2067), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n713), .A2(G1996), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1134), .A2(new_n1135), .B1(new_n1131), .B2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n803), .A2(new_n805), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n803), .A2(new_n805), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1131), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g718(.A(G290), .B(G1986), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1143), .B1(new_n1131), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1130), .A2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1132), .A2(G1996), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(KEYINPUT46), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1131), .B1(new_n1136), .B2(new_n713), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n1149), .B(KEYINPUT126), .ZN(new_n1150));
  OR3_X1    g725(.A1(new_n1148), .A2(new_n1150), .A3(KEYINPUT47), .ZN(new_n1151));
  OAI21_X1  g726(.A(KEYINPUT47), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1143), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1132), .A2(G1986), .A3(G290), .ZN(new_n1154));
  XOR2_X1   g729(.A(new_n1154), .B(KEYINPUT48), .Z(new_n1155));
  AOI22_X1  g730(.A1(new_n1151), .A2(new_n1152), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n734), .A2(G2067), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1157), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1158));
  OR3_X1    g733(.A1(new_n1158), .A2(KEYINPUT125), .A3(new_n1132), .ZN(new_n1159));
  OAI21_X1  g734(.A(KEYINPUT125), .B1(new_n1158), .B2(new_n1132), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1156), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1146), .A2(new_n1161), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g737(.A(KEYINPUT127), .ZN(new_n1164));
  OAI21_X1  g738(.A(G319), .B1(new_n650), .B2(new_n651), .ZN(new_n1165));
  NOR2_X1   g739(.A1(G227), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g740(.A(new_n1164), .B1(new_n703), .B2(new_n1166), .ZN(new_n1167));
  AND3_X1   g741(.A1(new_n703), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1168));
  OAI211_X1 g742(.A(new_n924), .B(new_n875), .C1(new_n1167), .C2(new_n1168), .ZN(G225));
  INV_X1    g743(.A(G225), .ZN(G308));
endmodule


