//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 1 0 0 1 1 0 0 0 1 0 1 1 0 0 1 0 1 1 1 0 1 1 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n548, new_n549, new_n551, new_n552,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT67), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n458), .A2(G2105), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G101), .ZN(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G137), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n461), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(KEYINPUT68), .B1(new_n466), .B2(new_n462), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n468), .A2(new_n470), .A3(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n462), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n465), .B1(new_n467), .B2(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n468), .A2(new_n470), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(new_n462), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT69), .ZN(new_n480));
  NOR2_X1   g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT70), .Z(new_n482));
  INV_X1    g057(.A(G112), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n458), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n477), .A2(G2105), .ZN(new_n485));
  AOI22_X1  g060(.A1(new_n482), .A2(new_n484), .B1(new_n485), .B2(G136), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n480), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT71), .ZN(G162));
  NAND4_X1  g063(.A1(new_n468), .A2(new_n470), .A3(G126), .A4(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n468), .A2(new_n470), .A3(G138), .A4(new_n462), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n461), .A2(new_n496), .A3(G138), .A4(new_n462), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n493), .B1(new_n495), .B2(new_n497), .ZN(G164));
  XNOR2_X1  g073(.A(KEYINPUT5), .B(G543), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n499), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g077(.A(new_n502), .B(KEYINPUT73), .ZN(new_n503));
  OR2_X1    g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n506), .A2(new_n499), .ZN(new_n507));
  XOR2_X1   g082(.A(KEYINPUT72), .B(G88), .Z(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n509), .B1(new_n504), .B2(new_n505), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n507), .A2(new_n508), .B1(G50), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n503), .A2(new_n511), .ZN(G303));
  INV_X1    g087(.A(G303), .ZN(G166));
  NAND3_X1  g088(.A1(new_n499), .A2(G63), .A3(G651), .ZN(new_n514));
  INV_X1    g089(.A(new_n510), .ZN(new_n515));
  INV_X1    g090(.A(G51), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT74), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT74), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n514), .B(new_n519), .C1(new_n515), .C2(new_n516), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n507), .A2(G89), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n518), .A2(new_n520), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT75), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n523), .A2(new_n522), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n527), .A2(KEYINPUT75), .A3(new_n518), .A4(new_n520), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(new_n528), .ZN(G168));
  NAND2_X1  g104(.A1(new_n510), .A2(G52), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n506), .A2(new_n499), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n499), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n535), .A2(new_n536), .B1(new_n501), .B2(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  AOI22_X1  g114(.A1(new_n499), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n501), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n510), .A2(G43), .ZN(new_n543));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n544), .B2(new_n532), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT77), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n548), .A2(new_n552), .ZN(G188));
  NAND2_X1  g128(.A1(new_n510), .A2(G53), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT78), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(KEYINPUT9), .ZN(new_n556));
  MUX2_X1   g131(.A(KEYINPUT9), .B(new_n556), .S(KEYINPUT79), .Z(new_n557));
  NOR2_X1   g132(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n510), .A2(G53), .B1(new_n555), .B2(KEYINPUT9), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n499), .A2(G65), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n563), .A2(G651), .B1(new_n507), .B2(G91), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n560), .A2(new_n564), .ZN(G299));
  INV_X1    g140(.A(G168), .ZN(G286));
  NAND2_X1  g141(.A1(new_n510), .A2(G49), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT80), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n499), .A2(G74), .ZN(new_n569));
  AOI22_X1  g144(.A1(G651), .A2(new_n569), .B1(new_n507), .B2(G87), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(G288));
  AOI22_X1  g146(.A1(new_n507), .A2(G86), .B1(G48), .B2(new_n510), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n499), .A2(G61), .ZN(new_n573));
  NAND2_X1  g148(.A1(G73), .A2(G543), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n501), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(KEYINPUT81), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT81), .ZN(new_n577));
  AOI211_X1 g152(.A(new_n577), .B(new_n501), .C1(new_n573), .C2(new_n574), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n572), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT82), .ZN(G305));
  NAND2_X1  g155(.A1(new_n510), .A2(G47), .ZN(new_n581));
  INV_X1    g156(.A(G85), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n582), .B2(new_n532), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n499), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n501), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  XOR2_X1   g163(.A(new_n588), .B(KEYINPUT83), .Z(new_n589));
  XNOR2_X1  g164(.A(KEYINPUT84), .B(KEYINPUT10), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n507), .A2(G92), .A3(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n590), .ZN(new_n592));
  INV_X1    g167(.A(G92), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n532), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n591), .A2(new_n594), .B1(G54), .B2(new_n510), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT85), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(G66), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(G66), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n499), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT86), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n599), .A2(KEYINPUT86), .A3(new_n600), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n603), .A2(G651), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n595), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(KEYINPUT87), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT87), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n595), .A2(new_n605), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n589), .B1(G868), .B2(new_n610), .ZN(G284));
  OAI21_X1  g186(.A(new_n589), .B1(G868), .B2(new_n610), .ZN(G321));
  NOR2_X1   g187(.A1(G299), .A2(G868), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g189(.A(new_n613), .B1(G168), .B2(G868), .ZN(G280));
  XNOR2_X1  g190(.A(KEYINPUT88), .B(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n610), .B1(G860), .B2(new_n616), .ZN(G148));
  INV_X1    g192(.A(new_n546), .ZN(new_n618));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AND2_X1   g195(.A1(new_n610), .A2(new_n616), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n619), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g198(.A1(new_n463), .A2(new_n458), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT89), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  INV_X1    g202(.A(G2100), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n485), .A2(G135), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n478), .A2(G123), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n462), .A2(G111), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n631), .B(new_n632), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2096), .Z(new_n636));
  NAND3_X1  g211(.A1(new_n629), .A2(new_n630), .A3(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(KEYINPUT14), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT90), .B(KEYINPUT16), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2451), .B(G2454), .Z(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n645), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(KEYINPUT91), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n649), .A2(new_n650), .ZN(new_n654));
  INV_X1    g229(.A(G14), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G401));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT92), .Z(new_n660));
  XNOR2_X1  g235(.A(G2072), .B(G2078), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n661), .B(KEYINPUT17), .Z(new_n666));
  OAI211_X1 g241(.A(new_n663), .B(new_n665), .C1(new_n660), .C2(new_n666), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n664), .A2(new_n659), .A3(new_n661), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT18), .Z(new_n669));
  NAND3_X1  g244(.A1(new_n660), .A2(new_n666), .A3(new_n664), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n667), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(new_n628), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT93), .B(G2096), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT19), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n680), .A2(new_n681), .ZN(new_n684));
  NOR3_X1   g259(.A1(new_n679), .A2(new_n684), .A3(new_n682), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n679), .A2(new_n684), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT94), .B(KEYINPUT20), .Z(new_n687));
  AOI211_X1 g262(.A(new_n683), .B(new_n685), .C1(new_n686), .C2(new_n687), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(new_n686), .B2(new_n687), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n689), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1991), .B(G1996), .Z(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n692), .A2(new_n693), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n676), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n692), .A2(new_n693), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n698), .A2(new_n675), .A3(new_n694), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(G229));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n702), .A2(G33), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT25), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G139), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(new_n463), .ZN(new_n708));
  NAND2_X1  g283(.A1(G115), .A2(G2104), .ZN(new_n709));
  INV_X1    g284(.A(G127), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n477), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n708), .B1(G2105), .B2(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT97), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n703), .B1(new_n713), .B2(G29), .ZN(new_n714));
  INV_X1    g289(.A(G2072), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT24), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n702), .B1(new_n716), .B2(G34), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(KEYINPUT98), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(KEYINPUT98), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n716), .B2(G34), .ZN(new_n720));
  AOI22_X1  g295(.A1(G160), .A2(G29), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  OAI22_X1  g296(.A1(new_n714), .A2(new_n715), .B1(G2084), .B2(new_n721), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n714), .A2(new_n715), .ZN(new_n723));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G20), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT23), .Z(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G299), .B2(G16), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(G1956), .Z(new_n728));
  OR3_X1    g303(.A1(new_n722), .A2(new_n723), .A3(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(G29), .A2(G35), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G162), .B2(G29), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT29), .B(G2090), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n702), .A2(G32), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n485), .A2(G141), .B1(G105), .B2(new_n459), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n478), .A2(G129), .ZN(new_n736));
  NAND3_X1  g311(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT26), .Z(new_n738));
  AND3_X1   g313(.A1(new_n735), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n734), .B1(new_n739), .B2(new_n702), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT27), .B(G1996), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n740), .A2(new_n742), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT30), .B(G28), .ZN(new_n745));
  OR2_X1    g320(.A1(KEYINPUT31), .A2(G11), .ZN(new_n746));
  NAND2_X1  g321(.A1(KEYINPUT31), .A2(G11), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n745), .A2(new_n702), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n635), .B2(new_n702), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n744), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(G27), .A2(G29), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G164), .B2(G29), .ZN(new_n752));
  INV_X1    g327(.A(G2078), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n733), .A2(new_n743), .A3(new_n750), .A4(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n731), .A2(new_n732), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n721), .A2(G2084), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT99), .ZN(new_n758));
  NOR4_X1   g333(.A1(new_n729), .A2(new_n755), .A3(new_n756), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n724), .A2(G21), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G168), .B2(new_n724), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G1966), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT100), .Z(new_n763));
  OR2_X1    g338(.A1(new_n761), .A2(G1966), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n724), .A2(G5), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G171), .B2(new_n724), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT101), .ZN(new_n767));
  INV_X1    g342(.A(G1961), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n759), .A2(new_n763), .A3(new_n764), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n724), .A2(G19), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n546), .B2(new_n724), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(G1341), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n702), .A2(G26), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT28), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n485), .A2(G140), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n478), .A2(G128), .ZN(new_n777));
  OR2_X1    g352(.A1(G104), .A2(G2105), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n778), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n775), .B1(new_n781), .B2(new_n702), .ZN(new_n782));
  INV_X1    g357(.A(G2067), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n724), .A2(G4), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n610), .B2(new_n724), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n773), .B(new_n784), .C1(G1348), .C2(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G1348), .B2(new_n786), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT96), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n770), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT36), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n724), .A2(G23), .ZN(new_n793));
  INV_X1    g368(.A(G288), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(new_n724), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT33), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G1976), .ZN(new_n797));
  NOR2_X1   g372(.A1(G16), .A2(G22), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G166), .B2(G16), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(G1971), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(G6), .A2(G16), .ZN(new_n802));
  INV_X1    g377(.A(G305), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(G16), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT32), .B(G1981), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NOR3_X1   g381(.A1(new_n801), .A2(KEYINPUT34), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n724), .A2(G24), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n586), .B2(new_n724), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G1986), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n702), .A2(G25), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n478), .A2(G119), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT95), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n462), .A2(G107), .ZN(new_n814));
  OAI21_X1  g389(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n485), .A2(G131), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n811), .B1(new_n819), .B2(new_n702), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT35), .B(G1991), .Z(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n820), .B(new_n822), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n807), .A2(new_n810), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(KEYINPUT34), .B1(new_n801), .B2(new_n806), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n792), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n824), .A2(new_n792), .A3(new_n825), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n791), .B1(new_n827), .B2(new_n828), .ZN(G311));
  INV_X1    g404(.A(new_n828), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n790), .B1(new_n830), .B2(new_n826), .ZN(G150));
  AOI22_X1  g406(.A1(new_n507), .A2(G93), .B1(G55), .B2(new_n510), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n499), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n501), .B2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT102), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(G860), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT37), .Z(new_n837));
  NOR2_X1   g412(.A1(new_n618), .A2(new_n834), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(new_n835), .B2(new_n618), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT38), .Z(new_n840));
  NAND2_X1  g415(.A1(new_n610), .A2(G559), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT39), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(G860), .B1(new_n842), .B2(new_n843), .ZN(new_n845));
  AND3_X1   g420(.A1(new_n844), .A2(KEYINPUT103), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(KEYINPUT103), .B1(new_n844), .B2(new_n845), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n837), .B1(new_n846), .B2(new_n847), .ZN(G145));
  XNOR2_X1  g423(.A(G162), .B(new_n635), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(G160), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n713), .B(new_n739), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n485), .A2(G142), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n478), .A2(G130), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n462), .A2(G118), .ZN(new_n854));
  OAI21_X1  g429(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n852), .B(new_n853), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT104), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(new_n626), .Z(new_n858));
  OR2_X1    g433(.A1(new_n851), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n495), .A2(new_n497), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n489), .A2(new_n492), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n780), .B(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n818), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n851), .A2(new_n858), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n859), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n864), .B1(new_n859), .B2(new_n865), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n850), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  INV_X1    g445(.A(G160), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n849), .B(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n872), .A3(new_n866), .ZN(new_n873));
  INV_X1    g448(.A(G37), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n869), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(KEYINPUT40), .Z(G395));
  INV_X1    g451(.A(KEYINPUT105), .ZN(new_n877));
  NAND2_X1  g452(.A1(G299), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n560), .A2(new_n564), .A3(KEYINPUT105), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n878), .A2(new_n605), .A3(new_n595), .A4(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n606), .A2(new_n877), .A3(G299), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n882), .A2(KEYINPUT41), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(KEYINPUT41), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n883), .A2(KEYINPUT106), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT106), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n882), .A2(new_n886), .A3(KEYINPUT41), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n621), .B(new_n839), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n882), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n803), .A2(new_n586), .ZN(new_n893));
  NAND2_X1  g468(.A1(G305), .A2(G290), .ZN(new_n894));
  XNOR2_X1  g469(.A(G303), .B(G288), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n895), .B1(new_n893), .B2(new_n894), .ZN(new_n897));
  OAI21_X1  g472(.A(KEYINPUT42), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OR3_X1    g473(.A1(new_n896), .A2(new_n897), .A3(KEYINPUT42), .ZN(new_n899));
  AND4_X1   g474(.A1(new_n890), .A2(new_n892), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  AOI22_X1  g475(.A1(new_n890), .A2(new_n892), .B1(new_n899), .B2(new_n898), .ZN(new_n901));
  OAI21_X1  g476(.A(G868), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT107), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n835), .A2(new_n619), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n903), .B1(new_n902), .B2(new_n904), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(G295));
  NAND2_X1  g482(.A1(new_n902), .A2(new_n904), .ZN(G331));
  INV_X1    g483(.A(KEYINPUT108), .ZN(new_n909));
  XNOR2_X1  g484(.A(G168), .B(G171), .ZN(new_n910));
  INV_X1    g485(.A(new_n839), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(G168), .B(G301), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n839), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(new_n887), .A3(new_n885), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n896), .A2(new_n897), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n912), .A2(new_n914), .A3(new_n891), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n874), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n917), .B1(new_n916), .B2(new_n918), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n909), .B(KEYINPUT43), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT43), .ZN(new_n923));
  INV_X1    g498(.A(new_n920), .ZN(new_n924));
  INV_X1    g499(.A(new_n921), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n918), .ZN(new_n927));
  AOI22_X1  g502(.A1(new_n912), .A2(new_n914), .B1(new_n884), .B2(new_n883), .ZN(new_n928));
  OAI22_X1  g503(.A1(new_n927), .A2(new_n928), .B1(new_n896), .B2(new_n897), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n929), .A2(new_n919), .A3(new_n874), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT108), .B1(new_n930), .B2(KEYINPUT43), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n922), .B1(new_n926), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n924), .A2(new_n923), .A3(new_n925), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(KEYINPUT109), .A3(KEYINPUT43), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(new_n934), .A3(KEYINPUT44), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT109), .B1(new_n930), .B2(KEYINPUT43), .ZN(new_n936));
  OAI22_X1  g511(.A1(new_n932), .A2(KEYINPUT44), .B1(new_n935), .B2(new_n936), .ZN(G397));
  INV_X1    g512(.A(KEYINPUT45), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(G164), .B2(G1384), .ZN(new_n939));
  AOI22_X1  g514(.A1(new_n485), .A2(G137), .B1(G101), .B2(new_n459), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n471), .A2(new_n472), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n474), .B1(new_n941), .B2(G2105), .ZN(new_n942));
  AOI211_X1 g517(.A(KEYINPUT68), .B(new_n462), .C1(new_n471), .C2(new_n472), .ZN(new_n943));
  OAI211_X1 g518(.A(G40), .B(new_n940), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n939), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(G1986), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(new_n946), .A3(new_n586), .ZN(new_n947));
  XNOR2_X1  g522(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n947), .A2(new_n948), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n819), .A2(new_n821), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n780), .B(new_n783), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n739), .B(G1996), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n818), .A2(new_n822), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n951), .A2(new_n952), .A3(new_n953), .A4(new_n954), .ZN(new_n955));
  AOI211_X1 g530(.A(new_n949), .B(new_n950), .C1(new_n945), .C2(new_n955), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n939), .A2(new_n944), .A3(G1996), .ZN(new_n957));
  OR2_X1    g532(.A1(new_n957), .A2(KEYINPUT46), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n952), .A2(new_n739), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n945), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n957), .A2(KEYINPUT46), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n962), .B(KEYINPUT125), .ZN(new_n963));
  XOR2_X1   g538(.A(new_n963), .B(KEYINPUT47), .Z(new_n964));
  NAND2_X1  g539(.A1(new_n953), .A2(new_n952), .ZN(new_n965));
  OAI22_X1  g540(.A1(new_n965), .A2(new_n951), .B1(G2067), .B2(new_n780), .ZN(new_n966));
  AOI211_X1 g541(.A(new_n956), .B(new_n964), .C1(new_n945), .C2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT123), .ZN(new_n968));
  INV_X1    g543(.A(new_n944), .ZN(new_n969));
  INV_X1    g544(.A(G2084), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n971));
  INV_X1    g546(.A(G1384), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n862), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n969), .A2(new_n970), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(G1384), .B1(new_n860), .B2(new_n861), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n976), .A2(KEYINPUT45), .ZN(new_n977));
  AOI211_X1 g552(.A(new_n938), .B(G1384), .C1(new_n860), .C2(new_n861), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n977), .A2(new_n978), .A3(new_n944), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n975), .B1(new_n979), .B2(G1966), .ZN(new_n980));
  OAI211_X1 g555(.A(KEYINPUT121), .B(G8), .C1(new_n980), .C2(G286), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT51), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G8), .ZN(new_n984));
  INV_X1    g559(.A(G1966), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n976), .A2(KEYINPUT45), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n939), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n985), .B1(new_n987), .B2(new_n944), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n984), .B1(new_n988), .B2(new_n975), .ZN(new_n989));
  NOR2_X1   g564(.A1(G168), .A2(new_n984), .ZN(new_n990));
  OAI211_X1 g565(.A(KEYINPUT121), .B(KEYINPUT51), .C1(new_n989), .C2(new_n990), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n983), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n980), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n968), .B(KEYINPUT62), .C1(new_n992), .C2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT110), .B1(new_n976), .B2(KEYINPUT45), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n997), .B(new_n938), .C1(G164), .C2(G1384), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n996), .A2(new_n969), .A3(new_n998), .A4(new_n986), .ZN(new_n999));
  XNOR2_X1  g574(.A(KEYINPUT111), .B(G1971), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT112), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n974), .A2(new_n973), .A3(G40), .A4(G160), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1002), .B1(new_n1003), .B2(G2090), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n862), .A2(new_n972), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n944), .B1(KEYINPUT50), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G2090), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1006), .A2(KEYINPUT112), .A3(new_n1007), .A4(new_n973), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1001), .A2(new_n1004), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n1011));
  AOI211_X1 g586(.A(new_n1011), .B(new_n984), .C1(new_n503), .C2(new_n511), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1009), .B(G8), .C1(new_n1010), .C2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n978), .A2(new_n944), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1014), .A2(new_n753), .A3(new_n998), .A4(new_n996), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n1016));
  AOI22_X1  g591(.A1(new_n1015), .A2(new_n1016), .B1(new_n768), .B2(new_n1003), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n979), .A2(KEYINPUT53), .A3(new_n753), .ZN(new_n1018));
  AOI21_X1  g593(.A(G301), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n944), .A2(new_n1005), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1020), .A2(new_n984), .ZN(new_n1021));
  INV_X1    g596(.A(G1976), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT52), .B1(G288), .B2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1021), .B(new_n1023), .C1(new_n1022), .C2(G288), .ZN(new_n1024));
  INV_X1    g599(.A(new_n572), .ZN(new_n1025));
  OAI21_X1  g600(.A(G1981), .B1(new_n1025), .B2(new_n575), .ZN(new_n1026));
  INV_X1    g601(.A(G1981), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1027), .B(new_n572), .C1(new_n576), .C2(new_n578), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT49), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1026), .A2(new_n1028), .A3(KEYINPUT49), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1031), .A2(new_n1021), .A3(new_n1032), .ZN(new_n1033));
  OAI221_X1 g608(.A(G8), .B1(new_n944), .B2(new_n1005), .C1(G288), .C2(new_n1022), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT52), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n1024), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1003), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1007), .A2(new_n1038), .B1(new_n999), .B2(new_n1000), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1037), .B1(new_n1039), .B2(new_n984), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1013), .A2(new_n1019), .A3(new_n1036), .A4(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n994), .B1(new_n983), .B2(new_n991), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT62), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1041), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT123), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n995), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1033), .A2(new_n1022), .A3(new_n794), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1028), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1021), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1036), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1049), .B1(new_n1013), .B2(new_n1050), .ZN(new_n1051));
  XOR2_X1   g626(.A(KEYINPUT114), .B(KEYINPUT63), .Z(new_n1052));
  NAND2_X1  g627(.A1(new_n989), .A2(G168), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT113), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n989), .A2(new_n1055), .A3(G168), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1013), .A2(new_n1036), .A3(new_n1040), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1052), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1013), .A2(new_n1036), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1009), .A2(G8), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n1037), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1061), .A2(new_n1057), .A3(KEYINPUT63), .A4(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1051), .B1(new_n1060), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G1348), .ZN(new_n1066));
  NAND4_X1  g641(.A1(G160), .A2(G40), .A3(new_n783), .A4(new_n976), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1003), .A2(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1020), .A2(KEYINPUT116), .A3(new_n783), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g646(.A(KEYINPUT56), .B(G2072), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1014), .A2(new_n998), .A3(new_n996), .A4(new_n1072), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT115), .B(G1956), .Z(new_n1074));
  NAND2_X1  g649(.A1(new_n1003), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n554), .A2(new_n556), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1076), .B1(new_n554), .B2(new_n557), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n499), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n1078));
  INV_X1    g653(.A(G91), .ZN(new_n1079));
  OAI22_X1  g654(.A1(new_n1078), .A2(new_n501), .B1(new_n532), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT57), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n560), .A2(new_n564), .A3(new_n1082), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1073), .A2(new_n1075), .A3(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1071), .A2(new_n1085), .A3(new_n610), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1081), .A2(new_n1083), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1088), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1087), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1086), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT118), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1086), .A2(new_n1095), .A3(new_n1092), .ZN(new_n1096));
  INV_X1    g671(.A(G1996), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1014), .A2(new_n1097), .A3(new_n998), .A4(new_n996), .ZN(new_n1098));
  XOR2_X1   g673(.A(KEYINPUT58), .B(G1341), .Z(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n944), .B2(new_n1005), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT59), .B1(new_n1101), .B2(new_n546), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n1103));
  AOI211_X1 g678(.A(new_n1103), .B(new_n618), .C1(new_n1098), .C2(new_n1100), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT61), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1106), .B1(new_n1087), .B2(new_n1091), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1085), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1073), .A2(new_n1075), .A3(new_n1084), .A4(KEYINPUT119), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1107), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1085), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1084), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1106), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1105), .A2(new_n1111), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT60), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1003), .A2(new_n1066), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1117), .A2(new_n1070), .A3(KEYINPUT60), .A4(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT120), .B1(new_n607), .B2(new_n609), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1069), .A2(new_n1120), .A3(KEYINPUT60), .A4(new_n1070), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n607), .A2(KEYINPUT120), .A3(new_n609), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1116), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1094), .B(new_n1096), .C1(new_n1115), .C2(new_n1126), .ZN(new_n1127));
  XOR2_X1   g702(.A(G301), .B(KEYINPUT54), .Z(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1003), .A2(new_n768), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1130), .A2(new_n1131), .A3(new_n1018), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n753), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1134));
  OR4_X1    g709(.A1(new_n465), .A2(new_n987), .A3(new_n473), .A4(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1017), .A2(new_n1128), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1042), .A2(new_n1059), .A3(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1127), .B1(new_n1138), .B2(KEYINPUT122), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n1140));
  NOR4_X1   g715(.A1(new_n1042), .A2(new_n1059), .A3(new_n1137), .A4(new_n1140), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1046), .B(new_n1065), .C1(new_n1139), .C2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n586), .B(new_n946), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n945), .B1(new_n955), .B2(new_n1143), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1142), .A2(KEYINPUT124), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT124), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n967), .B1(new_n1145), .B2(new_n1146), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g722(.A(G319), .ZN(new_n1149));
  OAI21_X1  g723(.A(KEYINPUT127), .B1(G227), .B2(new_n1149), .ZN(new_n1150));
  OR3_X1    g724(.A1(G227), .A2(KEYINPUT127), .A3(new_n1149), .ZN(new_n1151));
  NAND4_X1  g725(.A1(new_n700), .A2(new_n657), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  NOR2_X1   g726(.A1(new_n875), .A2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g727(.A(new_n1153), .B(new_n922), .C1(new_n926), .C2(new_n931), .ZN(G225));
  INV_X1    g728(.A(G225), .ZN(G308));
endmodule


