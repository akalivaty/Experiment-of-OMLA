//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 0 1 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1216, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G97), .A2(G257), .ZN(new_n207));
  INV_X1    g0007(.A(G87), .ZN(new_n208));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  OAI21_X1  g0009(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AOI21_X1  g0010(.A(new_n210), .B1(G68), .B2(G238), .ZN(new_n211));
  INV_X1    g0011(.A(G107), .ZN(new_n212));
  INV_X1    g0012(.A(G264), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n214), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G77), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G58), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n206), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT0), .Z(new_n228));
  INV_X1    g0028(.A(G68), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n221), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NOR3_X1   g0032(.A1(new_n231), .A2(new_n204), .A3(new_n232), .ZN(new_n233));
  NOR3_X1   g0033(.A1(new_n225), .A2(new_n228), .A3(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G264), .ZN(new_n240));
  INV_X1    g0040(.A(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n238), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT64), .ZN(new_n245));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(new_n212), .ZN(new_n249));
  INV_X1    g0049(.A(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n247), .B(new_n251), .ZN(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n232), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  OAI22_X1  g0056(.A1(new_n256), .A2(new_n216), .B1(new_n204), .B2(G68), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n204), .A2(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(new_n218), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n254), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(KEYINPUT11), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n254), .B1(new_n203), .B2(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G68), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n263), .B(KEYINPUT70), .ZN(new_n264));
  INV_X1    g0064(.A(G13), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G1), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(G20), .A3(new_n229), .ZN(new_n267));
  XNOR2_X1  g0067(.A(new_n267), .B(KEYINPUT12), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n261), .A2(new_n264), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G169), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT65), .B(G45), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n203), .B(G274), .C1(new_n272), .C2(G41), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT69), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n273), .B(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n232), .B1(G33), .B2(G41), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n222), .A2(G1698), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n277), .B1(G226), .B2(G1698), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT66), .ZN(new_n279));
  AND2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT3), .ZN(new_n283));
  INV_X1    g0083(.A(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(KEYINPUT66), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n278), .B1(new_n282), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G33), .A2(G97), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n276), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n232), .ZN(new_n292));
  INV_X1    g0092(.A(G41), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n292), .B1(new_n284), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G238), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n275), .A2(new_n291), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT13), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT13), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n275), .A2(new_n301), .A3(new_n291), .A4(new_n298), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n271), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT14), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n300), .A2(G179), .A3(new_n302), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT71), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n305), .B(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n270), .B1(new_n304), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n300), .A2(G190), .A3(new_n302), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n270), .ZN(new_n310));
  INV_X1    g0110(.A(G200), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(new_n300), .B2(new_n302), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(G20), .B1(new_n230), .B2(G50), .ZN(new_n315));
  INV_X1    g0115(.A(G150), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT8), .B(G58), .ZN(new_n317));
  OAI221_X1 g0117(.A(new_n315), .B1(new_n316), .B2(new_n256), .C1(new_n258), .C2(new_n317), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n318), .A2(new_n254), .B1(G50), .B2(new_n262), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n266), .A2(G20), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(G50), .B2(new_n320), .ZN(new_n321));
  XNOR2_X1  g0121(.A(new_n321), .B(KEYINPUT9), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n282), .A2(new_n287), .ZN(new_n323));
  INV_X1    g0123(.A(G1698), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G222), .ZN(new_n325));
  NAND2_X1  g0125(.A1(G223), .A2(G1698), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n323), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n327), .B(new_n276), .C1(G77), .C2(new_n323), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n328), .B(new_n273), .C1(new_n217), .C2(new_n296), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G200), .ZN(new_n330));
  INV_X1    g0130(.A(G190), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n322), .B(new_n330), .C1(new_n331), .C2(new_n329), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT10), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(new_n330), .B2(KEYINPUT68), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n332), .B(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n329), .A2(new_n271), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n336), .B(new_n321), .C1(G179), .C2(new_n329), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n320), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n317), .ZN(new_n340));
  INV_X1    g0140(.A(new_n262), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n340), .B1(new_n341), .B2(new_n317), .ZN(new_n342));
  XOR2_X1   g0142(.A(KEYINPUT72), .B(KEYINPUT7), .Z(new_n343));
  NOR2_X1   g0143(.A1(new_n280), .A2(new_n281), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n343), .A2(new_n204), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n285), .A2(new_n286), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT7), .B1(new_n346), .B2(G20), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n345), .A2(new_n347), .A3(G68), .ZN(new_n348));
  XNOR2_X1  g0148(.A(G58), .B(G68), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n349), .A2(G20), .B1(G159), .B2(new_n255), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n348), .A2(KEYINPUT16), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n254), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT7), .ZN(new_n354));
  NOR4_X1   g0154(.A1(new_n280), .A2(new_n281), .A3(new_n354), .A4(G20), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n282), .A2(new_n287), .A3(new_n204), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n355), .B1(new_n356), .B2(new_n343), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n350), .B1(new_n357), .B2(new_n229), .ZN(new_n358));
  XOR2_X1   g0158(.A(KEYINPUT73), .B(KEYINPUT16), .Z(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n342), .B1(new_n353), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n217), .A2(G1698), .ZN(new_n362));
  OAI221_X1 g0162(.A(new_n362), .B1(G223), .B2(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n363));
  NAND2_X1  g0163(.A1(G33), .A2(G87), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(KEYINPUT74), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT74), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n363), .A2(new_n367), .A3(new_n364), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n366), .A2(new_n276), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n297), .A2(G232), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n273), .ZN(new_n372));
  OAI21_X1  g0172(.A(G200), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n372), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n374), .A2(G190), .A3(new_n369), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n361), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT17), .ZN(new_n377));
  XNOR2_X1  g0177(.A(new_n376), .B(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT18), .ZN(new_n379));
  OAI21_X1  g0179(.A(G169), .B1(new_n370), .B2(new_n372), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n374), .A2(G179), .A3(new_n369), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n379), .B1(new_n382), .B2(new_n361), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n380), .A2(new_n381), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n352), .B1(new_n358), .B2(new_n359), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n384), .B(KEYINPUT18), .C1(new_n385), .C2(new_n342), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n378), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G238), .A2(G1698), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n323), .B(new_n389), .C1(new_n222), .C2(G1698), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n390), .B(new_n276), .C1(G107), .C2(new_n323), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n391), .B(new_n273), .C1(new_n219), .C2(new_n296), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n271), .ZN(new_n393));
  INV_X1    g0193(.A(new_n317), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n394), .A2(new_n255), .B1(G20), .B2(G77), .ZN(new_n395));
  XOR2_X1   g0195(.A(KEYINPUT15), .B(G87), .Z(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n395), .B1(new_n258), .B2(new_n397), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n398), .A2(new_n254), .B1(G77), .B2(new_n262), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n339), .A2(new_n218), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n393), .B(new_n401), .C1(G179), .C2(new_n392), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n392), .A2(G200), .ZN(new_n403));
  INV_X1    g0203(.A(new_n401), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n403), .B(new_n404), .C1(new_n331), .C2(new_n392), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  XOR2_X1   g0206(.A(new_n406), .B(KEYINPUT67), .Z(new_n407));
  AND4_X1   g0207(.A1(new_n314), .A2(new_n338), .A3(new_n388), .A4(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n356), .A2(new_n343), .ZN(new_n409));
  INV_X1    g0209(.A(new_n355), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT75), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n412), .A3(G107), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n212), .A2(KEYINPUT6), .A3(G97), .ZN(new_n414));
  XOR2_X1   g0214(.A(G97), .B(G107), .Z(new_n415));
  OAI21_X1  g0215(.A(new_n414), .B1(new_n415), .B2(KEYINPUT6), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n416), .A2(G20), .B1(G77), .B2(new_n255), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT75), .B1(new_n357), .B2(new_n212), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n413), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n254), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n324), .A2(G244), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT4), .ZN(new_n422));
  OAI22_X1  g0222(.A1(new_n421), .A2(new_n422), .B1(new_n209), .B2(new_n324), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n323), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n421), .B1(new_n285), .B2(new_n286), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT77), .B1(new_n425), .B2(KEYINPUT4), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G283), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT77), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n428), .B(new_n422), .C1(new_n344), .C2(new_n421), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n424), .A2(new_n426), .A3(new_n427), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n276), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT5), .B(G41), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n203), .A2(G45), .A3(G274), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n432), .A2(new_n203), .A3(G45), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n436), .A2(G257), .A3(new_n294), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n431), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(G200), .ZN(new_n440));
  INV_X1    g0240(.A(G97), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n320), .A2(new_n441), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n253), .A2(new_n232), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n203), .A2(G33), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(new_n320), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n442), .B1(new_n446), .B2(new_n441), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT76), .ZN(new_n448));
  OR2_X1    g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n448), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n437), .B1(new_n430), .B2(new_n276), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n452), .A2(G190), .A3(new_n435), .ZN(new_n453));
  AND4_X1   g0253(.A1(new_n420), .A2(new_n440), .A3(new_n451), .A4(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G179), .ZN(new_n455));
  AND4_X1   g0255(.A1(new_n455), .A2(new_n431), .A3(new_n435), .A4(new_n438), .ZN(new_n456));
  AOI21_X1  g0256(.A(G169), .B1(new_n452), .B2(new_n435), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n420), .A2(new_n451), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT78), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n419), .A2(new_n254), .B1(new_n449), .B2(new_n450), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n431), .A2(new_n455), .A3(new_n435), .A4(new_n438), .ZN(new_n463));
  INV_X1    g0263(.A(new_n435), .ZN(new_n464));
  AOI211_X1 g0264(.A(new_n464), .B(new_n437), .C1(new_n430), .C2(new_n276), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n463), .B1(new_n465), .B2(G169), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT78), .B1(new_n462), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n454), .B1(new_n461), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n282), .A2(new_n287), .A3(G303), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n213), .A2(G1698), .ZN(new_n470));
  OAI221_X1 g0270(.A(new_n470), .B1(G257), .B2(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT81), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT81), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n469), .A2(new_n474), .A3(new_n471), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n473), .A2(new_n276), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n436), .A2(new_n294), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n435), .B1(new_n477), .B2(new_n241), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n446), .A2(G116), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n339), .A2(new_n250), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n253), .A2(new_n232), .B1(G20), .B2(new_n250), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n427), .B(new_n204), .C1(G33), .C2(new_n441), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT20), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n483), .A2(KEYINPUT20), .A3(new_n484), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n481), .B(new_n482), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n480), .A2(new_n488), .A3(new_n455), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n469), .A2(new_n474), .A3(new_n471), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n474), .B1(new_n469), .B2(new_n471), .ZN(new_n491));
  NOR3_X1   g0291(.A1(new_n490), .A2(new_n491), .A3(new_n294), .ZN(new_n492));
  OAI211_X1 g0292(.A(G169), .B(new_n487), .C1(new_n492), .C2(new_n478), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT21), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT21), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n480), .A2(new_n495), .A3(G169), .A4(new_n487), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n489), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n323), .A2(new_n204), .A3(G87), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT22), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n346), .A2(KEYINPUT22), .A3(G87), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G116), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n204), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n212), .A2(G20), .ZN(new_n505));
  XOR2_X1   g0305(.A(new_n505), .B(KEYINPUT23), .Z(new_n506));
  NAND3_X1  g0306(.A1(new_n500), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT24), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n500), .A2(KEYINPUT24), .A3(new_n504), .A4(new_n506), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n509), .A2(new_n254), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n446), .A2(G107), .ZN(new_n512));
  INV_X1    g0312(.A(new_n266), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n513), .A2(new_n505), .ZN(new_n514));
  XNOR2_X1  g0314(.A(new_n514), .B(KEYINPUT25), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n511), .A2(new_n512), .A3(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n477), .A2(new_n213), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n209), .A2(new_n324), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n346), .B(new_n518), .C1(G257), .C2(new_n324), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G294), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n294), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n517), .A2(new_n521), .A3(new_n464), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n522), .A2(G169), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n523), .B1(new_n455), .B2(new_n522), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n516), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n492), .A2(new_n478), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n487), .B1(new_n526), .B2(G190), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(new_n311), .B2(new_n526), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n497), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  OR2_X1    g0329(.A1(G238), .A2(G1698), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n219), .A2(G1698), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n530), .B(new_n531), .C1(new_n280), .C2(new_n281), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n502), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n276), .ZN(new_n534));
  INV_X1    g0334(.A(G45), .ZN(new_n535));
  OAI21_X1  g0335(.A(G250), .B1(new_n535), .B2(G1), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n276), .B1(new_n433), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n311), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n294), .B1(new_n532), .B2(new_n502), .ZN(new_n540));
  NOR3_X1   g0340(.A1(new_n540), .A2(new_n537), .A3(new_n331), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n446), .A2(G87), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n204), .B(G68), .C1(new_n280), .C2(new_n281), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT19), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(new_n258), .B2(new_n441), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n204), .ZN(new_n549));
  NOR2_X1   g0349(.A1(G87), .A2(G97), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n550), .A2(KEYINPUT79), .A3(new_n212), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT79), .B1(new_n550), .B2(new_n212), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n549), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n443), .B1(new_n547), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n396), .A2(new_n320), .ZN(new_n556));
  NOR3_X1   g0356(.A1(new_n555), .A2(KEYINPUT80), .A3(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT80), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n550), .A2(new_n212), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT79), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n561), .A2(new_n551), .B1(new_n204), .B2(new_n548), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n544), .A2(new_n546), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n254), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n556), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n558), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n542), .B(new_n543), .C1(new_n557), .C2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(KEYINPUT80), .B1(new_n555), .B2(new_n556), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n564), .A2(new_n558), .A3(new_n565), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n568), .A2(new_n569), .B1(new_n396), .B2(new_n446), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n540), .A2(new_n537), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G179), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(new_n271), .B2(new_n571), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n567), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n522), .A2(G190), .ZN(new_n576));
  AND4_X1   g0376(.A1(new_n512), .A2(new_n511), .A3(new_n515), .A4(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n522), .A2(new_n311), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n575), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  AND4_X1   g0380(.A1(new_n408), .A2(new_n468), .A3(new_n529), .A4(new_n580), .ZN(G372));
  INV_X1    g0381(.A(KEYINPUT14), .ZN(new_n582));
  OR2_X1    g0382(.A1(new_n303), .A2(new_n582), .ZN(new_n583));
  OR2_X1    g0383(.A1(new_n305), .A2(KEYINPUT71), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n303), .A2(new_n582), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n305), .A2(KEYINPUT71), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n583), .A2(new_n584), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n269), .ZN(new_n588));
  AOI211_X1 g0388(.A(new_n313), .B(new_n378), .C1(new_n588), .C2(new_n402), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n383), .A2(new_n386), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT83), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n383), .A2(new_n386), .A3(KEYINPUT83), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n335), .B1(new_n589), .B2(new_n594), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n595), .A2(new_n337), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n570), .A2(new_n574), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n497), .A2(new_n525), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n580), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n461), .A2(new_n467), .ZN(new_n601));
  INV_X1    g0401(.A(new_n454), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n598), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT82), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n575), .A2(new_n462), .A3(new_n466), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n605), .B1(new_n606), .B2(KEYINPUT26), .ZN(new_n607));
  OAI22_X1  g0407(.A1(new_n557), .A2(new_n566), .B1(new_n397), .B2(new_n445), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n568), .A2(new_n569), .B1(G87), .B2(new_n446), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n608), .A2(new_n573), .B1(new_n609), .B2(new_n542), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n610), .A2(new_n459), .A3(new_n458), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT26), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(KEYINPUT82), .A3(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n461), .A2(new_n467), .A3(KEYINPUT26), .A4(new_n610), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n607), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n408), .B1(new_n604), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n596), .A2(new_n616), .ZN(G369));
  OR3_X1    g0417(.A1(new_n513), .A2(KEYINPUT27), .A3(G20), .ZN(new_n618));
  OAI21_X1  g0418(.A(KEYINPUT27), .B1(new_n513), .B2(G20), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n618), .A2(G213), .A3(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(G343), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n525), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n577), .A2(new_n579), .B1(new_n516), .B2(new_n622), .ZN(new_n625));
  INV_X1    g0425(.A(new_n525), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n497), .A2(new_n622), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n624), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n487), .A2(new_n622), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n497), .B(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n633), .A2(new_n528), .ZN(new_n634));
  XOR2_X1   g0434(.A(KEYINPUT84), .B(G330), .Z(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n631), .B1(new_n636), .B2(new_n637), .ZN(G399));
  INV_X1    g0438(.A(new_n226), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n639), .A2(G41), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(G1), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n561), .A2(new_n250), .A3(new_n551), .ZN(new_n643));
  OAI22_X1  g0443(.A1(new_n642), .A2(new_n643), .B1(new_n231), .B2(new_n641), .ZN(new_n644));
  XOR2_X1   g0444(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n645));
  XNOR2_X1  g0445(.A(new_n644), .B(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n622), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n511), .A2(new_n512), .A3(new_n515), .A4(new_n576), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n610), .B1(new_n648), .B2(new_n578), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(new_n497), .B2(new_n525), .ZN(new_n650));
  AOI211_X1 g0450(.A(KEYINPUT91), .B(new_n454), .C1(new_n467), .C2(new_n461), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT91), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n652), .B1(new_n601), .B2(new_n602), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n650), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n597), .B(KEYINPUT89), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n461), .A2(new_n467), .A3(new_n610), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT90), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(new_n658), .A3(new_n612), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n658), .B1(new_n657), .B2(new_n612), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n611), .A2(new_n612), .ZN(new_n662));
  NOR3_X1   g0462(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  OAI211_X1 g0463(.A(KEYINPUT29), .B(new_n647), .C1(new_n656), .C2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT92), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n597), .B1(new_n650), .B2(new_n468), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n607), .A2(new_n613), .A3(new_n614), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n622), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT88), .B1(new_n669), .B2(KEYINPUT29), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n647), .B1(new_n615), .B2(new_n604), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT88), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT29), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n657), .A2(new_n612), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(KEYINPUT90), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n659), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n654), .B(new_n655), .C1(new_n678), .C2(new_n662), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n679), .A2(KEYINPUT92), .A3(KEYINPUT29), .A4(new_n647), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n666), .A2(new_n675), .A3(new_n680), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n529), .A2(new_n468), .A3(new_n580), .A4(new_n647), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(KEYINPUT31), .ZN(new_n683));
  INV_X1    g0483(.A(new_n572), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n526), .A2(new_n452), .A3(new_n522), .A4(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n686), .A2(KEYINPUT87), .A3(KEYINPUT30), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT87), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT30), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n688), .B1(new_n685), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n526), .A2(new_n522), .ZN(new_n692));
  INV_X1    g0492(.A(new_n571), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n692), .A2(new_n455), .A3(new_n439), .A4(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n685), .A2(new_n689), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n647), .B1(new_n691), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n683), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n691), .B1(KEYINPUT86), .B2(new_n696), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n696), .A2(KEYINPUT86), .ZN(new_n702));
  OAI211_X1 g0502(.A(KEYINPUT31), .B(new_n622), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n635), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n681), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n646), .B1(new_n706), .B2(G1), .ZN(G364));
  NOR2_X1   g0507(.A1(new_n634), .A2(new_n635), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT93), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n265), .A2(G20), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G45), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n641), .A2(G1), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n709), .A2(new_n636), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n232), .B1(G20), .B2(new_n271), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n331), .A2(G20), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT96), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n718), .A2(G179), .A3(new_n311), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n212), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n718), .A2(G179), .A3(G200), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(G159), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n723), .A2(KEYINPUT32), .A3(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n204), .A2(new_n455), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n726), .A2(new_n331), .A3(new_n311), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n727), .A2(KEYINPUT95), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(KEYINPUT95), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  AOI211_X1 g0531(.A(new_n721), .B(new_n725), .C1(G77), .C2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G179), .A2(G200), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n204), .B1(new_n733), .B2(G190), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n726), .A2(G190), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n311), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI221_X1 g0537(.A(new_n323), .B1(new_n441), .B2(new_n734), .C1(new_n737), .C2(new_n216), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT32), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n739), .B1(new_n722), .B2(G159), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n726), .A2(new_n331), .A3(G200), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI211_X1 g0542(.A(new_n738), .B(new_n740), .C1(G68), .C2(new_n742), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n732), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n735), .A2(G200), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n311), .A2(G179), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n747), .A2(G20), .A3(G190), .ZN(new_n748));
  OAI221_X1 g0548(.A(new_n744), .B1(new_n221), .B2(new_n746), .C1(new_n208), .C2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n323), .ZN(new_n750));
  INV_X1    g0550(.A(G294), .ZN(new_n751));
  INV_X1    g0551(.A(G322), .ZN(new_n752));
  OAI221_X1 g0552(.A(new_n750), .B1(new_n751), .B2(new_n734), .C1(new_n746), .C2(new_n752), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n722), .A2(G329), .B1(G326), .B2(new_n736), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n748), .B(KEYINPUT97), .Z(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G303), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g0557(.A(KEYINPUT33), .B(G317), .ZN(new_n758));
  AOI211_X1 g0558(.A(new_n753), .B(new_n757), .C1(new_n742), .C2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G283), .ZN(new_n760));
  INV_X1    g0560(.A(G311), .ZN(new_n761));
  OAI221_X1 g0561(.A(new_n759), .B1(new_n760), .B2(new_n720), .C1(new_n761), .C2(new_n727), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n715), .B1(new_n749), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G13), .A2(G33), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n714), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n323), .A2(new_n226), .A3(G355), .ZN(new_n768));
  AND2_X1   g0568(.A1(new_n247), .A2(G45), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n639), .A2(new_n346), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(new_n231), .B2(new_n272), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n768), .B1(G116), .B2(new_n226), .C1(new_n769), .C2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n763), .B1(new_n767), .B2(new_n772), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n712), .B(KEYINPUT94), .Z(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n766), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n773), .B(new_n775), .C1(new_n634), .C2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n713), .A2(new_n777), .ZN(G396));
  OAI21_X1  g0578(.A(new_n405), .B1(new_n404), .B2(new_n647), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n402), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n402), .A2(new_n622), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n669), .A2(new_n783), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n622), .B(new_n782), .C1(new_n667), .C2(new_n668), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(new_n705), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n712), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G143), .A2(new_n745), .B1(new_n742), .B2(G150), .ZN(new_n789));
  INV_X1    g0589(.A(G137), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n789), .B1(new_n790), .B2(new_n737), .C1(new_n730), .C2(new_n724), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n791), .B(KEYINPUT34), .Z(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n344), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n755), .A2(G50), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n722), .A2(G132), .ZN(new_n795));
  INV_X1    g0595(.A(new_n734), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n719), .A2(G68), .B1(G58), .B2(new_n796), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n793), .A2(new_n794), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n745), .A2(G294), .B1(G97), .B2(new_n796), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT98), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n323), .B(new_n800), .C1(G116), .C2(new_n731), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n755), .A2(G107), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n720), .A2(new_n208), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(G303), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n723), .A2(new_n761), .B1(new_n805), .B2(new_n737), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(G283), .B2(new_n742), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n801), .A2(new_n802), .A3(new_n804), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n798), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n774), .B1(new_n809), .B2(new_n714), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n714), .A2(new_n764), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n810), .B1(G77), .B2(new_n812), .C1(new_n783), .C2(new_n765), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n788), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(G384));
  INV_X1    g0615(.A(new_n620), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n384), .A2(new_n816), .B1(new_n385), .B2(new_n342), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT37), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n817), .A2(new_n818), .A3(new_n376), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT100), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n817), .A2(new_n376), .A3(KEYINPUT100), .A4(new_n818), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n348), .A2(new_n350), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n359), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n342), .B1(new_n353), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n816), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n828), .B(new_n376), .C1(new_n382), .C2(new_n826), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(KEYINPUT37), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n823), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n816), .B(new_n827), .C1(new_n378), .C2(new_n387), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n831), .A2(new_n832), .A3(KEYINPUT38), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n376), .B(KEYINPUT17), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n592), .A2(new_n834), .A3(new_n593), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n361), .A2(new_n620), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n817), .A2(new_n376), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(KEYINPUT37), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n835), .A2(new_n836), .B1(new_n823), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n833), .B1(new_n839), .B2(KEYINPUT38), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT39), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT38), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n821), .A2(new_n822), .B1(KEYINPUT37), .B2(new_n829), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n828), .B1(new_n834), .B2(new_n590), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n833), .A2(new_n846), .A3(KEYINPUT39), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n842), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n588), .A2(new_n622), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n833), .A2(new_n846), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n269), .A2(new_n622), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n853), .B(KEYINPUT99), .Z(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n308), .B2(new_n313), .ZN(new_n856));
  INV_X1    g0656(.A(new_n313), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n588), .A2(new_n857), .A3(new_n854), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n781), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n852), .B(new_n859), .C1(new_n785), .C2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n594), .A2(new_n620), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT101), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n861), .A2(KEYINPUT101), .A3(new_n862), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n851), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n666), .A2(new_n675), .A3(new_n408), .A4(new_n680), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n596), .ZN(new_n868));
  XOR2_X1   g0668(.A(new_n866), .B(new_n868), .Z(new_n869));
  INV_X1    g0669(.A(KEYINPUT40), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n782), .B1(new_n856), .B2(new_n858), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n698), .B1(new_n682), .B2(KEYINPUT31), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n698), .A2(KEYINPUT31), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n833), .A2(new_n846), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n870), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OR2_X1    g0676(.A1(new_n872), .A2(new_n873), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n840), .A2(new_n877), .A3(KEYINPUT40), .A4(new_n871), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n408), .A2(new_n877), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n879), .B(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n635), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n869), .B(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n203), .B2(new_n710), .ZN(new_n884));
  OAI211_X1 g0684(.A(G20), .B(new_n292), .C1(new_n416), .C2(KEYINPUT35), .ZN(new_n885));
  AOI211_X1 g0685(.A(new_n250), .B(new_n885), .C1(KEYINPUT35), .C2(new_n416), .ZN(new_n886));
  XOR2_X1   g0686(.A(new_n886), .B(KEYINPUT36), .Z(new_n887));
  OAI21_X1  g0687(.A(G77), .B1(new_n221), .B2(new_n229), .ZN(new_n888));
  OAI22_X1  g0688(.A1(new_n231), .A2(new_n888), .B1(G50), .B2(new_n229), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n889), .A2(G1), .A3(new_n265), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n884), .A2(new_n887), .A3(new_n890), .ZN(G367));
  INV_X1    g0691(.A(new_n770), .ZN(new_n892));
  OAI221_X1 g0692(.A(new_n767), .B1(new_n226), .B2(new_n397), .C1(new_n242), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n775), .A2(new_n893), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n894), .B(KEYINPUT108), .Z(new_n895));
  OAI22_X1  g0695(.A1(new_n730), .A2(new_n216), .B1(new_n724), .B2(new_n741), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n323), .B1(new_n720), .B2(new_n218), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n896), .B(new_n897), .C1(G68), .C2(new_n796), .ZN(new_n898));
  INV_X1    g0698(.A(new_n748), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n736), .A2(G143), .B1(new_n899), .B2(G58), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  OAI221_X1 g0701(.A(new_n901), .B1(new_n790), .B2(new_n723), .C1(new_n316), .C2(new_n746), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n741), .A2(new_n751), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT46), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n748), .B2(new_n250), .ZN(new_n905));
  OAI221_X1 g0705(.A(new_n905), .B1(new_n746), .B2(new_n805), .C1(new_n761), .C2(new_n737), .ZN(new_n906));
  AOI211_X1 g0706(.A(new_n346), .B(new_n906), .C1(G317), .C2(new_n722), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n755), .A2(KEYINPUT46), .A3(G116), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n908), .B(KEYINPUT109), .Z(new_n909));
  NAND2_X1  g0709(.A1(new_n796), .A2(G107), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n731), .A2(G283), .B1(new_n719), .B2(G97), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n907), .A2(new_n909), .A3(new_n910), .A4(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n902), .B1(new_n903), .B2(new_n912), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n913), .B(KEYINPUT47), .Z(new_n914));
  OAI21_X1  g0714(.A(new_n895), .B1(new_n914), .B2(new_n715), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT110), .Z(new_n916));
  NOR2_X1   g0716(.A1(new_n609), .A2(new_n647), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n597), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n575), .B2(new_n917), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n916), .B1(new_n776), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n711), .A2(G1), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT106), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n468), .B(new_n652), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n459), .A2(new_n622), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(KEYINPUT102), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT102), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n923), .A2(new_n927), .A3(new_n924), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n458), .A2(new_n459), .A3(new_n622), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n926), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n631), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(KEYINPUT45), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n926), .A2(new_n928), .ZN(new_n933));
  XOR2_X1   g0733(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n934));
  NAND4_X1  g0734(.A1(new_n933), .A2(new_n630), .A3(new_n929), .A4(new_n934), .ZN(new_n935));
  OAI211_X1 g0735(.A(KEYINPUT105), .B(KEYINPUT44), .C1(new_n930), .C2(new_n631), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT45), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n930), .A2(new_n937), .A3(new_n631), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n932), .A2(new_n935), .A3(new_n936), .A4(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n636), .A2(new_n637), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n922), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n637), .B(new_n628), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(new_n636), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n681), .A2(new_n705), .A3(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT107), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n939), .A2(new_n940), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(KEYINPUT106), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n943), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n706), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n640), .B(KEYINPUT41), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n921), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT42), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n637), .A2(new_n629), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n954), .B1(new_n930), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n930), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n601), .B1(new_n957), .B2(new_n525), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n956), .B1(new_n958), .B2(new_n647), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n930), .A2(new_n954), .A3(new_n955), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(KEYINPUT103), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT103), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n930), .A2(new_n962), .A3(new_n954), .A4(new_n955), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n959), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n919), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT43), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(KEYINPUT104), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT104), .ZN(new_n970));
  INV_X1    g0770(.A(new_n968), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n959), .A2(new_n970), .A3(new_n971), .A4(new_n964), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n919), .A2(KEYINPUT43), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n965), .A2(new_n968), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n930), .A2(new_n940), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n973), .A2(new_n940), .A3(new_n930), .A4(new_n975), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n920), .B1(new_n953), .B2(new_n980), .ZN(G387));
  NOR2_X1   g0781(.A1(new_n748), .A2(new_n218), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n719), .A2(G97), .B1(G50), .B2(new_n745), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n983), .B1(new_n316), .B2(new_n723), .C1(new_n317), .C2(new_n741), .ZN(new_n984));
  INV_X1    g0784(.A(new_n727), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n982), .B(new_n984), .C1(G68), .C2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n796), .A2(new_n396), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n736), .A2(G159), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n986), .A2(new_n346), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  AOI22_X1  g0789(.A1(G317), .A2(new_n745), .B1(new_n742), .B2(G311), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(new_n752), .B2(new_n737), .C1(new_n730), .C2(new_n805), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT48), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n992), .B1(new_n760), .B2(new_n734), .C1(new_n751), .C2(new_n748), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT49), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n719), .A2(G116), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n722), .A2(G326), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n995), .A2(new_n344), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n993), .A2(new_n994), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n989), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n714), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n394), .A2(new_n216), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT50), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n229), .A2(new_n218), .ZN(new_n1004));
  NOR4_X1   g0804(.A1(new_n1003), .A2(G45), .A3(new_n1004), .A4(new_n643), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n272), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n770), .B1(new_n238), .B2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n643), .A2(new_n226), .A3(new_n323), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1005), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n226), .A2(G107), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n767), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1001), .A2(new_n775), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n637), .B2(new_n766), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n945), .B2(new_n921), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n947), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n706), .B2(new_n945), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1014), .B1(new_n1016), .B2(new_n641), .ZN(G393));
  OR2_X1    g0817(.A1(new_n941), .A2(new_n942), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n1015), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n950), .A2(new_n1019), .A3(new_n640), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n921), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n957), .A2(new_n766), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT111), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n767), .B1(new_n441), .B2(new_n226), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n251), .B2(new_n770), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n804), .B1(new_n218), .B2(new_n734), .C1(new_n317), .C2(new_n730), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G150), .A2(new_n736), .B1(new_n745), .B2(G159), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT51), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n346), .B1(new_n741), .B2(new_n216), .ZN(new_n1030));
  NOR3_X1   g0830(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n229), .B2(new_n748), .ZN(new_n1032));
  AND2_X1   g0832(.A1(new_n722), .A2(G143), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n734), .A2(new_n250), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n721), .B1(G303), .B2(new_n742), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(G311), .A2(new_n745), .B1(new_n736), .B2(G317), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT52), .Z(new_n1037));
  NAND2_X1  g0837(.A1(new_n985), .A2(G294), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n750), .B1(new_n760), .B2(new_n748), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G322), .B2(new_n722), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1035), .A2(new_n1037), .A3(new_n1038), .A4(new_n1040), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n1032), .A2(new_n1033), .B1(new_n1034), .B2(new_n1041), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n774), .B(new_n1026), .C1(new_n1042), .C2(new_n714), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1024), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1020), .A2(new_n1022), .A3(new_n1044), .ZN(G390));
  NOR2_X1   g0845(.A1(new_n748), .A2(new_n316), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT53), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n722), .A2(G125), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1047), .A2(new_n1048), .A3(new_n323), .ZN(new_n1049));
  XOR2_X1   g0849(.A(KEYINPUT54), .B(G143), .Z(new_n1050));
  AOI21_X1  g0850(.A(new_n1049), .B1(new_n731), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n736), .A2(G128), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n719), .A2(G50), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n742), .A2(G137), .B1(new_n796), .B2(G159), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(G132), .B2(new_n745), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n737), .A2(new_n760), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n745), .A2(G116), .B1(G77), .B2(new_n796), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT114), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n731), .A2(G97), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n323), .B1(G107), .B2(new_n742), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n755), .A2(G87), .B1(new_n719), .B2(G68), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1057), .B(new_n1063), .C1(G294), .C2(new_n722), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n714), .B1(new_n1056), .B2(new_n1064), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n1065), .A2(new_n775), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(new_n394), .B2(new_n812), .C1(new_n849), .C2(new_n765), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n850), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n859), .B1(new_n785), .B2(new_n860), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1068), .A2(new_n1069), .B1(new_n842), .B2(new_n847), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n647), .B(new_n780), .C1(new_n656), .C2(new_n663), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n781), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n859), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT112), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n840), .A2(new_n1068), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n859), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n1071), .B2(new_n781), .ZN(new_n1079));
  OAI21_X1  g0879(.A(KEYINPUT112), .B1(new_n1079), .B2(new_n1075), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1070), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n877), .A2(G330), .A3(new_n871), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n704), .A2(new_n635), .A3(new_n783), .A4(new_n859), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1085), .B(new_n1070), .C1(new_n1077), .C2(new_n1080), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1067), .B1(new_n1087), .B2(new_n1021), .ZN(new_n1088));
  OAI211_X1 g0888(.A(G330), .B(new_n783), .C1(new_n872), .C2(new_n873), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n1078), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1085), .A2(new_n1090), .A3(new_n781), .A4(new_n1071), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(KEYINPUT113), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1071), .A2(new_n781), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT113), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1093), .A2(new_n1094), .A3(new_n1085), .A4(new_n1090), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n703), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n635), .B(new_n783), .C1(new_n1096), .C2(new_n872), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n1078), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n1082), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n781), .B1(new_n671), .B2(new_n782), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1092), .A2(new_n1095), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n880), .A2(G330), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n867), .A2(new_n596), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1087), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1070), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1074), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1108));
  NOR3_X1   g0908(.A1(new_n1079), .A2(KEYINPUT112), .A3(new_n1075), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1107), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n1082), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1085), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1107), .B(new_n1112), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1105), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1114), .A2(new_n641), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1088), .B1(new_n1106), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(G378));
  NAND3_X1  g0917(.A1(new_n876), .A2(G330), .A3(new_n878), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1119));
  XOR2_X1   g0919(.A(new_n1119), .B(KEYINPUT120), .Z(new_n1120));
  XNOR2_X1  g0920(.A(new_n338), .B(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n321), .A2(new_n816), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1120), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n338), .B(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n1122), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1118), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1130), .A2(G330), .A3(new_n876), .A4(new_n878), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n866), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n865), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1134), .A2(new_n863), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1135), .A2(new_n851), .A3(new_n1131), .A4(new_n1129), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n921), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n742), .A2(G97), .B1(new_n985), .B2(new_n396), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n293), .B(new_n344), .C1(new_n748), .C2(new_n218), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n1139), .A2(KEYINPUT116), .B1(KEYINPUT115), .B2(new_n1140), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n736), .A2(G116), .B1(G68), .B2(new_n796), .ZN(new_n1142));
  XOR2_X1   g0942(.A(new_n1142), .B(KEYINPUT117), .Z(new_n1143));
  NAND2_X1  g0943(.A1(new_n1140), .A2(KEYINPUT115), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n719), .A2(G58), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n1141), .B(new_n1146), .C1(KEYINPUT116), .C2(new_n1139), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1147), .B1(new_n212), .B2(new_n746), .C1(new_n760), .C2(new_n723), .ZN(new_n1148));
  XOR2_X1   g0948(.A(new_n1148), .B(KEYINPUT58), .Z(new_n1149));
  OAI21_X1  g0949(.A(new_n216), .B1(new_n280), .B2(G41), .ZN(new_n1150));
  AOI21_X1  g0950(.A(G33), .B1(new_n722), .B2(G124), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1151), .B(new_n293), .C1(new_n724), .C2(new_n720), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT118), .Z(new_n1153));
  AOI22_X1  g0953(.A1(G128), .A2(new_n745), .B1(new_n985), .B2(G137), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n736), .A2(G125), .B1(new_n899), .B2(new_n1050), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n796), .A2(G150), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n742), .A2(G132), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT59), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1150), .B1(new_n1153), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n714), .B1(new_n1149), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n712), .B1(new_n216), .B2(new_n811), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT119), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1161), .B(new_n1163), .C1(new_n1128), .C2(new_n765), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n1164), .B(KEYINPUT121), .Z(new_n1165));
  NAND2_X1  g0965(.A1(new_n1138), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n867), .A2(new_n596), .A3(new_n1103), .ZN(new_n1168));
  OAI211_X1 g0968(.A(KEYINPUT57), .B(new_n1137), .C1(new_n1114), .C2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n640), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n1104), .ZN(new_n1173));
  AOI21_X1  g0973(.A(KEYINPUT57), .B1(new_n1173), .B2(new_n1137), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1167), .B1(new_n1170), .B2(new_n1174), .ZN(G375));
  AND2_X1   g0975(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT122), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1176), .A2(new_n1177), .A3(new_n1101), .A4(new_n1168), .ZN(new_n1178));
  OAI21_X1  g0978(.A(KEYINPUT122), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1180), .A2(new_n952), .A3(new_n1105), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1078), .A2(new_n764), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n812), .A2(G68), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n722), .A2(G128), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G132), .A2(new_n736), .B1(new_n745), .B2(G137), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1145), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n755), .A2(G159), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n346), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1186), .B(new_n1188), .C1(new_n742), .C2(new_n1050), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1189), .B1(new_n216), .B2(new_n734), .C1(new_n316), .C2(new_n727), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n987), .B1(new_n746), .B2(new_n760), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT123), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n323), .B(new_n1192), .C1(G116), .C2(new_n742), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n755), .A2(G97), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n731), .A2(G107), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(G77), .A2(new_n719), .B1(new_n722), .B2(G303), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n737), .A2(new_n751), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1190), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n774), .B(new_n1183), .C1(new_n1199), .C2(new_n714), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1102), .A2(new_n921), .B1(new_n1182), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1181), .A2(new_n1201), .ZN(G381));
  INV_X1    g1002(.A(G390), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n952), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n950), .B2(new_n706), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n978), .B(new_n979), .C1(new_n1205), .C2(new_n921), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1203), .A2(new_n1206), .A3(new_n920), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(G381), .A2(G384), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(G393), .A2(G396), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  OR2_X1    g1011(.A1(new_n1211), .A2(KEYINPUT124), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(G375), .A2(G378), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1211), .A2(KEYINPUT124), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(G407));
  INV_X1    g1015(.A(new_n1213), .ZN(new_n1216));
  OAI211_X1 g1016(.A(G407), .B(G213), .C1(G343), .C2(new_n1216), .ZN(G409));
  XNOR2_X1  g1017(.A(G393), .B(G396), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1203), .B1(new_n1206), .B2(new_n920), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1219), .B1(new_n1208), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(G387), .A2(G390), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1222), .A2(new_n1207), .A3(new_n1218), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(G375), .A2(G378), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n621), .A2(G213), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n1172), .B2(new_n1104), .ZN(new_n1228));
  AOI21_X1  g1028(.A(KEYINPUT125), .B1(new_n1228), .B2(new_n952), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1113), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1168), .B1(new_n1230), .B2(new_n1171), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT125), .ZN(new_n1232));
  NOR4_X1   g1032(.A1(new_n1231), .A2(new_n1232), .A3(new_n1204), .A4(new_n1227), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1116), .B(new_n1167), .C1(new_n1229), .C2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1201), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT60), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n1102), .A2(new_n1104), .A3(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1236), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1237), .B1(new_n1180), .B2(new_n1239), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n814), .B(new_n1235), .C1(new_n1240), .C2(new_n640), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1092), .A2(new_n1101), .A3(new_n1095), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1177), .B1(new_n1242), .B2(new_n1168), .ZN(new_n1243));
  NOR3_X1   g1043(.A1(new_n1102), .A2(new_n1104), .A3(KEYINPUT122), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1239), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1237), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1245), .A2(new_n640), .A3(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(G384), .B1(new_n1247), .B2(new_n1201), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1241), .A2(new_n1248), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1225), .A2(new_n1226), .A3(new_n1234), .A4(new_n1249), .ZN(new_n1250));
  OR2_X1    g1050(.A1(new_n1250), .A2(KEYINPUT62), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(KEYINPUT62), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1224), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT127), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1238), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1255), .A2(new_n641), .A3(new_n1237), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n814), .B1(new_n1256), .B2(new_n1235), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1247), .A2(G384), .A3(new_n1201), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n621), .A2(G213), .A3(G2897), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1259), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n641), .B1(new_n1228), .B2(KEYINPUT57), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT57), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n1231), .B2(new_n1227), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1166), .B1(new_n1263), .B2(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1234), .B(new_n1226), .C1(new_n1266), .C2(new_n1116), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1262), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT61), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1254), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  AOI211_X1 g1070(.A(KEYINPUT127), .B(KEYINPUT61), .C1(new_n1262), .C2(new_n1267), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT63), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1250), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(KEYINPUT126), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT61), .B1(new_n1262), .B2(new_n1267), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1277), .A2(KEYINPUT63), .A3(new_n1234), .A4(new_n1249), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT126), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1250), .A2(new_n1279), .A3(new_n1273), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1275), .A2(new_n1276), .A3(new_n1278), .A4(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1224), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n1253), .A2(new_n1272), .B1(new_n1281), .B2(new_n1282), .ZN(G405));
  AND2_X1   g1083(.A1(new_n1216), .A2(new_n1225), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n1222), .A2(new_n1207), .A3(new_n1218), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1218), .B1(new_n1222), .B2(new_n1207), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1284), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1216), .A2(new_n1225), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1221), .A2(new_n1223), .A3(new_n1288), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1287), .A2(new_n1249), .A3(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1249), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(G402));
endmodule


