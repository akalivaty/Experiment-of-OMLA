//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 1 1 0 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G119), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G128), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n187), .A2(KEYINPUT23), .A3(G119), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G110), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n192), .A2(new_n188), .ZN(new_n196));
  OR2_X1    g010(.A1(new_n196), .A2(KEYINPUT73), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(KEYINPUT73), .ZN(new_n198));
  XOR2_X1   g012(.A(KEYINPUT24), .B(G110), .Z(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G125), .ZN(new_n201));
  NOR3_X1   g015(.A1(new_n201), .A2(KEYINPUT16), .A3(G140), .ZN(new_n202));
  XNOR2_X1  g016(.A(G125), .B(G140), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(KEYINPUT16), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n204), .A2(G146), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n195), .B(new_n200), .C1(new_n206), .C2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT74), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(new_n204), .B(G146), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n211), .A2(KEYINPUT74), .A3(new_n195), .A4(new_n200), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n203), .B(KEYINPUT76), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n194), .A2(G110), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n217), .B(KEYINPUT75), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n199), .B1(new_n197), .B2(new_n198), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n205), .B(new_n216), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n213), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT22), .B(G137), .ZN(new_n222));
  INV_X1    g036(.A(G953), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(G221), .A3(G234), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n222), .B(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n221), .A2(new_n226), .ZN(new_n227));
  XOR2_X1   g041(.A(KEYINPUT72), .B(G902), .Z(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n213), .A2(new_n220), .A3(new_n225), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT25), .ZN(new_n232));
  INV_X1    g046(.A(G217), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n233), .B1(new_n229), .B2(G234), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT25), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n227), .A2(new_n235), .A3(new_n229), .A4(new_n230), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n232), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n227), .A2(new_n230), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n234), .A2(G902), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n237), .A2(KEYINPUT77), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(KEYINPUT77), .B1(new_n237), .B2(new_n240), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT1), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n215), .A2(G143), .ZN(new_n245));
  INV_X1    g059(.A(G143), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G146), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n245), .A2(new_n247), .A3(G128), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT64), .B1(new_n246), .B2(G146), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT64), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(new_n215), .A3(G143), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n249), .A2(new_n251), .A3(new_n247), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n246), .A2(G146), .ZN(new_n253));
  OAI21_X1  g067(.A(G128), .B1(new_n253), .B2(new_n244), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n244), .A2(new_n248), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT11), .ZN(new_n256));
  INV_X1    g070(.A(G134), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n256), .B1(new_n257), .B2(G137), .ZN(new_n258));
  INV_X1    g072(.A(G137), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(KEYINPUT11), .A3(G134), .ZN(new_n260));
  INV_X1    g074(.A(G131), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n257), .A2(G137), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n258), .A2(new_n260), .A3(new_n261), .A4(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n259), .A2(G134), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n257), .A2(G137), .ZN(new_n265));
  OAI21_X1  g079(.A(G131), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT67), .B1(new_n255), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n258), .A2(new_n262), .A3(new_n260), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G131), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n263), .ZN(new_n271));
  AND2_X1   g085(.A1(KEYINPUT0), .A2(G128), .ZN(new_n272));
  NOR2_X1   g086(.A1(KEYINPUT0), .A2(G128), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n245), .A2(new_n247), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n252), .A2(new_n274), .B1(new_n275), .B2(new_n272), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n271), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n252), .A2(new_n254), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n245), .A2(new_n247), .A3(new_n244), .A4(G128), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT67), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n263), .A2(new_n266), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n268), .A2(new_n277), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT30), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n277), .A2(KEYINPUT65), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT30), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT65), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n271), .A2(new_n276), .A3(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT66), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n267), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n263), .A2(new_n266), .A3(KEYINPUT66), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n280), .A3(new_n292), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n286), .A2(new_n287), .A3(new_n289), .A4(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n285), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n191), .A2(G116), .ZN(new_n296));
  INV_X1    g110(.A(G116), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G119), .ZN(new_n298));
  INV_X1    g112(.A(G113), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n299), .A2(KEYINPUT2), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n299), .A2(KEYINPUT2), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n296), .B(new_n298), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n296), .A2(new_n298), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT2), .B(G113), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n295), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n306), .B1(new_n271), .B2(new_n276), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n268), .A2(new_n308), .A3(new_n283), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT68), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT68), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n268), .A2(new_n308), .A3(new_n311), .A4(new_n283), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(G237), .A2(G953), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G210), .ZN(new_n316));
  INV_X1    g130(.A(G101), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n316), .B(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n318), .B(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n314), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT29), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT69), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n280), .A2(new_n282), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n308), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT28), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n324), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AOI211_X1 g142(.A(KEYINPUT69), .B(KEYINPUT28), .C1(new_n308), .C2(new_n325), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT71), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT71), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n332), .B1(new_n328), .B2(new_n329), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n284), .A2(new_n306), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n313), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(KEYINPUT70), .A3(KEYINPUT28), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT70), .ZN(new_n338));
  AOI22_X1  g152(.A1(new_n310), .A2(new_n312), .B1(new_n306), .B2(new_n284), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n338), .B1(new_n339), .B2(new_n327), .ZN(new_n340));
  INV_X1    g154(.A(new_n320), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n334), .A2(new_n337), .A3(new_n340), .A4(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n286), .A2(new_n289), .A3(new_n293), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n306), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n327), .B1(new_n313), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n330), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n320), .A2(KEYINPUT29), .ZN(new_n348));
  AOI22_X1  g162(.A1(new_n323), .A2(new_n342), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(G472), .B1(new_n349), .B2(new_n228), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n307), .A2(new_n341), .A3(new_n313), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT31), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n320), .B1(new_n345), .B2(new_n346), .ZN(new_n353));
  AOI22_X1  g167(.A1(new_n295), .A2(new_n306), .B1(new_n312), .B2(new_n310), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT31), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(new_n341), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n352), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(G472), .A2(G902), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT32), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT32), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n357), .A2(new_n361), .A3(new_n358), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n243), .B1(new_n350), .B2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT85), .B(G469), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(G110), .B(G140), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n367), .B(KEYINPUT79), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n223), .A2(G227), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n368), .B(new_n369), .ZN(new_n370));
  OR2_X1    g184(.A1(KEYINPUT80), .A2(G104), .ZN(new_n371));
  NAND2_X1  g185(.A1(KEYINPUT80), .A2(G104), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n373));
  INV_X1    g187(.A(G107), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n371), .A2(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n373), .A2(new_n374), .A3(G104), .ZN(new_n376));
  NAND2_X1  g190(.A1(KEYINPUT3), .A2(G107), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(G101), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  AND2_X1   g193(.A1(KEYINPUT80), .A2(G104), .ZN(new_n380));
  NOR2_X1   g194(.A1(KEYINPUT80), .A2(G104), .ZN(new_n381));
  OAI22_X1  g195(.A1(new_n380), .A2(new_n381), .B1(KEYINPUT3), .B2(G107), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n382), .A2(new_n317), .A3(new_n377), .A4(new_n376), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n379), .A2(KEYINPUT4), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT4), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n385), .B(G101), .C1(new_n375), .C2(new_n378), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n276), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT81), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n371), .A2(new_n388), .A3(new_n374), .A4(new_n372), .ZN(new_n389));
  NOR3_X1   g203(.A1(new_n380), .A2(new_n381), .A3(G107), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT81), .B1(new_n374), .B2(G104), .ZN(new_n391));
  OAI211_X1 g205(.A(G101), .B(new_n389), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n187), .B1(new_n245), .B2(KEYINPUT1), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n279), .B1(new_n275), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n383), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT10), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n280), .A2(KEYINPUT10), .A3(new_n383), .A4(new_n392), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n387), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n271), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT84), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n399), .A2(KEYINPUT84), .A3(new_n271), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n271), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n387), .A2(new_n397), .A3(new_n405), .A4(new_n398), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n370), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n370), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT82), .ZN(new_n409));
  AOI21_X1  g223(.A(KEYINPUT12), .B1(new_n271), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n392), .A2(new_n383), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n255), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n395), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n411), .B1(new_n414), .B2(new_n271), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n271), .A3(new_n411), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n408), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n229), .B(new_n366), .C1(new_n407), .C2(new_n418), .ZN(new_n419));
  AOI211_X1 g233(.A(new_n405), .B(new_n410), .C1(new_n395), .C2(new_n413), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n406), .B1(new_n420), .B2(new_n415), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT83), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n370), .ZN(new_n424));
  OAI211_X1 g238(.A(KEYINPUT83), .B(new_n406), .C1(new_n420), .C2(new_n415), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n404), .A2(new_n370), .A3(new_n406), .ZN(new_n427));
  AOI21_X1  g241(.A(G902), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G469), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n419), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  XOR2_X1   g244(.A(KEYINPUT9), .B(G234), .Z(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G221), .B1(new_n432), .B2(G902), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n433), .B(KEYINPUT78), .Z(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n430), .A2(KEYINPUT86), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT86), .B1(new_n430), .B2(new_n435), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n223), .A2(G952), .ZN(new_n439));
  NAND2_X1  g253(.A1(G234), .A2(G237), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n441), .B(KEYINPUT99), .ZN(new_n442));
  XOR2_X1   g256(.A(KEYINPUT21), .B(G898), .Z(new_n443));
  NAND3_X1  g257(.A1(new_n228), .A2(G953), .A3(new_n440), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(G214), .B1(G237), .B2(G902), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n278), .A2(new_n201), .A3(new_n279), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n447), .B1(new_n201), .B2(new_n276), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n223), .A2(G224), .ZN(new_n449));
  XOR2_X1   g263(.A(new_n449), .B(KEYINPUT88), .Z(new_n450));
  XNOR2_X1  g264(.A(new_n448), .B(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT6), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n384), .A2(new_n306), .A3(new_n386), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n296), .A2(new_n298), .A3(KEYINPUT5), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n454), .B(G113), .C1(KEYINPUT5), .C2(new_n296), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n392), .A2(new_n302), .A3(new_n383), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT87), .ZN(new_n458));
  XOR2_X1   g272(.A(G110), .B(G122), .Z(new_n459));
  INV_X1    g273(.A(KEYINPUT87), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n453), .A2(new_n460), .A3(new_n456), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n458), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  OR2_X1    g276(.A1(new_n457), .A2(new_n459), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n452), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n453), .A2(new_n460), .A3(new_n456), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n460), .B1(new_n453), .B2(new_n456), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(KEYINPUT6), .B1(new_n467), .B2(new_n459), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n451), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT89), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n455), .A2(new_n302), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n412), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n470), .B1(new_n412), .B2(new_n471), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n456), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  XOR2_X1   g288(.A(new_n459), .B(KEYINPUT8), .Z(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n449), .A2(KEYINPUT7), .ZN(new_n477));
  OR2_X1    g291(.A1(new_n477), .A2(KEYINPUT90), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n447), .B(new_n478), .C1(new_n201), .C2(new_n276), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(KEYINPUT90), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n479), .B(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n476), .A2(new_n463), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(G902), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT91), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n483), .A2(KEYINPUT91), .A3(new_n484), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n469), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(G210), .B1(G237), .B2(G902), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n469), .A2(new_n487), .A3(new_n490), .A4(new_n488), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n445), .B(new_n446), .C1(new_n492), .C2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G237), .ZN(new_n496));
  AND4_X1   g310(.A1(G143), .A2(new_n496), .A3(new_n223), .A4(G214), .ZN(new_n497));
  AOI21_X1  g311(.A(G143), .B1(new_n315), .B2(G214), .ZN(new_n498));
  OAI21_X1  g312(.A(G131), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT93), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n496), .A2(new_n223), .A3(G214), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n246), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n315), .A2(G143), .A3(G214), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT93), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(new_n505), .A3(G131), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n500), .A2(KEYINPUT17), .A3(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT94), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n500), .A2(new_n506), .A3(KEYINPUT94), .A4(KEYINPUT17), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n211), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT95), .ZN(new_n514));
  INV_X1    g328(.A(new_n504), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n500), .A2(new_n506), .B1(new_n261), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT95), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n511), .A2(new_n519), .A3(new_n512), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n514), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(G113), .B(G122), .ZN(new_n522));
  XOR2_X1   g336(.A(new_n522), .B(G104), .Z(new_n523));
  NAND2_X1  g337(.A1(new_n515), .A2(KEYINPUT92), .ZN(new_n524));
  NAND2_X1  g338(.A1(KEYINPUT18), .A2(G131), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n524), .B(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n216), .B1(new_n215), .B2(new_n203), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n521), .A2(new_n523), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n523), .B1(new_n521), .B2(new_n528), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n484), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(G475), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n432), .A2(new_n233), .A3(G953), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT96), .ZN(new_n535));
  INV_X1    g349(.A(G122), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n535), .B1(new_n536), .B2(G116), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n297), .A2(KEYINPUT96), .A3(G122), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n297), .A2(G122), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n540), .A2(G107), .A3(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(G128), .B(G143), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(G134), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n539), .A2(KEYINPUT14), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT97), .ZN(new_n546));
  INV_X1    g360(.A(new_n541), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT14), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n540), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n549), .B1(new_n537), .B2(new_n538), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT97), .B1(new_n551), .B2(new_n541), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n548), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  AOI211_X1 g367(.A(new_n542), .B(new_n544), .C1(new_n553), .C2(G107), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n543), .A2(KEYINPUT13), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n246), .A2(G128), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n555), .B(G134), .C1(KEYINPUT13), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n543), .A2(new_n257), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n374), .B1(new_n539), .B2(new_n547), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n557), .B(new_n558), .C1(new_n542), .C2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n534), .B1(new_n554), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT98), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n553), .A2(G107), .ZN(new_n564));
  INV_X1    g378(.A(new_n542), .ZN(new_n565));
  INV_X1    g379(.A(new_n544), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n560), .A3(new_n533), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n562), .A2(new_n563), .A3(new_n568), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n567), .A2(KEYINPUT98), .A3(new_n560), .A4(new_n533), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(new_n229), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(G478), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(KEYINPUT15), .ZN(new_n573));
  XOR2_X1   g387(.A(new_n571), .B(new_n573), .Z(new_n574));
  INV_X1    g388(.A(KEYINPUT20), .ZN(new_n575));
  INV_X1    g389(.A(new_n516), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT19), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n214), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n577), .B2(new_n203), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n576), .B(new_n205), .C1(new_n579), .C2(G146), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n580), .A2(new_n528), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(new_n523), .ZN(new_n582));
  INV_X1    g396(.A(new_n528), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n519), .B1(new_n511), .B2(new_n512), .ZN(new_n584));
  AOI211_X1 g398(.A(KEYINPUT95), .B(new_n211), .C1(new_n509), .C2(new_n510), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n583), .B1(new_n586), .B2(new_n518), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n582), .B1(new_n587), .B2(new_n523), .ZN(new_n588));
  NOR2_X1   g402(.A1(G475), .A2(G902), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n575), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n521), .A2(new_n523), .A3(new_n528), .ZN(new_n592));
  OR2_X1    g406(.A1(new_n581), .A2(new_n523), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n594), .A2(KEYINPUT20), .A3(new_n589), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n532), .A2(new_n574), .A3(new_n591), .A4(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n495), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n364), .A2(new_n438), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(G101), .ZN(G3));
  NOR3_X1   g413(.A1(new_n436), .A2(new_n243), .A3(new_n437), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n532), .A2(new_n591), .A3(new_n595), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n571), .A2(new_n572), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT101), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT33), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n569), .A2(new_n604), .A3(new_n570), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n562), .A2(KEYINPUT33), .A3(new_n568), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT100), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n228), .A2(new_n572), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n562), .A2(KEYINPUT100), .A3(new_n568), .A4(KEYINPUT33), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n605), .A2(new_n608), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT101), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n571), .A2(new_n612), .A3(new_n572), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n603), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n601), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(new_n495), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n357), .A2(new_n229), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n617), .A2(G472), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n358), .B2(new_n357), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n600), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT34), .B(G104), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G6));
  XOR2_X1   g436(.A(new_n445), .B(KEYINPUT102), .Z(new_n623));
  OAI211_X1 g437(.A(new_n446), .B(new_n623), .C1(new_n492), .C2(new_n494), .ZN(new_n624));
  AOI21_X1  g438(.A(KEYINPUT20), .B1(new_n594), .B2(new_n589), .ZN(new_n625));
  AOI211_X1 g439(.A(new_n575), .B(new_n590), .C1(new_n592), .C2(new_n593), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n574), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(new_n628), .A3(new_n532), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n600), .A2(new_n619), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT35), .B(G107), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  NOR2_X1   g447(.A1(new_n226), .A2(KEYINPUT36), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n221), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n239), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n237), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n438), .A2(new_n597), .A3(new_n619), .A4(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT37), .B(G110), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G12));
  OAI21_X1  g454(.A(new_n442), .B1(G900), .B2(new_n444), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n629), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n637), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n363), .B2(new_n350), .ZN(new_n645));
  INV_X1    g459(.A(new_n446), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n489), .A2(new_n491), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n646), .B1(new_n647), .B2(new_n493), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n438), .A2(new_n643), .A3(new_n645), .A4(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT103), .B(G128), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G30));
  INV_X1    g465(.A(new_n438), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n641), .B(KEYINPUT39), .Z(new_n653));
  NOR2_X1   g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n637), .B1(new_n655), .B2(KEYINPUT40), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n647), .A2(new_n493), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n657), .B(KEYINPUT38), .Z(new_n658));
  NAND2_X1  g472(.A1(new_n314), .A2(new_n341), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n659), .B(new_n484), .C1(new_n341), .C2(new_n336), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(G472), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n363), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n601), .A2(new_n628), .ZN(new_n664));
  NOR4_X1   g478(.A1(new_n658), .A2(new_n663), .A3(new_n646), .A4(new_n664), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n656), .B(new_n665), .C1(KEYINPUT40), .C2(new_n655), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G143), .ZN(G45));
  NAND3_X1  g481(.A1(new_n438), .A2(new_n648), .A3(new_n645), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n591), .A2(new_n595), .ZN(new_n669));
  INV_X1    g483(.A(G475), .ZN(new_n670));
  INV_X1    g484(.A(new_n530), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n592), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n670), .B1(new_n672), .B2(new_n484), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n614), .B(new_n641), .C1(new_n669), .C2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(KEYINPUT104), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT104), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n601), .A2(new_n676), .A3(new_n614), .A4(new_n641), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n668), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(new_n215), .ZN(G48));
  INV_X1    g494(.A(new_n403), .ZN(new_n681));
  AOI21_X1  g495(.A(KEYINPUT84), .B1(new_n399), .B2(new_n271), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n406), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n418), .B1(new_n683), .B2(new_n424), .ZN(new_n684));
  OAI21_X1  g498(.A(G469), .B1(new_n684), .B2(new_n228), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n419), .A3(new_n435), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT105), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n685), .A2(new_n419), .A3(KEYINPUT105), .A4(new_n435), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n364), .A2(new_n616), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT41), .B(G113), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G15));
  NAND3_X1  g507(.A1(new_n364), .A2(new_n630), .A3(new_n690), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G116), .ZN(G18));
  NAND3_X1  g509(.A1(new_n597), .A2(new_n645), .A3(new_n690), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  INV_X1    g511(.A(new_n623), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n664), .A2(new_n698), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n352), .A2(new_n356), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n334), .A2(new_n337), .A3(new_n340), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n320), .ZN(new_n702));
  AOI211_X1 g516(.A(G472), .B(G902), .C1(new_n700), .C2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n237), .A2(new_n240), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n703), .A2(new_n618), .A3(new_n704), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n648), .A2(new_n688), .A3(new_n689), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n699), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT106), .B(G122), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G24));
  NOR3_X1   g523(.A1(new_n703), .A2(new_n618), .A3(new_n644), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n675), .A2(new_n677), .A3(new_n706), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G125), .ZN(G27));
  NAND2_X1  g526(.A1(new_n430), .A2(new_n435), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n657), .A2(new_n646), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n675), .A2(new_n714), .A3(new_n677), .A4(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n364), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n704), .B1(new_n363), .B2(new_n350), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT42), .ZN(new_n720));
  OAI22_X1  g534(.A1(new_n718), .A2(KEYINPUT42), .B1(new_n716), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT107), .B(G131), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G33));
  AND4_X1   g537(.A1(new_n364), .A2(new_n714), .A3(new_n643), .A4(new_n715), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT108), .B(G134), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G36));
  NOR2_X1   g540(.A1(new_n619), .A2(new_n644), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT110), .ZN(new_n728));
  INV_X1    g542(.A(new_n601), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n614), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(KEYINPUT43), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n728), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(KEYINPUT112), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n426), .A2(new_n427), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT45), .ZN(new_n739));
  OAI21_X1  g553(.A(G469), .B1(new_n739), .B2(G902), .ZN(new_n740));
  XOR2_X1   g554(.A(new_n740), .B(KEYINPUT46), .Z(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n419), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n435), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n653), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n715), .B1(new_n734), .B2(new_n735), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n737), .A2(new_n744), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G137), .ZN(G39));
  NAND2_X1  g564(.A1(new_n363), .A2(new_n350), .ZN(new_n751));
  INV_X1    g565(.A(new_n243), .ZN(new_n752));
  INV_X1    g566(.A(new_n715), .ZN(new_n753));
  NOR4_X1   g567(.A1(new_n678), .A2(new_n751), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  XOR2_X1   g568(.A(new_n754), .B(KEYINPUT113), .Z(new_n755));
  INV_X1    g569(.A(KEYINPUT47), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n743), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n742), .A2(KEYINPUT47), .A3(new_n435), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G140), .ZN(G42));
  INV_X1    g575(.A(new_n442), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n733), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n705), .A3(new_n706), .ZN(new_n764));
  INV_X1    g578(.A(new_n690), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(new_n753), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n763), .A2(new_n719), .A3(new_n766), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n767), .A2(KEYINPUT48), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n766), .A2(new_n752), .A3(new_n762), .A4(new_n663), .ZN(new_n769));
  OAI221_X1 g583(.A(new_n439), .B1(new_n615), .B2(new_n769), .C1(new_n767), .C2(KEYINPUT48), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n763), .A2(new_n705), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n685), .A2(new_n419), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n435), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n771), .B(new_n715), .C1(new_n759), .C2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n763), .A2(new_n710), .A3(new_n766), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OR3_X1    g590(.A1(new_n769), .A2(new_n601), .A3(new_n614), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n690), .A2(KEYINPUT119), .A3(new_n646), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT119), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n779), .B1(new_n765), .B2(new_n446), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n780), .A2(new_n658), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n763), .A2(new_n705), .A3(new_n778), .A4(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n776), .A2(new_n777), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n774), .A2(KEYINPUT120), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT51), .ZN(new_n787));
  AOI211_X1 g601(.A(new_n768), .B(new_n770), .C1(new_n785), .C2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n691), .A2(new_n694), .A3(new_n707), .A4(new_n696), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n789), .A2(KEYINPUT118), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n791), .B1(new_n615), .B2(new_n624), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n603), .A2(new_n611), .A3(new_n613), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n793), .B1(new_n627), .B2(new_n532), .ZN(new_n794));
  AOI211_X1 g608(.A(new_n646), .B(new_n698), .C1(new_n647), .C2(new_n493), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n795), .A3(KEYINPUT114), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n600), .A2(new_n792), .A3(new_n619), .A4(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n797), .A2(new_n631), .A3(new_n598), .A4(new_n638), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n789), .A2(KEYINPUT118), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n790), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n647), .A2(new_n446), .A3(new_n493), .A4(new_n641), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n802), .B1(new_n363), .B2(new_n350), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n438), .A2(new_n574), .A3(new_n803), .A4(new_n729), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n703), .A2(new_n618), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n804), .B1(new_n716), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n724), .B1(new_n806), .B2(new_n637), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n721), .A2(KEYINPUT53), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n801), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n711), .B(new_n649), .C1(new_n668), .C2(new_n678), .ZN(new_n812));
  INV_X1    g626(.A(new_n648), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n664), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n637), .A2(new_n642), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n814), .A2(new_n714), .A3(new_n662), .A4(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n811), .B1(new_n812), .B2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(KEYINPUT115), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n438), .A2(new_n648), .A3(new_n645), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n676), .B1(new_n794), .B2(new_n641), .ZN(new_n823));
  INV_X1    g637(.A(new_n677), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n822), .B1(new_n825), .B2(new_n643), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n826), .A2(KEYINPUT52), .A3(new_n711), .A4(new_n816), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT115), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n818), .A2(new_n820), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n821), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n819), .B1(new_n812), .B2(new_n817), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n832), .A2(new_n827), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n798), .A2(new_n789), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n834), .A2(new_n721), .A3(new_n807), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n831), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT117), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n838), .B(new_n831), .C1(new_n833), .C2(new_n835), .ZN(new_n839));
  AOI221_X4 g653(.A(KEYINPUT54), .B1(new_n810), .B2(new_n830), .C1(new_n837), .C2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n832), .A2(new_n827), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(new_n721), .A3(new_n807), .A4(new_n834), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT53), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n830), .A2(new_n831), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n843), .B1(new_n844), .B2(new_n835), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n840), .B1(KEYINPUT54), .B2(new_n846), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n785), .A2(new_n787), .ZN(new_n848));
  AND4_X1   g662(.A1(new_n764), .A2(new_n788), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(G952), .A2(G953), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT121), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n772), .A2(KEYINPUT49), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n704), .B1(new_n772), .B2(KEYINPUT49), .ZN(new_n853));
  AND4_X1   g667(.A1(new_n435), .A2(new_n852), .A3(new_n853), .A4(new_n446), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n854), .A2(new_n658), .A3(new_n663), .ZN(new_n855));
  OAI22_X1  g669(.A1(new_n849), .A2(new_n851), .B1(new_n730), .B2(new_n855), .ZN(G75));
  NOR2_X1   g670(.A1(new_n464), .A2(new_n468), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(new_n451), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n858), .B(KEYINPUT55), .Z(new_n859));
  NAND2_X1  g673(.A1(new_n810), .A2(new_n830), .ZN(new_n860));
  INV_X1    g674(.A(new_n839), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n838), .B1(new_n842), .B2(new_n831), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n228), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n490), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n859), .B1(new_n865), .B2(KEYINPUT56), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n223), .A2(G952), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n863), .A2(KEYINPUT122), .A3(new_n228), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n491), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n859), .A2(KEYINPUT56), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n869), .B1(new_n873), .B2(new_n874), .ZN(G51));
  NAND2_X1  g689(.A1(G469), .A2(G902), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n876), .B(KEYINPUT57), .Z(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n863), .A2(KEYINPUT54), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n837), .A2(new_n839), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n880), .A2(new_n881), .A3(new_n860), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n878), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT123), .B1(new_n883), .B2(new_n684), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n881), .B1(new_n880), .B2(new_n860), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n877), .B1(new_n840), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT123), .ZN(new_n887));
  INV_X1    g701(.A(new_n684), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n871), .A2(G469), .A3(new_n739), .A4(new_n872), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n884), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n891), .A2(new_n868), .ZN(G54));
  AND2_X1   g706(.A1(KEYINPUT58), .A2(G475), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n871), .A2(new_n872), .A3(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT124), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n894), .A2(new_n895), .A3(new_n588), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n895), .B1(new_n894), .B2(new_n588), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n871), .A2(new_n594), .A3(new_n872), .A4(new_n893), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n868), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n896), .A2(new_n897), .A3(new_n899), .ZN(G60));
  NAND2_X1  g714(.A1(G478), .A2(G902), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT59), .Z(new_n902));
  NOR2_X1   g716(.A1(new_n847), .A2(new_n902), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n605), .A2(new_n608), .A3(new_n610), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n868), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n902), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n879), .B2(new_n882), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n905), .A2(new_n908), .ZN(G63));
  NAND2_X1  g723(.A1(G217), .A2(G902), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT60), .Z(new_n911));
  NAND3_X1  g725(.A1(new_n863), .A2(new_n635), .A3(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n863), .A2(new_n911), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n868), .B(new_n912), .C1(new_n913), .C2(new_n238), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT61), .B1(new_n912), .B2(KEYINPUT125), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n914), .B(new_n915), .ZN(G66));
  NAND2_X1  g730(.A1(new_n443), .A2(G224), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(G953), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n918), .B1(new_n834), .B2(G953), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n857), .B1(G898), .B2(new_n223), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(G69));
  INV_X1    g735(.A(new_n812), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n666), .A2(new_n922), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT62), .Z(new_n924));
  NAND2_X1  g738(.A1(new_n615), .A2(new_n629), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n654), .A2(new_n364), .A3(new_n715), .A4(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n924), .A2(new_n749), .A3(new_n760), .A4(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n223), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n295), .B(new_n579), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n223), .A2(G900), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT126), .Z(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n724), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n744), .A2(new_n719), .A3(new_n814), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n935), .A2(new_n721), .A3(new_n922), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n749), .A2(new_n934), .A3(new_n760), .A4(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n933), .B1(new_n937), .B2(new_n223), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n930), .B1(new_n938), .B2(new_n929), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n223), .B1(G227), .B2(G900), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n940), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n930), .B(new_n942), .C1(new_n929), .C2(new_n938), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n941), .A2(new_n943), .ZN(G72));
  NAND2_X1  g758(.A1(G472), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT63), .Z(new_n946));
  INV_X1    g760(.A(new_n834), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n927), .B2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n659), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n867), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n946), .B1(new_n937), .B2(new_n947), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n951), .A2(new_n320), .A3(new_n354), .ZN(new_n952));
  INV_X1    g766(.A(new_n351), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n321), .B(KEYINPUT127), .Z(new_n954));
  OAI211_X1 g768(.A(new_n846), .B(new_n946), .C1(new_n953), .C2(new_n954), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n950), .A2(new_n952), .A3(new_n955), .ZN(G57));
endmodule


