//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n545, new_n546, new_n547, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n563, new_n564, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n831, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1181;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AND2_X1   g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  AOI21_X1  g032(.A(new_n457), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n460), .A2(new_n462), .A3(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT65), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(new_n466), .A3(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n464), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n460), .A2(new_n462), .A3(G137), .A4(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G101), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(G2104), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n460), .A2(new_n462), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(new_n471), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n479), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NAND4_X1  g062(.A1(new_n460), .A2(new_n462), .A3(G126), .A4(G2105), .ZN(new_n488));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n489), .A2(new_n491), .A3(G2104), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n460), .A2(new_n462), .A3(G138), .A4(new_n471), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n465), .A2(new_n496), .A3(G138), .A4(new_n471), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n493), .B1(new_n495), .B2(new_n497), .ZN(G164));
  XNOR2_X1  g073(.A(KEYINPUT5), .B(G543), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n499), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT6), .B(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G50), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n501), .A2(KEYINPUT6), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G651), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n507), .A2(new_n509), .A3(new_n510), .A4(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n504), .A2(new_n505), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n502), .A2(new_n515), .ZN(G166));
  NAND3_X1  g091(.A1(new_n499), .A2(new_n503), .A3(G89), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n503), .A2(G51), .A3(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OR2_X1    g094(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AND2_X1   g099(.A1(G63), .A2(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n499), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n523), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n527), .A2(new_n520), .A3(new_n521), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n524), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n519), .A2(new_n529), .ZN(G168));
  AOI22_X1  g105(.A1(new_n499), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n531), .A2(new_n501), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n499), .A2(new_n503), .A3(G90), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n503), .A2(G52), .A3(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n532), .A2(new_n535), .ZN(G171));
  NAND3_X1  g111(.A1(new_n503), .A2(G43), .A3(G543), .ZN(new_n537));
  INV_X1    g112(.A(G81), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n499), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  OAI221_X1 g114(.A(new_n537), .B1(new_n538), .B2(new_n513), .C1(new_n539), .C2(new_n501), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  AND3_X1   g117(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G36), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  XOR2_X1   g122(.A(new_n547), .B(KEYINPUT67), .Z(G188));
  INV_X1    g123(.A(new_n513), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n507), .A2(new_n509), .A3(G65), .ZN(new_n550));
  NAND2_X1  g125(.A1(G78), .A2(G543), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n549), .A2(G91), .B1(new_n552), .B2(G651), .ZN(new_n553));
  INV_X1    g128(.A(G53), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(KEYINPUT68), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n555), .A2(new_n510), .A3(new_n512), .A4(G543), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT9), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT9), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n503), .A2(new_n558), .A3(G543), .A4(new_n555), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n553), .A2(new_n560), .ZN(G299));
  OAI211_X1 g136(.A(new_n534), .B(new_n533), .C1(new_n531), .C2(new_n501), .ZN(G301));
  AND2_X1   g137(.A1(new_n520), .A2(new_n521), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n563), .A2(new_n527), .B1(new_n499), .B2(new_n525), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n564), .A2(new_n524), .A3(new_n517), .A4(new_n518), .ZN(G286));
  INV_X1    g140(.A(G166), .ZN(G303));
  OAI21_X1  g141(.A(G651), .B1(new_n499), .B2(G74), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n499), .A2(new_n503), .A3(G87), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n503), .A2(G49), .A3(G543), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(KEYINPUT69), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT69), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n567), .A2(new_n568), .A3(new_n569), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(G288));
  NAND3_X1  g149(.A1(new_n499), .A2(new_n503), .A3(G86), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n503), .A2(G48), .A3(G543), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n499), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n575), .B(new_n576), .C1(new_n577), .C2(new_n501), .ZN(G305));
  AOI22_X1  g153(.A1(new_n499), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n579), .A2(new_n501), .ZN(new_n580));
  INV_X1    g155(.A(G47), .ZN(new_n581));
  INV_X1    g156(.A(G85), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n504), .A2(new_n581), .B1(new_n513), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  XNOR2_X1  g161(.A(KEYINPUT70), .B(KEYINPUT10), .ZN(new_n587));
  INV_X1    g162(.A(G92), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n513), .B2(new_n588), .ZN(new_n589));
  XOR2_X1   g164(.A(KEYINPUT70), .B(KEYINPUT10), .Z(new_n590));
  NAND4_X1  g165(.A1(new_n590), .A2(G92), .A3(new_n499), .A4(new_n503), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n503), .A2(G54), .A3(G543), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n499), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n594), .B2(new_n501), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n586), .B1(new_n596), .B2(G868), .ZN(G321));
  XOR2_X1   g172(.A(G321), .B(KEYINPUT71), .Z(G284));
  NAND2_X1  g173(.A1(G286), .A2(G868), .ZN(new_n599));
  AND2_X1   g174(.A1(new_n557), .A2(new_n559), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n499), .A2(new_n503), .A3(G91), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n499), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(new_n501), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n599), .B1(new_n604), .B2(G868), .ZN(G297));
  OAI21_X1  g180(.A(new_n599), .B1(new_n604), .B2(G868), .ZN(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n596), .B1(new_n607), .B2(G860), .ZN(G148));
  NOR2_X1   g183(.A1(new_n541), .A2(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n596), .A2(new_n607), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n609), .B1(new_n611), .B2(KEYINPUT72), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(KEYINPUT72), .B2(new_n611), .ZN(G323));
  XOR2_X1   g188(.A(KEYINPUT73), .B(KEYINPUT11), .Z(new_n614));
  XNOR2_X1  g189(.A(G323), .B(new_n614), .ZN(G282));
  INV_X1    g190(.A(new_n474), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n465), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT12), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2100), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT74), .B(KEYINPUT13), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n480), .A2(G123), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n482), .A2(G135), .ZN(new_n623));
  OR2_X1    g198(.A1(G99), .A2(G2105), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n624), .B(G2104), .C1(G111), .C2(new_n471), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n622), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(G2096), .Z(new_n627));
  NAND2_X1  g202(.A1(new_n619), .A2(new_n620), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n621), .A2(new_n627), .A3(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2435), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n633), .A2(KEYINPUT14), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G1341), .B(G1348), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT76), .ZN(new_n643));
  XOR2_X1   g218(.A(G2443), .B(G2446), .Z(new_n644));
  XOR2_X1   g219(.A(new_n643), .B(new_n644), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n639), .A2(new_n640), .A3(new_n645), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(G14), .A3(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2072), .B(G2078), .Z(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT77), .B(KEYINPUT18), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n651), .A2(new_n652), .ZN(new_n658));
  INV_X1    g233(.A(new_n654), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n658), .B1(KEYINPUT17), .B2(new_n659), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n660), .B(new_n653), .C1(KEYINPUT17), .C2(new_n659), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n654), .A2(KEYINPUT78), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n654), .A2(KEYINPUT78), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n662), .A2(new_n658), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n657), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2096), .B(G2100), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT79), .B(KEYINPUT19), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n672), .A2(new_n673), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n671), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n674), .A2(KEYINPUT80), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(KEYINPUT80), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n677), .A2(new_n670), .A3(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n680));
  OAI221_X1 g255(.A(new_n676), .B1(new_n671), .B2(new_n675), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n680), .B2(new_n679), .ZN(new_n682));
  XOR2_X1   g257(.A(G1991), .B(G1996), .Z(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT81), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n682), .B(new_n688), .Z(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G229));
  NAND2_X1  g265(.A1(G162), .A2(G29), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(G29), .B2(G35), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G2090), .ZN(new_n696));
  NAND2_X1  g271(.A1(G115), .A2(G2104), .ZN(new_n697));
  INV_X1    g272(.A(G127), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n479), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G2105), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n482), .A2(G139), .ZN(new_n701));
  INV_X1    g276(.A(G103), .ZN(new_n702));
  OAI21_X1  g277(.A(KEYINPUT25), .B1(new_n474), .B2(new_n702), .ZN(new_n703));
  OR3_X1    g278(.A1(new_n474), .A2(KEYINPUT25), .A3(new_n702), .ZN(new_n704));
  AND4_X1   g279(.A1(new_n700), .A2(new_n701), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT89), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G29), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G29), .B2(G33), .ZN(new_n709));
  INV_X1    g284(.A(G2072), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n695), .A2(new_n696), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G19), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(new_n541), .B2(new_n712), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT85), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G1341), .ZN(new_n716));
  NAND2_X1  g291(.A1(G168), .A2(G16), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G16), .B2(G21), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT92), .B(G1966), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n626), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT31), .B(G11), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT93), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT30), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n722), .B1(new_n726), .B2(G28), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n726), .B2(G28), .ZN(new_n728));
  NOR3_X1   g303(.A1(new_n723), .A2(new_n725), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n718), .A2(new_n720), .ZN(new_n730));
  NAND2_X1  g305(.A1(G171), .A2(G16), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G5), .B2(G16), .ZN(new_n732));
  INV_X1    g307(.A(G1961), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n721), .A2(new_n729), .A3(new_n730), .A4(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(G29), .A2(G32), .ZN(new_n736));
  NAND3_X1  g311(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT26), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G105), .B2(new_n616), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n480), .A2(G129), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n482), .A2(G141), .ZN(new_n741));
  AND3_X1   g316(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n736), .B1(new_n742), .B2(G29), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT27), .B(G1996), .Z(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n733), .B2(new_n732), .ZN(new_n747));
  NOR3_X1   g322(.A1(new_n735), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n712), .A2(G4), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n596), .B2(new_n712), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT84), .B(G1348), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n750), .B(new_n751), .Z(new_n752));
  NOR2_X1   g327(.A1(G27), .A2(G29), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G164), .B2(G29), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G2078), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n711), .A2(new_n716), .A3(new_n748), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n712), .A2(G20), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT95), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT23), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n604), .B2(new_n712), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT96), .B(G1956), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n694), .B2(G2090), .ZN(new_n764));
  AND2_X1   g339(.A1(KEYINPUT24), .A2(G34), .ZN(new_n765));
  NOR2_X1   g340(.A1(KEYINPUT24), .A2(G34), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n722), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT90), .Z(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n477), .B2(new_n722), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT91), .Z(new_n770));
  INV_X1    g345(.A(G2084), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n764), .B(new_n772), .C1(new_n710), .C2(new_n709), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n722), .A2(G26), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT87), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT28), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n480), .A2(G128), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n482), .A2(G140), .ZN(new_n778));
  OR2_X1    g353(.A1(G104), .A2(G2105), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n779), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n777), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT86), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n776), .B1(new_n783), .B2(G29), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT88), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(G2067), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n770), .A2(new_n771), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n785), .A2(G2067), .ZN(new_n789));
  NOR4_X1   g364(.A1(new_n757), .A2(new_n773), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n712), .A2(G6), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n575), .A2(new_n576), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n507), .A2(new_n509), .A3(G61), .ZN(new_n793));
  NAND2_X1  g368(.A1(G73), .A2(G543), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n501), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n791), .B1(new_n796), .B2(new_n712), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT32), .B(G1981), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(G16), .A2(G23), .ZN(new_n800));
  INV_X1    g375(.A(new_n570), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(G16), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT33), .B(G1976), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n799), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n712), .A2(G22), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G166), .B2(new_n712), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1971), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT34), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n722), .A2(G25), .ZN(new_n811));
  OR2_X1    g386(.A1(G95), .A2(G2105), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n812), .B(G2104), .C1(G107), .C2(new_n471), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT82), .ZN(new_n814));
  AOI22_X1  g389(.A1(G119), .A2(new_n480), .B1(new_n482), .B2(G131), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n811), .B1(new_n817), .B2(new_n722), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT35), .B(G1991), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT83), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n818), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n712), .A2(G24), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n584), .B2(new_n712), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(G1986), .Z(new_n824));
  AND2_X1   g399(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n810), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n826), .A2(KEYINPUT36), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n826), .A2(KEYINPUT36), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n790), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(G311));
  INV_X1    g405(.A(KEYINPUT97), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n790), .B(KEYINPUT97), .C1(new_n827), .C2(new_n828), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(G150));
  NAND3_X1  g409(.A1(new_n503), .A2(G55), .A3(G543), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n499), .A2(new_n503), .A3(G93), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n499), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n835), .B(new_n836), .C1(new_n837), .C2(new_n501), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(G860), .ZN(new_n839));
  XOR2_X1   g414(.A(KEYINPUT99), .B(KEYINPUT37), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n596), .A2(G559), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT39), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT98), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n540), .B(new_n838), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(G860), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n845), .B2(new_n847), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n841), .B1(new_n848), .B2(new_n850), .ZN(G145));
  XNOR2_X1  g426(.A(new_n707), .B(new_n618), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n482), .A2(G142), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n471), .A2(G118), .ZN(new_n854));
  OAI21_X1  g429(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(G130), .B2(new_n480), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n783), .B(new_n857), .Z(new_n858));
  AND2_X1   g433(.A1(new_n852), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n852), .A2(new_n858), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n477), .B(new_n626), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n486), .B(G164), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n742), .B(new_n816), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n865), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n861), .A2(new_n868), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n866), .B(new_n867), .C1(new_n859), .C2(new_n860), .ZN(new_n870));
  XNOR2_X1  g445(.A(KEYINPUT100), .B(G37), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g448(.A(KEYINPUT105), .ZN(new_n874));
  XNOR2_X1  g449(.A(G166), .B(G305), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n584), .B(new_n570), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n875), .A2(new_n876), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(KEYINPUT42), .A3(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n881));
  INV_X1    g456(.A(new_n879), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n881), .B1(new_n882), .B2(new_n877), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(new_n596), .B2(G299), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n499), .A2(G66), .ZN(new_n887));
  AND2_X1   g462(.A1(G79), .A2(G543), .ZN(new_n888));
  OAI21_X1  g463(.A(G651), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n889), .A2(new_n593), .A3(new_n591), .A4(new_n589), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n604), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n596), .A2(G299), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n886), .B1(new_n893), .B2(new_n885), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT102), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(KEYINPUT101), .B1(new_n891), .B2(new_n892), .ZN(new_n897));
  OAI21_X1  g472(.A(KEYINPUT102), .B1(new_n897), .B2(new_n886), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n846), .B(new_n610), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n900), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT41), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n893), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n893), .A2(new_n885), .ZN(new_n905));
  INV_X1    g480(.A(new_n886), .ZN(new_n906));
  XNOR2_X1  g481(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n902), .A2(new_n904), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n884), .A2(new_n901), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(KEYINPUT104), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n901), .A2(new_n909), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n912), .A2(new_n880), .A3(new_n883), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT104), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n884), .A2(new_n901), .A3(new_n909), .A4(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n911), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(G868), .ZN(new_n917));
  INV_X1    g492(.A(new_n838), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n918), .A2(G868), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n874), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  AOI211_X1 g496(.A(KEYINPUT105), .B(new_n919), .C1(new_n916), .C2(G868), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(G295));
  NAND2_X1  g498(.A1(new_n917), .A2(new_n920), .ZN(G331));
  INV_X1    g499(.A(new_n907), .ZN(new_n925));
  NOR3_X1   g500(.A1(new_n897), .A2(new_n886), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n904), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT106), .B1(G171), .B2(G286), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT106), .ZN(new_n929));
  NAND3_X1  g504(.A1(G168), .A2(new_n929), .A3(G301), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(G171), .A2(G286), .A3(KEYINPUT107), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(G168), .B2(G301), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n931), .A2(new_n846), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n846), .B1(new_n931), .B2(new_n935), .ZN(new_n937));
  OAI22_X1  g512(.A1(new_n926), .A2(new_n927), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n878), .A2(new_n879), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n931), .A2(new_n935), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n847), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n931), .A2(new_n846), .A3(new_n935), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n941), .B(new_n942), .C1(new_n897), .C2(new_n886), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n938), .A2(new_n939), .A3(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n939), .ZN(new_n946));
  AOI22_X1  g521(.A1(new_n908), .A2(new_n904), .B1(new_n941), .B2(new_n942), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n936), .A2(new_n937), .A3(new_n894), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G37), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n945), .B1(new_n951), .B2(KEYINPUT108), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n949), .A2(new_n953), .A3(new_n950), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT43), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n936), .A2(new_n937), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n899), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n941), .A2(new_n942), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n891), .A2(new_n892), .A3(KEYINPUT41), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(KEYINPUT109), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n925), .B1(new_n897), .B2(new_n886), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n959), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n958), .A2(new_n963), .A3(new_n946), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n944), .A2(new_n871), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT110), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n958), .A2(new_n963), .A3(new_n946), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT110), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n967), .A2(new_n968), .A3(new_n871), .A4(new_n944), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n956), .B1(new_n966), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT44), .B1(new_n955), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n956), .B1(new_n952), .B2(new_n954), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n964), .A2(new_n965), .A3(KEYINPUT43), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n971), .A2(new_n975), .ZN(G397));
  NAND2_X1  g551(.A1(new_n495), .A2(new_n497), .ZN(new_n977));
  INV_X1    g552(.A(new_n493), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(KEYINPUT111), .B(G1384), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n470), .A2(G40), .A3(new_n476), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G2067), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n783), .B(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n742), .B(G1996), .ZN(new_n988));
  OR2_X1    g563(.A1(new_n817), .A2(new_n820), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n817), .A2(new_n820), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n987), .A2(new_n988), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  XOR2_X1   g566(.A(new_n584), .B(G1986), .Z(new_n992));
  OAI21_X1  g567(.A(new_n985), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G40), .ZN(new_n994));
  AOI211_X1 g569(.A(new_n994), .B(new_n475), .C1(new_n469), .C2(G2105), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT50), .ZN(new_n997));
  INV_X1    g572(.A(G1384), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n979), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n995), .A2(new_n996), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G1956), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI211_X1 g577(.A(KEYINPUT116), .B(KEYINPUT57), .C1(new_n600), .C2(new_n603), .ZN(new_n1003));
  OR2_X1    g578(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n1004));
  NAND2_X1  g579(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n553), .A2(new_n560), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n982), .B1(G164), .B2(G1384), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n979), .A2(KEYINPUT45), .A3(new_n980), .ZN(new_n1009));
  XNOR2_X1  g584(.A(KEYINPUT56), .B(G2072), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n995), .A2(new_n1008), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1002), .A2(new_n1007), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT117), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1002), .A2(new_n1011), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1007), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  AOI211_X1 g591(.A(KEYINPUT117), .B(new_n1007), .C1(new_n1002), .C2(new_n1011), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1000), .A2(new_n751), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n979), .A2(new_n998), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n984), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n986), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n890), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1012), .B1(new_n1018), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT61), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1012), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1012), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1007), .B1(new_n1002), .B2(new_n1011), .ZN(new_n1028));
  OAI22_X1  g603(.A1(new_n1027), .A2(new_n1028), .B1(KEYINPUT120), .B2(new_n1025), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1025), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT120), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1031), .B(new_n1025), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1032));
  INV_X1    g607(.A(G1996), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n995), .A2(new_n1008), .A3(new_n1009), .A4(new_n1033), .ZN(new_n1034));
  XOR2_X1   g609(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n1035));
  XNOR2_X1  g610(.A(new_n1035), .B(G1341), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1036), .B1(new_n984), .B2(new_n1020), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1034), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n541), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT119), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1038), .A2(KEYINPUT119), .A3(new_n541), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(KEYINPUT59), .A3(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT119), .B1(new_n1038), .B2(new_n541), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT59), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n751), .A2(new_n1000), .B1(new_n1021), .B2(new_n986), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n890), .A2(KEYINPUT60), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1044), .A2(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1019), .A2(new_n890), .A3(new_n1022), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT60), .B1(new_n1049), .B2(new_n1023), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1032), .A2(new_n1043), .A3(new_n1048), .A4(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1024), .B1(new_n1030), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n1053));
  INV_X1    g628(.A(G2078), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n995), .A2(new_n1008), .A3(new_n1009), .A4(new_n1054), .ZN(new_n1055));
  XOR2_X1   g630(.A(KEYINPUT122), .B(KEYINPUT53), .Z(new_n1056));
  AOI22_X1  g631(.A1(new_n1055), .A2(new_n1056), .B1(new_n1000), .B2(new_n733), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n475), .A2(KEYINPUT123), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n475), .A2(KEYINPUT123), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1054), .A2(KEYINPUT53), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1060), .A2(new_n994), .ZN(new_n1061));
  AND4_X1   g636(.A1(new_n470), .A2(new_n1058), .A3(new_n1059), .A4(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1062), .A2(new_n1009), .A3(new_n983), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1057), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1053), .B1(new_n1064), .B2(G171), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n979), .A2(KEYINPUT45), .A3(new_n998), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n995), .A2(new_n1008), .A3(new_n1066), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n1067), .A2(new_n1060), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1057), .A2(new_n1068), .A3(KEYINPUT124), .A4(G301), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1057), .A2(G301), .A3(new_n1068), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT124), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1065), .A2(new_n1069), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT125), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1065), .A2(new_n1072), .A3(KEYINPUT125), .A4(new_n1069), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G8), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n995), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT112), .B(G1971), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n995), .A2(new_n996), .A3(new_n999), .A4(new_n696), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1078), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(G303), .A2(G8), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT55), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1084), .B(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT113), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1083), .A2(KEYINPUT113), .A3(new_n1086), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(G168), .A2(new_n1078), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT51), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1000), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1096), .A2(new_n771), .B1(new_n1067), .B2(new_n720), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1092), .B(new_n1095), .C1(new_n1097), .C2(new_n1078), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1067), .A2(new_n720), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(G2084), .B2(new_n1000), .ZN(new_n1100));
  OAI211_X1 g675(.A(G8), .B(new_n1094), .C1(new_n1100), .C2(G286), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1091), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1098), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1057), .A2(G301), .A3(new_n1063), .ZN(new_n1104));
  AOI21_X1  g679(.A(G301), .B1(new_n1057), .B2(new_n1068), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1053), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G1981), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT115), .B1(new_n796), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT49), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1109), .B(G1981), .C1(new_n792), .C2(new_n795), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1109), .B1(G305), .B2(G1981), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1108), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(G164), .A2(G1384), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1078), .B1(new_n995), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT49), .B1(new_n796), .B2(new_n1107), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT115), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(G305), .B2(G1981), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1116), .A2(new_n1118), .A3(new_n1110), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1113), .A2(new_n1115), .A3(new_n1119), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT114), .B(G1976), .Z(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT52), .B1(G288), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n801), .A2(G1976), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1115), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  OAI211_X1 g699(.A(G8), .B(new_n1123), .C1(new_n984), .C2(new_n1020), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT52), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1120), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(G8), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1086), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1127), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  AND4_X1   g706(.A1(new_n1090), .A2(new_n1103), .A3(new_n1106), .A4(new_n1131), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1052), .A2(new_n1077), .A3(new_n1132), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1097), .A2(new_n1078), .A3(G286), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1089), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1131), .B(new_n1134), .C1(new_n1135), .C2(new_n1087), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT63), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1090), .A2(KEYINPUT63), .A3(new_n1131), .A4(new_n1134), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1127), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1141), .B1(new_n1086), .B2(new_n1083), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1142), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1103), .A2(KEYINPUT62), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT62), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1098), .A2(new_n1101), .A3(new_n1145), .A4(new_n1102), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1143), .A2(new_n1144), .A3(new_n1105), .A4(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1090), .ZN(new_n1148));
  NOR2_X1   g723(.A1(G288), .A2(G1976), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1120), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1150), .B1(G1981), .B2(G305), .ZN(new_n1151));
  AOI22_X1  g726(.A1(new_n1148), .A2(new_n1141), .B1(new_n1115), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1140), .A2(new_n1147), .A3(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n993), .B1(new_n1133), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n987), .A2(new_n742), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT46), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1155), .A2(new_n985), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n985), .A2(new_n1033), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1159), .B1(KEYINPUT126), .B2(KEYINPUT46), .ZN(new_n1160));
  AOI211_X1 g735(.A(new_n1156), .B(new_n1157), .C1(new_n985), .C2(new_n1033), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1158), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT47), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n987), .A2(new_n988), .ZN(new_n1164));
  OAI22_X1  g739(.A1(new_n1164), .A2(new_n990), .B1(G2067), .B2(new_n783), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(new_n985), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n991), .A2(new_n985), .ZN(new_n1167));
  NOR4_X1   g742(.A1(new_n983), .A2(new_n984), .A3(G290), .A4(G1986), .ZN(new_n1168));
  XOR2_X1   g743(.A(new_n1168), .B(KEYINPUT48), .Z(new_n1169));
  NAND2_X1  g744(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  AND3_X1   g745(.A1(new_n1163), .A2(new_n1166), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1154), .A2(new_n1171), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g747(.A1(new_n973), .A2(new_n974), .ZN(new_n1174));
  AOI211_X1 g748(.A(G227), .B(new_n457), .C1(G567), .C2(new_n454), .ZN(new_n1175));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n1176));
  AND3_X1   g750(.A1(new_n649), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g751(.A(new_n1176), .B1(new_n649), .B2(new_n1175), .ZN(new_n1178));
  OAI211_X1 g752(.A(new_n872), .B(new_n689), .C1(new_n1177), .C2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g753(.A1(new_n1174), .A2(new_n1179), .ZN(G308));
  AND2_X1   g754(.A1(new_n872), .A2(new_n689), .ZN(new_n1181));
  OAI221_X1 g755(.A(new_n1181), .B1(new_n1178), .B2(new_n1177), .C1(new_n973), .C2(new_n974), .ZN(G225));
endmodule


