

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U547 ( .A1(n626), .A2(n510), .ZN(n509) );
  XOR2_X1 U548 ( .A(KEYINPUT27), .B(n625), .Z(n510) );
  AND2_X1 U549 ( .A1(n624), .A2(G1996), .ZN(n611) );
  XNOR2_X1 U550 ( .A(KEYINPUT97), .B(KEYINPUT28), .ZN(n630) );
  XNOR2_X1 U551 ( .A(n631), .B(n630), .ZN(n632) );
  NOR2_X1 U552 ( .A1(n584), .A2(n684), .ZN(n624) );
  NOR2_X1 U553 ( .A1(G164), .A2(G1384), .ZN(n685) );
  NOR2_X2 U554 ( .A1(G2105), .A2(n515), .ZN(n862) );
  NOR2_X1 U555 ( .A1(G651), .A2(n573), .ZN(n771) );
  NOR2_X1 U556 ( .A1(n540), .A2(n539), .ZN(G160) );
  INV_X1 U557 ( .A(G2104), .ZN(n515) );
  NAND2_X1 U558 ( .A1(n862), .A2(G102), .ZN(n511) );
  XNOR2_X1 U559 ( .A(n511), .B(KEYINPUT88), .ZN(n514) );
  NOR2_X1 U560 ( .A1(G2104), .A2(G2105), .ZN(n512) );
  XOR2_X2 U561 ( .A(KEYINPUT17), .B(n512), .Z(n860) );
  NAND2_X1 U562 ( .A1(G138), .A2(n860), .ZN(n513) );
  NAND2_X1 U563 ( .A1(n514), .A2(n513), .ZN(n519) );
  AND2_X1 U564 ( .A1(n515), .A2(G2105), .ZN(n856) );
  NAND2_X1 U565 ( .A1(G126), .A2(n856), .ZN(n517) );
  AND2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n857) );
  NAND2_X1 U567 ( .A1(G114), .A2(n857), .ZN(n516) );
  NAND2_X1 U568 ( .A1(n517), .A2(n516), .ZN(n518) );
  NOR2_X1 U569 ( .A1(n519), .A2(n518), .ZN(G164) );
  INV_X1 U570 ( .A(G651), .ZN(n525) );
  NOR2_X1 U571 ( .A1(G543), .A2(n525), .ZN(n520) );
  XOR2_X1 U572 ( .A(KEYINPUT1), .B(n520), .Z(n775) );
  NAND2_X1 U573 ( .A1(G63), .A2(n775), .ZN(n522) );
  XOR2_X1 U574 ( .A(G543), .B(KEYINPUT0), .Z(n573) );
  NAND2_X1 U575 ( .A1(G51), .A2(n771), .ZN(n521) );
  NAND2_X1 U576 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U577 ( .A(KEYINPUT6), .B(n523), .ZN(n530) );
  NOR2_X1 U578 ( .A1(G651), .A2(G543), .ZN(n772) );
  NAND2_X1 U579 ( .A1(n772), .A2(G89), .ZN(n524) );
  XNOR2_X1 U580 ( .A(n524), .B(KEYINPUT4), .ZN(n527) );
  NOR2_X1 U581 ( .A1(n573), .A2(n525), .ZN(n769) );
  NAND2_X1 U582 ( .A1(G76), .A2(n769), .ZN(n526) );
  NAND2_X1 U583 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U584 ( .A(n528), .B(KEYINPUT5), .Z(n529) );
  NOR2_X1 U585 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U586 ( .A(KEYINPUT76), .B(n531), .Z(n532) );
  XNOR2_X1 U587 ( .A(KEYINPUT7), .B(n532), .ZN(G168) );
  NAND2_X1 U588 ( .A1(G113), .A2(n857), .ZN(n533) );
  XNOR2_X1 U589 ( .A(n533), .B(KEYINPUT64), .ZN(n536) );
  NAND2_X1 U590 ( .A1(G101), .A2(n862), .ZN(n534) );
  XOR2_X1 U591 ( .A(KEYINPUT23), .B(n534), .Z(n535) );
  NAND2_X1 U592 ( .A1(n536), .A2(n535), .ZN(n540) );
  NAND2_X1 U593 ( .A1(G125), .A2(n856), .ZN(n538) );
  NAND2_X1 U594 ( .A1(G137), .A2(n860), .ZN(n537) );
  NAND2_X1 U595 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U596 ( .A1(G64), .A2(n775), .ZN(n542) );
  NAND2_X1 U597 ( .A1(G52), .A2(n771), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n542), .A2(n541), .ZN(n547) );
  NAND2_X1 U599 ( .A1(G90), .A2(n772), .ZN(n544) );
  NAND2_X1 U600 ( .A1(G77), .A2(n769), .ZN(n543) );
  NAND2_X1 U601 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U602 ( .A(KEYINPUT9), .B(n545), .Z(n546) );
  NOR2_X1 U603 ( .A1(n547), .A2(n546), .ZN(G171) );
  NAND2_X1 U604 ( .A1(G53), .A2(n771), .ZN(n548) );
  XNOR2_X1 U605 ( .A(n548), .B(KEYINPUT68), .ZN(n555) );
  NAND2_X1 U606 ( .A1(G65), .A2(n775), .ZN(n550) );
  NAND2_X1 U607 ( .A1(G91), .A2(n772), .ZN(n549) );
  NAND2_X1 U608 ( .A1(n550), .A2(n549), .ZN(n553) );
  NAND2_X1 U609 ( .A1(G78), .A2(n769), .ZN(n551) );
  XNOR2_X1 U610 ( .A(KEYINPUT67), .B(n551), .ZN(n552) );
  NOR2_X1 U611 ( .A1(n553), .A2(n552), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n555), .A2(n554), .ZN(G299) );
  XOR2_X1 U613 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U614 ( .A1(G88), .A2(n772), .ZN(n557) );
  NAND2_X1 U615 ( .A1(G75), .A2(n769), .ZN(n556) );
  NAND2_X1 U616 ( .A1(n557), .A2(n556), .ZN(n560) );
  NAND2_X1 U617 ( .A1(G62), .A2(n775), .ZN(n558) );
  XNOR2_X1 U618 ( .A(KEYINPUT83), .B(n558), .ZN(n559) );
  NOR2_X1 U619 ( .A1(n560), .A2(n559), .ZN(n562) );
  NAND2_X1 U620 ( .A1(n771), .A2(G50), .ZN(n561) );
  NAND2_X1 U621 ( .A1(n562), .A2(n561), .ZN(G303) );
  NAND2_X1 U622 ( .A1(G61), .A2(n775), .ZN(n564) );
  NAND2_X1 U623 ( .A1(G86), .A2(n772), .ZN(n563) );
  NAND2_X1 U624 ( .A1(n564), .A2(n563), .ZN(n567) );
  NAND2_X1 U625 ( .A1(n769), .A2(G73), .ZN(n565) );
  XOR2_X1 U626 ( .A(KEYINPUT2), .B(n565), .Z(n566) );
  NOR2_X1 U627 ( .A1(n567), .A2(n566), .ZN(n569) );
  NAND2_X1 U628 ( .A1(n771), .A2(G48), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n569), .A2(n568), .ZN(G305) );
  NAND2_X1 U630 ( .A1(G49), .A2(n771), .ZN(n571) );
  NAND2_X1 U631 ( .A1(G74), .A2(G651), .ZN(n570) );
  NAND2_X1 U632 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U633 ( .A1(n775), .A2(n572), .ZN(n575) );
  NAND2_X1 U634 ( .A1(n573), .A2(G87), .ZN(n574) );
  NAND2_X1 U635 ( .A1(n575), .A2(n574), .ZN(G288) );
  NAND2_X1 U636 ( .A1(n775), .A2(G60), .ZN(n576) );
  XOR2_X1 U637 ( .A(KEYINPUT65), .B(n576), .Z(n578) );
  NAND2_X1 U638 ( .A1(n771), .A2(G47), .ZN(n577) );
  NAND2_X1 U639 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U640 ( .A(KEYINPUT66), .B(n579), .Z(n583) );
  NAND2_X1 U641 ( .A1(G85), .A2(n772), .ZN(n581) );
  NAND2_X1 U642 ( .A1(G72), .A2(n769), .ZN(n580) );
  AND2_X1 U643 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U644 ( .A1(n583), .A2(n582), .ZN(G290) );
  INV_X1 U645 ( .A(n685), .ZN(n584) );
  NAND2_X1 U646 ( .A1(G160), .A2(G40), .ZN(n684) );
  INV_X1 U647 ( .A(n624), .ZN(n640) );
  NAND2_X1 U648 ( .A1(G8), .A2(n640), .ZN(n672) );
  NOR2_X1 U649 ( .A1(G1966), .A2(n672), .ZN(n653) );
  NOR2_X1 U650 ( .A1(G2084), .A2(n640), .ZN(n650) );
  NOR2_X1 U651 ( .A1(n653), .A2(n650), .ZN(n585) );
  NAND2_X1 U652 ( .A1(G8), .A2(n585), .ZN(n586) );
  XNOR2_X1 U653 ( .A(KEYINPUT30), .B(n586), .ZN(n587) );
  NOR2_X1 U654 ( .A1(G168), .A2(n587), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G1961), .B(KEYINPUT95), .ZN(n972) );
  NAND2_X1 U656 ( .A1(n640), .A2(n972), .ZN(n589) );
  XNOR2_X1 U657 ( .A(G2078), .B(KEYINPUT25), .ZN(n924) );
  NAND2_X1 U658 ( .A1(n624), .A2(n924), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n589), .A2(n588), .ZN(n635) );
  NOR2_X1 U660 ( .A1(G171), .A2(n635), .ZN(n590) );
  NOR2_X1 U661 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U662 ( .A(KEYINPUT31), .B(n592), .Z(n639) );
  NAND2_X1 U663 ( .A1(G66), .A2(n775), .ZN(n594) );
  NAND2_X1 U664 ( .A1(G92), .A2(n772), .ZN(n593) );
  NAND2_X1 U665 ( .A1(n594), .A2(n593), .ZN(n598) );
  NAND2_X1 U666 ( .A1(G54), .A2(n771), .ZN(n596) );
  NAND2_X1 U667 ( .A1(G79), .A2(n769), .ZN(n595) );
  NAND2_X1 U668 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U669 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U670 ( .A(KEYINPUT15), .B(n599), .Z(n600) );
  XOR2_X1 U671 ( .A(KEYINPUT74), .B(n600), .Z(n747) );
  INV_X1 U672 ( .A(n747), .ZN(n939) );
  NAND2_X1 U673 ( .A1(G56), .A2(n775), .ZN(n601) );
  XOR2_X1 U674 ( .A(KEYINPUT14), .B(n601), .Z(n608) );
  NAND2_X1 U675 ( .A1(G81), .A2(n772), .ZN(n602) );
  XOR2_X1 U676 ( .A(KEYINPUT71), .B(n602), .Z(n603) );
  XNOR2_X1 U677 ( .A(n603), .B(KEYINPUT12), .ZN(n605) );
  NAND2_X1 U678 ( .A1(G68), .A2(n769), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U680 ( .A(KEYINPUT13), .B(n606), .Z(n607) );
  NOR2_X1 U681 ( .A1(n608), .A2(n607), .ZN(n610) );
  NAND2_X1 U682 ( .A1(n771), .A2(G43), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n610), .A2(n609), .ZN(n948) );
  XOR2_X1 U684 ( .A(n611), .B(KEYINPUT26), .Z(n613) );
  NAND2_X1 U685 ( .A1(n640), .A2(G1341), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U687 ( .A1(n948), .A2(n614), .ZN(n615) );
  OR2_X1 U688 ( .A1(n939), .A2(n615), .ZN(n622) );
  NAND2_X1 U689 ( .A1(n615), .A2(n939), .ZN(n620) );
  NAND2_X1 U690 ( .A1(n640), .A2(G1348), .ZN(n616) );
  XNOR2_X1 U691 ( .A(n616), .B(KEYINPUT98), .ZN(n618) );
  NAND2_X1 U692 ( .A1(n624), .A2(G2067), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U694 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n622), .A2(n621), .ZN(n628) );
  INV_X1 U696 ( .A(G299), .ZN(n784) );
  NAND2_X1 U697 ( .A1(G1956), .A2(n640), .ZN(n623) );
  XNOR2_X1 U698 ( .A(n623), .B(KEYINPUT96), .ZN(n626) );
  NAND2_X1 U699 ( .A1(n624), .A2(G2072), .ZN(n625) );
  NAND2_X1 U700 ( .A1(n784), .A2(n509), .ZN(n627) );
  NAND2_X1 U701 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U702 ( .A(KEYINPUT99), .B(n629), .ZN(n633) );
  OR2_X1 U703 ( .A1(n509), .A2(n784), .ZN(n631) );
  NOR2_X1 U704 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U705 ( .A(n634), .B(KEYINPUT29), .ZN(n637) );
  NAND2_X1 U706 ( .A1(G171), .A2(n635), .ZN(n636) );
  NAND2_X1 U707 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U708 ( .A1(n639), .A2(n638), .ZN(n651) );
  NAND2_X1 U709 ( .A1(n651), .A2(G286), .ZN(n645) );
  NOR2_X1 U710 ( .A1(G1971), .A2(n672), .ZN(n642) );
  NOR2_X1 U711 ( .A1(G2090), .A2(n640), .ZN(n641) );
  NOR2_X1 U712 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U713 ( .A1(n643), .A2(G303), .ZN(n644) );
  NAND2_X1 U714 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U715 ( .A(KEYINPUT100), .B(n646), .ZN(n647) );
  NAND2_X1 U716 ( .A1(n647), .A2(G8), .ZN(n649) );
  XOR2_X1 U717 ( .A(KEYINPUT32), .B(KEYINPUT101), .Z(n648) );
  XNOR2_X1 U718 ( .A(n649), .B(n648), .ZN(n657) );
  NAND2_X1 U719 ( .A1(G8), .A2(n650), .ZN(n655) );
  INV_X1 U720 ( .A(n651), .ZN(n652) );
  NOR2_X1 U721 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U722 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U723 ( .A1(n657), .A2(n656), .ZN(n667) );
  NOR2_X1 U724 ( .A1(G2090), .A2(G303), .ZN(n658) );
  NAND2_X1 U725 ( .A1(G8), .A2(n658), .ZN(n659) );
  NAND2_X1 U726 ( .A1(n667), .A2(n659), .ZN(n660) );
  NAND2_X1 U727 ( .A1(n660), .A2(n672), .ZN(n683) );
  XNOR2_X1 U728 ( .A(KEYINPUT24), .B(KEYINPUT94), .ZN(n661) );
  XNOR2_X1 U729 ( .A(n661), .B(KEYINPUT93), .ZN(n663) );
  NOR2_X1 U730 ( .A1(G1981), .A2(G305), .ZN(n662) );
  XNOR2_X1 U731 ( .A(n663), .B(n662), .ZN(n664) );
  NOR2_X1 U732 ( .A1(n672), .A2(n664), .ZN(n681) );
  XNOR2_X1 U733 ( .A(G1981), .B(G305), .ZN(n956) );
  NOR2_X1 U734 ( .A1(G1976), .A2(G288), .ZN(n940) );
  NOR2_X1 U735 ( .A1(G1971), .A2(G303), .ZN(n665) );
  NOR2_X1 U736 ( .A1(n940), .A2(n665), .ZN(n666) );
  NAND2_X1 U737 ( .A1(n667), .A2(n666), .ZN(n670) );
  NAND2_X1 U738 ( .A1(G288), .A2(G1976), .ZN(n668) );
  XOR2_X1 U739 ( .A(KEYINPUT102), .B(n668), .Z(n944) );
  NOR2_X1 U740 ( .A1(n672), .A2(n944), .ZN(n669) );
  NAND2_X1 U741 ( .A1(n670), .A2(n669), .ZN(n671) );
  INV_X1 U742 ( .A(KEYINPUT33), .ZN(n675) );
  NAND2_X1 U743 ( .A1(n671), .A2(n675), .ZN(n678) );
  INV_X1 U744 ( .A(n672), .ZN(n673) );
  NAND2_X1 U745 ( .A1(n673), .A2(n940), .ZN(n674) );
  NOR2_X1 U746 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U747 ( .A(n676), .B(KEYINPUT103), .ZN(n677) );
  NAND2_X1 U748 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U749 ( .A1(n956), .A2(n679), .ZN(n680) );
  NOR2_X1 U750 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U751 ( .A1(n683), .A2(n682), .ZN(n718) );
  NOR2_X1 U752 ( .A1(n685), .A2(n684), .ZN(n728) );
  XNOR2_X1 U753 ( .A(G2067), .B(KEYINPUT37), .ZN(n726) );
  NAND2_X1 U754 ( .A1(G128), .A2(n856), .ZN(n687) );
  NAND2_X1 U755 ( .A1(G116), .A2(n857), .ZN(n686) );
  NAND2_X1 U756 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U757 ( .A(n688), .B(KEYINPUT35), .ZN(n693) );
  NAND2_X1 U758 ( .A1(G104), .A2(n862), .ZN(n690) );
  NAND2_X1 U759 ( .A1(G140), .A2(n860), .ZN(n689) );
  NAND2_X1 U760 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U761 ( .A(KEYINPUT34), .B(n691), .Z(n692) );
  NAND2_X1 U762 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U763 ( .A(n694), .B(KEYINPUT36), .Z(n875) );
  OR2_X1 U764 ( .A1(n726), .A2(n875), .ZN(n695) );
  XOR2_X1 U765 ( .A(KEYINPUT90), .B(n695), .Z(n908) );
  NAND2_X1 U766 ( .A1(n728), .A2(n908), .ZN(n724) );
  NAND2_X1 U767 ( .A1(G119), .A2(n856), .ZN(n697) );
  NAND2_X1 U768 ( .A1(G131), .A2(n860), .ZN(n696) );
  NAND2_X1 U769 ( .A1(n697), .A2(n696), .ZN(n700) );
  NAND2_X1 U770 ( .A1(G107), .A2(n857), .ZN(n698) );
  XNOR2_X1 U771 ( .A(KEYINPUT91), .B(n698), .ZN(n699) );
  NOR2_X1 U772 ( .A1(n700), .A2(n699), .ZN(n702) );
  NAND2_X1 U773 ( .A1(n862), .A2(G95), .ZN(n701) );
  NAND2_X1 U774 ( .A1(n702), .A2(n701), .ZN(n870) );
  NAND2_X1 U775 ( .A1(G1991), .A2(n870), .ZN(n711) );
  NAND2_X1 U776 ( .A1(G129), .A2(n856), .ZN(n704) );
  NAND2_X1 U777 ( .A1(G141), .A2(n860), .ZN(n703) );
  NAND2_X1 U778 ( .A1(n704), .A2(n703), .ZN(n707) );
  NAND2_X1 U779 ( .A1(n862), .A2(G105), .ZN(n705) );
  XOR2_X1 U780 ( .A(KEYINPUT38), .B(n705), .Z(n706) );
  NOR2_X1 U781 ( .A1(n707), .A2(n706), .ZN(n709) );
  NAND2_X1 U782 ( .A1(n857), .A2(G117), .ZN(n708) );
  NAND2_X1 U783 ( .A1(n709), .A2(n708), .ZN(n871) );
  NAND2_X1 U784 ( .A1(G1996), .A2(n871), .ZN(n710) );
  NAND2_X1 U785 ( .A1(n711), .A2(n710), .ZN(n904) );
  NAND2_X1 U786 ( .A1(n904), .A2(n728), .ZN(n712) );
  XOR2_X1 U787 ( .A(KEYINPUT92), .B(n712), .Z(n721) );
  INV_X1 U788 ( .A(n721), .ZN(n713) );
  NAND2_X1 U789 ( .A1(n724), .A2(n713), .ZN(n716) );
  XOR2_X1 U790 ( .A(KEYINPUT89), .B(G1986), .Z(n714) );
  XNOR2_X1 U791 ( .A(G290), .B(n714), .ZN(n960) );
  AND2_X1 U792 ( .A1(n960), .A2(n728), .ZN(n715) );
  NOR2_X1 U793 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U794 ( .A1(n718), .A2(n717), .ZN(n731) );
  NOR2_X1 U795 ( .A1(G1996), .A2(n871), .ZN(n897) );
  NOR2_X1 U796 ( .A1(G1986), .A2(G290), .ZN(n719) );
  NOR2_X1 U797 ( .A1(G1991), .A2(n870), .ZN(n895) );
  NOR2_X1 U798 ( .A1(n719), .A2(n895), .ZN(n720) );
  NOR2_X1 U799 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U800 ( .A1(n897), .A2(n722), .ZN(n723) );
  XNOR2_X1 U801 ( .A(n723), .B(KEYINPUT39), .ZN(n725) );
  NAND2_X1 U802 ( .A1(n725), .A2(n724), .ZN(n727) );
  NAND2_X1 U803 ( .A1(n875), .A2(n726), .ZN(n909) );
  NAND2_X1 U804 ( .A1(n727), .A2(n909), .ZN(n729) );
  NAND2_X1 U805 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U806 ( .A1(n731), .A2(n730), .ZN(n733) );
  XNOR2_X1 U807 ( .A(KEYINPUT104), .B(KEYINPUT40), .ZN(n732) );
  XNOR2_X1 U808 ( .A(n733), .B(n732), .ZN(G329) );
  XOR2_X1 U809 ( .A(G2443), .B(G2446), .Z(n735) );
  XNOR2_X1 U810 ( .A(G2427), .B(G2451), .ZN(n734) );
  XNOR2_X1 U811 ( .A(n735), .B(n734), .ZN(n741) );
  XOR2_X1 U812 ( .A(G2430), .B(G2454), .Z(n737) );
  XNOR2_X1 U813 ( .A(G1348), .B(G1341), .ZN(n736) );
  XNOR2_X1 U814 ( .A(n737), .B(n736), .ZN(n739) );
  XOR2_X1 U815 ( .A(G2435), .B(G2438), .Z(n738) );
  XNOR2_X1 U816 ( .A(n739), .B(n738), .ZN(n740) );
  XOR2_X1 U817 ( .A(n741), .B(n740), .Z(n742) );
  AND2_X1 U818 ( .A1(G14), .A2(n742), .ZN(G401) );
  AND2_X1 U819 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U820 ( .A(G57), .ZN(G237) );
  XOR2_X1 U821 ( .A(KEYINPUT11), .B(KEYINPUT70), .Z(n746) );
  XOR2_X1 U822 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n744) );
  NAND2_X1 U823 ( .A1(G7), .A2(G661), .ZN(n743) );
  XOR2_X1 U824 ( .A(n744), .B(n743), .Z(n1004) );
  NAND2_X1 U825 ( .A1(G567), .A2(n1004), .ZN(n745) );
  XNOR2_X1 U826 ( .A(n746), .B(n745), .ZN(G234) );
  XOR2_X1 U827 ( .A(G860), .B(KEYINPUT72), .Z(n753) );
  OR2_X1 U828 ( .A1(n753), .A2(n948), .ZN(G153) );
  XNOR2_X1 U829 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  INV_X1 U830 ( .A(G868), .ZN(n782) );
  NOR2_X1 U831 ( .A1(n782), .A2(G301), .ZN(n749) );
  NOR2_X1 U832 ( .A1(n747), .A2(G868), .ZN(n748) );
  NOR2_X1 U833 ( .A1(n749), .A2(n748), .ZN(n750) );
  XOR2_X1 U834 ( .A(KEYINPUT75), .B(n750), .Z(G284) );
  NAND2_X1 U835 ( .A1(G868), .A2(G286), .ZN(n752) );
  NAND2_X1 U836 ( .A1(G299), .A2(n782), .ZN(n751) );
  NAND2_X1 U837 ( .A1(n752), .A2(n751), .ZN(G297) );
  NAND2_X1 U838 ( .A1(n753), .A2(G559), .ZN(n754) );
  NAND2_X1 U839 ( .A1(n754), .A2(n939), .ZN(n755) );
  XNOR2_X1 U840 ( .A(n755), .B(KEYINPUT77), .ZN(n756) );
  XOR2_X1 U841 ( .A(KEYINPUT16), .B(n756), .Z(G148) );
  NOR2_X1 U842 ( .A1(G868), .A2(n948), .ZN(n759) );
  NAND2_X1 U843 ( .A1(n939), .A2(G868), .ZN(n757) );
  NOR2_X1 U844 ( .A1(G559), .A2(n757), .ZN(n758) );
  NOR2_X1 U845 ( .A1(n759), .A2(n758), .ZN(G282) );
  NAND2_X1 U846 ( .A1(n856), .A2(G123), .ZN(n760) );
  XNOR2_X1 U847 ( .A(n760), .B(KEYINPUT18), .ZN(n762) );
  NAND2_X1 U848 ( .A1(G135), .A2(n860), .ZN(n761) );
  NAND2_X1 U849 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U850 ( .A(KEYINPUT78), .B(n763), .ZN(n767) );
  NAND2_X1 U851 ( .A1(G99), .A2(n862), .ZN(n765) );
  NAND2_X1 U852 ( .A1(G111), .A2(n857), .ZN(n764) );
  NAND2_X1 U853 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U854 ( .A1(n767), .A2(n766), .ZN(n900) );
  XNOR2_X1 U855 ( .A(n900), .B(G2096), .ZN(n768) );
  INV_X1 U856 ( .A(G2100), .ZN(n818) );
  NAND2_X1 U857 ( .A1(n768), .A2(n818), .ZN(G156) );
  NAND2_X1 U858 ( .A1(G80), .A2(n769), .ZN(n770) );
  XNOR2_X1 U859 ( .A(n770), .B(KEYINPUT80), .ZN(n780) );
  NAND2_X1 U860 ( .A1(G55), .A2(n771), .ZN(n774) );
  NAND2_X1 U861 ( .A1(G93), .A2(n772), .ZN(n773) );
  NAND2_X1 U862 ( .A1(n774), .A2(n773), .ZN(n778) );
  NAND2_X1 U863 ( .A1(G67), .A2(n775), .ZN(n776) );
  XNOR2_X1 U864 ( .A(KEYINPUT81), .B(n776), .ZN(n777) );
  NOR2_X1 U865 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U866 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U867 ( .A(KEYINPUT82), .B(n781), .ZN(n1001) );
  NAND2_X1 U868 ( .A1(n782), .A2(n1001), .ZN(n783) );
  XNOR2_X1 U869 ( .A(n783), .B(KEYINPUT84), .ZN(n794) );
  XNOR2_X1 U870 ( .A(n1001), .B(G290), .ZN(n789) );
  XOR2_X1 U871 ( .A(KEYINPUT19), .B(n784), .Z(n785) );
  XNOR2_X1 U872 ( .A(n785), .B(G288), .ZN(n786) );
  XOR2_X1 U873 ( .A(G303), .B(n786), .Z(n787) );
  XNOR2_X1 U874 ( .A(n787), .B(G305), .ZN(n788) );
  XNOR2_X1 U875 ( .A(n789), .B(n788), .ZN(n879) );
  XNOR2_X1 U876 ( .A(n948), .B(KEYINPUT79), .ZN(n791) );
  NAND2_X1 U877 ( .A1(n939), .A2(G559), .ZN(n790) );
  XOR2_X1 U878 ( .A(n791), .B(n790), .Z(n999) );
  XNOR2_X1 U879 ( .A(n879), .B(n999), .ZN(n792) );
  NAND2_X1 U880 ( .A1(G868), .A2(n792), .ZN(n793) );
  NAND2_X1 U881 ( .A1(n794), .A2(n793), .ZN(G295) );
  NAND2_X1 U882 ( .A1(G2078), .A2(G2084), .ZN(n795) );
  XOR2_X1 U883 ( .A(KEYINPUT20), .B(n795), .Z(n796) );
  NAND2_X1 U884 ( .A1(G2090), .A2(n796), .ZN(n797) );
  XNOR2_X1 U885 ( .A(KEYINPUT21), .B(n797), .ZN(n798) );
  NAND2_X1 U886 ( .A1(n798), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U887 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U888 ( .A(KEYINPUT85), .B(KEYINPUT22), .Z(n800) );
  NAND2_X1 U889 ( .A1(G132), .A2(G82), .ZN(n799) );
  XNOR2_X1 U890 ( .A(n800), .B(n799), .ZN(n801) );
  NOR2_X1 U891 ( .A1(n801), .A2(G218), .ZN(n802) );
  NAND2_X1 U892 ( .A1(G96), .A2(n802), .ZN(n1002) );
  NAND2_X1 U893 ( .A1(G2106), .A2(n1002), .ZN(n803) );
  XNOR2_X1 U894 ( .A(n803), .B(KEYINPUT86), .ZN(n807) );
  NAND2_X1 U895 ( .A1(G69), .A2(G120), .ZN(n804) );
  NOR2_X1 U896 ( .A1(G237), .A2(n804), .ZN(n805) );
  NAND2_X1 U897 ( .A1(G108), .A2(n805), .ZN(n1003) );
  NAND2_X1 U898 ( .A1(G567), .A2(n1003), .ZN(n806) );
  NAND2_X1 U899 ( .A1(n807), .A2(n806), .ZN(n884) );
  NAND2_X1 U900 ( .A1(G661), .A2(G483), .ZN(n808) );
  NOR2_X1 U901 ( .A1(n884), .A2(n808), .ZN(n812) );
  NAND2_X1 U902 ( .A1(G36), .A2(n812), .ZN(n809) );
  XOR2_X1 U903 ( .A(KEYINPUT87), .B(n809), .Z(G176) );
  NAND2_X1 U904 ( .A1(G2106), .A2(n1004), .ZN(G217) );
  AND2_X1 U905 ( .A1(G15), .A2(G2), .ZN(n810) );
  NAND2_X1 U906 ( .A1(G661), .A2(n810), .ZN(G259) );
  NAND2_X1 U907 ( .A1(G3), .A2(G1), .ZN(n811) );
  NAND2_X1 U908 ( .A1(n812), .A2(n811), .ZN(G188) );
  XNOR2_X1 U909 ( .A(G96), .B(KEYINPUT105), .ZN(G221) );
  XOR2_X1 U910 ( .A(G2678), .B(G2084), .Z(n814) );
  XNOR2_X1 U911 ( .A(G2067), .B(G2078), .ZN(n813) );
  XNOR2_X1 U912 ( .A(n814), .B(n813), .ZN(n815) );
  XOR2_X1 U913 ( .A(n815), .B(KEYINPUT107), .Z(n817) );
  XNOR2_X1 U914 ( .A(G2072), .B(KEYINPUT42), .ZN(n816) );
  XNOR2_X1 U915 ( .A(n817), .B(n816), .ZN(n822) );
  XNOR2_X1 U916 ( .A(n818), .B(G2096), .ZN(n820) );
  XNOR2_X1 U917 ( .A(G2090), .B(KEYINPUT43), .ZN(n819) );
  XNOR2_X1 U918 ( .A(n820), .B(n819), .ZN(n821) );
  XOR2_X1 U919 ( .A(n822), .B(n821), .Z(G227) );
  XOR2_X1 U920 ( .A(KEYINPUT109), .B(KEYINPUT108), .Z(n824) );
  XNOR2_X1 U921 ( .A(G1966), .B(G1961), .ZN(n823) );
  XNOR2_X1 U922 ( .A(n824), .B(n823), .ZN(n835) );
  INV_X1 U923 ( .A(G1996), .ZN(n825) );
  XNOR2_X1 U924 ( .A(KEYINPUT110), .B(n825), .ZN(n827) );
  XNOR2_X1 U925 ( .A(G1986), .B(G1991), .ZN(n826) );
  XNOR2_X1 U926 ( .A(n827), .B(n826), .ZN(n831) );
  XOR2_X1 U927 ( .A(G1976), .B(G1981), .Z(n829) );
  XNOR2_X1 U928 ( .A(G1956), .B(G1971), .ZN(n828) );
  XNOR2_X1 U929 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U930 ( .A(n831), .B(n830), .Z(n833) );
  XNOR2_X1 U931 ( .A(G2474), .B(KEYINPUT41), .ZN(n832) );
  XNOR2_X1 U932 ( .A(n833), .B(n832), .ZN(n834) );
  XNOR2_X1 U933 ( .A(n835), .B(n834), .ZN(G229) );
  NAND2_X1 U934 ( .A1(G124), .A2(n856), .ZN(n836) );
  XOR2_X1 U935 ( .A(KEYINPUT111), .B(n836), .Z(n837) );
  XNOR2_X1 U936 ( .A(n837), .B(KEYINPUT44), .ZN(n839) );
  NAND2_X1 U937 ( .A1(G100), .A2(n862), .ZN(n838) );
  NAND2_X1 U938 ( .A1(n839), .A2(n838), .ZN(n843) );
  NAND2_X1 U939 ( .A1(G136), .A2(n860), .ZN(n841) );
  NAND2_X1 U940 ( .A1(G112), .A2(n857), .ZN(n840) );
  NAND2_X1 U941 ( .A1(n841), .A2(n840), .ZN(n842) );
  NOR2_X1 U942 ( .A1(n843), .A2(n842), .ZN(G162) );
  XOR2_X1 U943 ( .A(KEYINPUT114), .B(KEYINPUT113), .Z(n845) );
  XNOR2_X1 U944 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U946 ( .A(n846), .B(G162), .Z(n855) );
  NAND2_X1 U947 ( .A1(G103), .A2(n862), .ZN(n848) );
  NAND2_X1 U948 ( .A1(G139), .A2(n860), .ZN(n847) );
  NAND2_X1 U949 ( .A1(n848), .A2(n847), .ZN(n853) );
  NAND2_X1 U950 ( .A1(G127), .A2(n856), .ZN(n850) );
  NAND2_X1 U951 ( .A1(G115), .A2(n857), .ZN(n849) );
  NAND2_X1 U952 ( .A1(n850), .A2(n849), .ZN(n851) );
  XOR2_X1 U953 ( .A(KEYINPUT47), .B(n851), .Z(n852) );
  NOR2_X1 U954 ( .A1(n853), .A2(n852), .ZN(n890) );
  XNOR2_X1 U955 ( .A(n890), .B(n900), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(n869) );
  NAND2_X1 U957 ( .A1(G130), .A2(n856), .ZN(n859) );
  NAND2_X1 U958 ( .A1(G118), .A2(n857), .ZN(n858) );
  NAND2_X1 U959 ( .A1(n859), .A2(n858), .ZN(n867) );
  NAND2_X1 U960 ( .A1(n860), .A2(G142), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n861), .B(KEYINPUT112), .ZN(n864) );
  NAND2_X1 U962 ( .A1(G106), .A2(n862), .ZN(n863) );
  NAND2_X1 U963 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U964 ( .A(n865), .B(KEYINPUT45), .Z(n866) );
  NOR2_X1 U965 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U966 ( .A(n869), .B(n868), .Z(n874) );
  XNOR2_X1 U967 ( .A(G160), .B(n870), .ZN(n872) );
  XNOR2_X1 U968 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U969 ( .A(n874), .B(n873), .Z(n877) );
  XOR2_X1 U970 ( .A(G164), .B(n875), .Z(n876) );
  XNOR2_X1 U971 ( .A(n877), .B(n876), .ZN(n878) );
  NOR2_X1 U972 ( .A1(G37), .A2(n878), .ZN(G395) );
  XNOR2_X1 U973 ( .A(G286), .B(n879), .ZN(n881) );
  XOR2_X1 U974 ( .A(G171), .B(n939), .Z(n880) );
  XNOR2_X1 U975 ( .A(n881), .B(n880), .ZN(n882) );
  XNOR2_X1 U976 ( .A(n882), .B(n948), .ZN(n883) );
  NOR2_X1 U977 ( .A1(G37), .A2(n883), .ZN(G397) );
  XOR2_X1 U978 ( .A(KEYINPUT106), .B(n884), .Z(G319) );
  NOR2_X1 U979 ( .A1(G227), .A2(G229), .ZN(n885) );
  XNOR2_X1 U980 ( .A(KEYINPUT49), .B(n885), .ZN(n886) );
  NOR2_X1 U981 ( .A1(G401), .A2(n886), .ZN(n888) );
  NOR2_X1 U982 ( .A1(G395), .A2(G397), .ZN(n887) );
  AND2_X1 U983 ( .A1(n888), .A2(n887), .ZN(n889) );
  NAND2_X1 U984 ( .A1(n889), .A2(G319), .ZN(G225) );
  XNOR2_X1 U985 ( .A(KEYINPUT115), .B(G225), .ZN(G308) );
  INV_X1 U987 ( .A(KEYINPUT55), .ZN(n913) );
  XOR2_X1 U988 ( .A(G2072), .B(n890), .Z(n892) );
  XOR2_X1 U989 ( .A(G164), .B(G2078), .Z(n891) );
  NOR2_X1 U990 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U991 ( .A(KEYINPUT50), .B(n893), .ZN(n906) );
  XOR2_X1 U992 ( .A(G2084), .B(G160), .Z(n894) );
  NOR2_X1 U993 ( .A1(n895), .A2(n894), .ZN(n902) );
  XOR2_X1 U994 ( .A(G2090), .B(G162), .Z(n896) );
  NOR2_X1 U995 ( .A1(n897), .A2(n896), .ZN(n898) );
  XNOR2_X1 U996 ( .A(n898), .B(KEYINPUT51), .ZN(n899) );
  NOR2_X1 U997 ( .A1(n900), .A2(n899), .ZN(n901) );
  NAND2_X1 U998 ( .A1(n902), .A2(n901), .ZN(n903) );
  NOR2_X1 U999 ( .A1(n904), .A2(n903), .ZN(n905) );
  NAND2_X1 U1000 ( .A1(n906), .A2(n905), .ZN(n907) );
  NOR2_X1 U1001 ( .A1(n908), .A2(n907), .ZN(n910) );
  NAND2_X1 U1002 ( .A1(n910), .A2(n909), .ZN(n911) );
  XOR2_X1 U1003 ( .A(KEYINPUT52), .B(n911), .Z(n912) );
  NAND2_X1 U1004 ( .A1(n913), .A2(n912), .ZN(n914) );
  NAND2_X1 U1005 ( .A1(n914), .A2(G29), .ZN(n997) );
  XNOR2_X1 U1006 ( .A(G2090), .B(G35), .ZN(n930) );
  XOR2_X1 U1007 ( .A(G1991), .B(G25), .Z(n915) );
  XNOR2_X1 U1008 ( .A(KEYINPUT116), .B(n915), .ZN(n916) );
  NAND2_X1 U1009 ( .A1(n916), .A2(G28), .ZN(n917) );
  XNOR2_X1 U1010 ( .A(n917), .B(KEYINPUT117), .ZN(n923) );
  XOR2_X1 U1011 ( .A(G32), .B(G1996), .Z(n919) );
  XOR2_X1 U1012 ( .A(G2072), .B(G33), .Z(n918) );
  NAND2_X1 U1013 ( .A1(n919), .A2(n918), .ZN(n921) );
  XNOR2_X1 U1014 ( .A(G26), .B(G2067), .ZN(n920) );
  NOR2_X1 U1015 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1016 ( .A1(n923), .A2(n922), .ZN(n927) );
  XOR2_X1 U1017 ( .A(G27), .B(n924), .Z(n925) );
  XNOR2_X1 U1018 ( .A(KEYINPUT118), .B(n925), .ZN(n926) );
  NOR2_X1 U1019 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1020 ( .A(KEYINPUT53), .B(n928), .ZN(n929) );
  NOR2_X1 U1021 ( .A1(n930), .A2(n929), .ZN(n933) );
  XOR2_X1 U1022 ( .A(G2084), .B(G34), .Z(n931) );
  XNOR2_X1 U1023 ( .A(KEYINPUT54), .B(n931), .ZN(n932) );
  NAND2_X1 U1024 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1025 ( .A(KEYINPUT55), .B(n934), .Z(n936) );
  INV_X1 U1026 ( .A(G29), .ZN(n935) );
  NAND2_X1 U1027 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1028 ( .A1(G11), .A2(n937), .ZN(n995) );
  INV_X1 U1029 ( .A(G16), .ZN(n991) );
  XOR2_X1 U1030 ( .A(n991), .B(KEYINPUT56), .Z(n964) );
  XOR2_X1 U1031 ( .A(G1956), .B(G299), .Z(n938) );
  XNOR2_X1 U1032 ( .A(n938), .B(KEYINPUT120), .ZN(n946) );
  XNOR2_X1 U1033 ( .A(G1348), .B(n939), .ZN(n942) );
  XNOR2_X1 U1034 ( .A(n940), .B(KEYINPUT121), .ZN(n941) );
  NAND2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1036 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1037 ( .A1(n946), .A2(n945), .ZN(n954) );
  XOR2_X1 U1038 ( .A(G1971), .B(G303), .Z(n947) );
  XNOR2_X1 U1039 ( .A(n947), .B(KEYINPUT122), .ZN(n952) );
  XOR2_X1 U1040 ( .A(G171), .B(G1961), .Z(n950) );
  XNOR2_X1 U1041 ( .A(n948), .B(G1341), .ZN(n949) );
  NOR2_X1 U1042 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1043 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1044 ( .A1(n954), .A2(n953), .ZN(n962) );
  XOR2_X1 U1045 ( .A(G168), .B(G1966), .Z(n955) );
  NOR2_X1 U1046 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1047 ( .A(KEYINPUT119), .B(n957), .Z(n958) );
  XNOR2_X1 U1048 ( .A(n958), .B(KEYINPUT57), .ZN(n959) );
  NOR2_X1 U1049 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1050 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1051 ( .A1(n964), .A2(n963), .ZN(n993) );
  XOR2_X1 U1052 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n971) );
  XNOR2_X1 U1053 ( .A(G1971), .B(G22), .ZN(n966) );
  XNOR2_X1 U1054 ( .A(G23), .B(G1976), .ZN(n965) );
  NOR2_X1 U1055 ( .A1(n966), .A2(n965), .ZN(n969) );
  XOR2_X1 U1056 ( .A(G1986), .B(KEYINPUT124), .Z(n967) );
  XNOR2_X1 U1057 ( .A(G24), .B(n967), .ZN(n968) );
  NAND2_X1 U1058 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1059 ( .A(n971), .B(n970), .ZN(n987) );
  XNOR2_X1 U1060 ( .A(G5), .B(n972), .ZN(n985) );
  XOR2_X1 U1061 ( .A(G1348), .B(KEYINPUT59), .Z(n973) );
  XNOR2_X1 U1062 ( .A(G4), .B(n973), .ZN(n980) );
  XOR2_X1 U1063 ( .A(G1981), .B(G6), .Z(n977) );
  XNOR2_X1 U1064 ( .A(G1956), .B(G20), .ZN(n975) );
  XNOR2_X1 U1065 ( .A(G1341), .B(G19), .ZN(n974) );
  NOR2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1068 ( .A(KEYINPUT123), .B(n978), .Z(n979) );
  NOR2_X1 U1069 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1070 ( .A(KEYINPUT60), .B(n981), .Z(n983) );
  XNOR2_X1 U1071 ( .A(G1966), .B(G21), .ZN(n982) );
  NOR2_X1 U1072 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1073 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1074 ( .A1(n987), .A2(n986), .ZN(n989) );
  XNOR2_X1 U1075 ( .A(KEYINPUT126), .B(KEYINPUT61), .ZN(n988) );
  XNOR2_X1 U1076 ( .A(n989), .B(n988), .ZN(n990) );
  NAND2_X1 U1077 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1078 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1079 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1080 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1081 ( .A(KEYINPUT62), .B(n998), .Z(G311) );
  XNOR2_X1 U1082 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  NOR2_X1 U1083 ( .A1(G860), .A2(n999), .ZN(n1000) );
  XOR2_X1 U1084 ( .A(n1001), .B(n1000), .Z(G145) );
  INV_X1 U1085 ( .A(G132), .ZN(G219) );
  INV_X1 U1086 ( .A(G120), .ZN(G236) );
  INV_X1 U1087 ( .A(G82), .ZN(G220) );
  INV_X1 U1088 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1089 ( .A1(n1003), .A2(n1002), .ZN(G325) );
  INV_X1 U1090 ( .A(G325), .ZN(G261) );
  INV_X1 U1091 ( .A(G108), .ZN(G238) );
  INV_X1 U1092 ( .A(n1004), .ZN(G223) );
  INV_X1 U1093 ( .A(G303), .ZN(G166) );
endmodule

