//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 0 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 1 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n795, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n997, new_n998;
  INV_X1    g000(.A(KEYINPUT107), .ZN(new_n202));
  XOR2_X1   g001(.A(G15gat), .B(G43gat), .Z(new_n203));
  XNOR2_X1  g002(.A(G71gat), .B(G99gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G227gat), .ZN(new_n206));
  INV_X1    g005(.A(G233gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G190gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT68), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT68), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G190gat), .ZN(new_n213));
  AOI21_X1  g012(.A(G183gat), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT24), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT23), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT67), .B(KEYINPUT23), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n221), .B(new_n223), .C1(new_n224), .C2(new_n222), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT25), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n227), .A2(KEYINPUT67), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n227), .A2(KEYINPUT67), .ZN(new_n229));
  OAI22_X1  g028(.A1(new_n228), .A2(new_n229), .B1(G169gat), .B2(G176gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT25), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n221), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT66), .B(G176gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n227), .A2(G169gat), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n217), .A2(KEYINPUT65), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n215), .A2(new_n237), .A3(new_n216), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT64), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n218), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n236), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  OAI22_X1  g040(.A1(new_n218), .A2(new_n239), .B1(G183gat), .B2(G190gat), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n230), .B(new_n235), .C1(new_n241), .C2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT28), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n244), .A2(KEYINPUT69), .ZN(new_n245));
  AND2_X1   g044(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT68), .B(G190gat), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n245), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n211), .A2(new_n213), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT27), .B(G183gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT26), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n222), .A2(new_n258), .ZN(new_n259));
  OAI211_X1 g058(.A(KEYINPUT70), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n257), .A2(new_n221), .A3(new_n259), .A4(new_n260), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n250), .A2(new_n254), .A3(new_n261), .A4(new_n215), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n226), .A2(new_n243), .A3(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(G127gat), .A2(G134gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT71), .B(G127gat), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n264), .B1(new_n265), .B2(G134gat), .ZN(new_n266));
  INV_X1    g065(.A(G113gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G120gat), .ZN(new_n268));
  INV_X1    g067(.A(G120gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(G113gat), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n268), .A2(new_n270), .A3(KEYINPUT72), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT72), .B1(new_n268), .B2(new_n270), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n266), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT73), .B(G120gat), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n268), .B1(new_n276), .B2(new_n267), .ZN(new_n277));
  INV_X1    g076(.A(new_n264), .ZN(new_n278));
  NAND2_X1  g077(.A1(G127gat), .A2(G134gat), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT1), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n263), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n270), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n286), .A2(new_n272), .A3(new_n271), .ZN(new_n287));
  AOI22_X1  g086(.A1(new_n287), .A2(new_n266), .B1(new_n277), .B2(new_n280), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n288), .A2(new_n243), .A3(new_n226), .A4(new_n262), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n209), .B1(new_n283), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT32), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n291), .A2(KEYINPUT33), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n205), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT74), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT74), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n295), .B(new_n205), .C1(new_n290), .C2(new_n292), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n290), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n291), .B1(new_n205), .B2(KEYINPUT33), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(KEYINPUT75), .B(KEYINPUT34), .Z(new_n302));
  NAND2_X1  g101(.A1(new_n283), .A2(new_n289), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n302), .B1(new_n303), .B2(new_n208), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n283), .A2(new_n209), .A3(new_n289), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n304), .B(KEYINPUT76), .C1(KEYINPUT34), .C2(new_n305), .ZN(new_n306));
  OR2_X1    g105(.A1(new_n304), .A2(KEYINPUT76), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n301), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT77), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n294), .A2(new_n296), .B1(new_n298), .B2(new_n299), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(new_n306), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n308), .A2(new_n309), .A3(new_n312), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n301), .A2(KEYINPUT77), .A3(new_n306), .A4(new_n307), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT29), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n263), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G226gat), .A2(G233gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n263), .A2(G226gat), .A3(G233gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT79), .ZN(new_n322));
  INV_X1    g121(.A(G211gat), .ZN(new_n323));
  INV_X1    g122(.A(G218gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G211gat), .A2(G218gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT78), .ZN(new_n328));
  INV_X1    g127(.A(G197gat), .ZN(new_n329));
  INV_X1    g128(.A(G204gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(G197gat), .A2(G204gat), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT22), .ZN(new_n333));
  AOI22_X1  g132(.A1(new_n331), .A2(new_n332), .B1(new_n333), .B2(new_n326), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT78), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n325), .A2(new_n335), .A3(new_n326), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n328), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n334), .B1(new_n328), .B2(new_n336), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n322), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n334), .ZN(new_n340));
  INV_X1    g139(.A(new_n336), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n335), .B1(new_n325), .B2(new_n326), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n328), .A2(new_n334), .A3(new_n336), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n343), .A2(KEYINPUT79), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n339), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n321), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT80), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n348), .B1(new_n317), .B2(new_n318), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n263), .A2(G226gat), .A3(G233gat), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n263), .A2(new_n316), .B1(G226gat), .B2(G233gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n350), .B1(new_n353), .B2(KEYINPUT80), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n347), .B1(new_n354), .B2(new_n346), .ZN(new_n355));
  XNOR2_X1  g154(.A(G8gat), .B(G36gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(G64gat), .B(G92gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n346), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n353), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n349), .B1(new_n321), .B2(new_n348), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n362), .B1(new_n363), .B2(new_n361), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n358), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n360), .A2(new_n365), .A3(KEYINPUT30), .ZN(new_n366));
  OR3_X1    g165(.A1(new_n364), .A2(KEYINPUT30), .A3(new_n358), .ZN(new_n367));
  NAND2_X1  g166(.A1(G225gat), .A2(G233gat), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G141gat), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT84), .B1(new_n370), .B2(G148gat), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT84), .ZN(new_n372));
  INV_X1    g171(.A(G148gat), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(new_n373), .A3(G141gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n370), .A2(G148gat), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n371), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(G155gat), .A2(G162gat), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT85), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(new_n378), .A3(KEYINPUT2), .ZN(new_n379));
  XNOR2_X1  g178(.A(G155gat), .B(G162gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n377), .A2(KEYINPUT2), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT85), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n376), .A2(new_n379), .A3(new_n380), .A4(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT83), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n377), .A2(KEYINPUT83), .A3(KEYINPUT2), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n373), .A2(G141gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n375), .A2(new_n387), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n385), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT82), .ZN(new_n390));
  INV_X1    g189(.A(G155gat), .ZN(new_n391));
  INV_X1    g190(.A(G162gat), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT82), .B1(G155gat), .B2(G162gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT81), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n377), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(KEYINPUT81), .A2(G155gat), .A3(G162gat), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n395), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n383), .B1(new_n389), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT86), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n385), .A2(new_n386), .A3(new_n388), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n403), .A2(new_n395), .A3(new_n397), .A4(new_n398), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n404), .A2(KEYINPUT86), .A3(new_n383), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n288), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n404), .A2(new_n275), .A3(new_n383), .A4(new_n281), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n369), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n407), .A2(KEYINPUT4), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT4), .ZN(new_n411));
  INV_X1    g210(.A(new_n399), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n382), .A2(new_n379), .A3(new_n380), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n412), .A2(new_n403), .B1(new_n413), .B2(new_n376), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n411), .B1(new_n414), .B2(new_n288), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n368), .B1(new_n410), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n282), .B1(new_n400), .B2(KEYINPUT3), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n405), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n417), .B1(new_n418), .B2(KEYINPUT3), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n409), .B(KEYINPUT5), .C1(new_n416), .C2(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n400), .A2(new_n401), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT86), .B1(new_n404), .B2(new_n383), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT3), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n417), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT87), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n426), .B1(new_n407), .B2(KEYINPUT4), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n414), .A2(new_n288), .A3(KEYINPUT87), .A4(new_n411), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n407), .A2(KEYINPUT4), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n369), .A2(KEYINPUT5), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n425), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n420), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(G1gat), .B(G29gat), .ZN(new_n434));
  INV_X1    g233(.A(G85gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(KEYINPUT0), .B(G57gat), .ZN(new_n437));
  XOR2_X1   g236(.A(new_n436), .B(new_n437), .Z(new_n438));
  NAND3_X1  g237(.A1(new_n433), .A2(KEYINPUT6), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n433), .A2(new_n438), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT6), .ZN(new_n441));
  INV_X1    g240(.A(new_n438), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n420), .A2(new_n432), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n440), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n366), .A2(new_n367), .B1(new_n439), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(G228gat), .A2(G233gat), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n343), .A2(new_n316), .A3(new_n344), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT3), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n400), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n316), .B1(new_n400), .B2(KEYINPUT3), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n451), .A2(KEYINPUT88), .B1(new_n346), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT88), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n450), .A2(new_n454), .A3(new_n400), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n447), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n446), .B1(new_n346), .B2(new_n452), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n418), .A2(new_n450), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(G22gat), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n451), .A2(KEYINPUT88), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n346), .A2(new_n452), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n455), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n446), .ZN(new_n464));
  INV_X1    g263(.A(G22gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n457), .A2(new_n458), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n460), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n459), .B1(new_n446), .B2(new_n463), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT89), .B1(new_n469), .B2(new_n465), .ZN(new_n470));
  XNOR2_X1  g269(.A(G78gat), .B(G106gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(KEYINPUT31), .B(G50gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n471), .B(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n468), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n460), .A2(new_n467), .A3(KEYINPUT89), .A4(new_n473), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n315), .A2(new_n445), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT35), .ZN(new_n479));
  AND2_X1   g278(.A1(new_n308), .A2(new_n312), .ZN(new_n480));
  XNOR2_X1  g279(.A(KEYINPUT95), .B(KEYINPUT35), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n480), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n445), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n480), .A2(KEYINPUT36), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT36), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n486), .B1(new_n313), .B2(new_n314), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT90), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT89), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n467), .A2(new_n489), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n490), .A2(new_n473), .B1(new_n467), .B2(new_n460), .ZN(new_n491));
  AND4_X1   g290(.A1(KEYINPUT89), .A2(new_n460), .A3(new_n467), .A4(new_n473), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n488), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n475), .A2(KEYINPUT90), .A3(new_n476), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI22_X1  g294(.A1(new_n485), .A2(new_n487), .B1(new_n495), .B2(new_n445), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT38), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT37), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n359), .B1(new_n355), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n364), .A2(KEYINPUT37), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n497), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n498), .B(new_n362), .C1(new_n363), .C2(new_n361), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n498), .B1(new_n353), .B2(new_n346), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n503), .B1(new_n363), .B2(new_n346), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n502), .A2(new_n504), .A3(new_n497), .A4(new_n358), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n444), .A2(new_n505), .A3(new_n439), .A4(new_n360), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n501), .B1(new_n506), .B2(KEYINPUT93), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n443), .A2(new_n441), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n442), .B1(new_n420), .B2(new_n432), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n439), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT93), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n512), .A2(new_n513), .A3(new_n360), .A4(new_n505), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n507), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n491), .A2(new_n492), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT92), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT40), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n425), .A2(new_n430), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT91), .B(KEYINPUT39), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(new_n369), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n442), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n368), .B1(new_n425), .B2(new_n430), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n418), .A2(new_n282), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n524), .A2(new_n407), .A3(new_n368), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT39), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n517), .B(new_n518), .C1(new_n522), .C2(new_n527), .ZN(new_n528));
  OR2_X1    g327(.A1(new_n523), .A2(new_n526), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n529), .A2(KEYINPUT40), .A3(new_n442), .A4(new_n521), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(new_n530), .A3(new_n440), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n529), .A2(new_n442), .A3(new_n521), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n517), .B1(new_n532), .B2(new_n518), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n366), .A2(new_n367), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n516), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n515), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n496), .B1(KEYINPUT94), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT94), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n515), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n484), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT103), .ZN(new_n542));
  XNOR2_X1  g341(.A(G15gat), .B(G22gat), .ZN(new_n543));
  INV_X1    g342(.A(G1gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT16), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n546), .B1(G1gat), .B2(new_n543), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n547), .A2(G8gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(G8gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AND2_X1   g349(.A1(G71gat), .A2(G78gat), .ZN(new_n551));
  NOR2_X1   g350(.A1(G71gat), .A2(G78gat), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(G57gat), .ZN(new_n554));
  INV_X1    g353(.A(G64gat), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n553), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n551), .B1(KEYINPUT9), .B2(new_n552), .ZN(new_n559));
  NAND2_X1  g358(.A1(KEYINPUT99), .A2(G57gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(new_n555), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n558), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT21), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n550), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n562), .B(KEYINPUT21), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n565), .B1(new_n550), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G231gat), .A2(G233gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(G183gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(new_n323), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n567), .B(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(G127gat), .B(G155gat), .Z(new_n572));
  XOR2_X1   g371(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n571), .A2(new_n574), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT17), .ZN(new_n579));
  XNOR2_X1  g378(.A(G43gat), .B(G50gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT15), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(G29gat), .A2(G36gat), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT14), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n580), .A2(KEYINPUT15), .ZN(new_n587));
  XNOR2_X1  g386(.A(KEYINPUT97), .B(G36gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(G29gat), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n583), .A2(new_n586), .A3(new_n587), .A4(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  AOI211_X1 g390(.A(new_n582), .B(new_n581), .C1(new_n586), .C2(new_n589), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n579), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n583), .A2(new_n586), .A3(new_n589), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n594), .A2(KEYINPUT15), .A3(new_n580), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n595), .A2(KEYINPUT17), .A3(new_n590), .ZN(new_n596));
  NAND2_X1  g395(.A1(G99gat), .A2(G106gat), .ZN(new_n597));
  INV_X1    g396(.A(G92gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(KEYINPUT8), .A2(new_n597), .B1(new_n435), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT7), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n600), .B1(new_n435), .B2(new_n598), .ZN(new_n601));
  NAND3_X1  g400(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(G99gat), .B(G106gat), .Z(new_n604));
  NAND3_X1  g403(.A1(new_n603), .A2(KEYINPUT101), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n604), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n599), .A2(new_n606), .A3(new_n601), .A4(new_n602), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT101), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n603), .A2(new_n604), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n593), .A2(new_n596), .A3(new_n605), .A4(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n590), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n605), .ZN(new_n613));
  NAND2_X1  g412(.A1(G232gat), .A2(G233gat), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n612), .A2(new_n613), .B1(KEYINPUT41), .B2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G190gat), .B(G218gat), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AND3_X1   g417(.A1(new_n611), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n618), .B1(new_n611), .B2(new_n616), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n615), .A2(KEYINPUT41), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(new_n392), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT100), .B(G134gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT102), .ZN(new_n625));
  OR3_X1    g424(.A1(new_n619), .A2(new_n620), .A3(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n624), .A2(KEYINPUT102), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n625), .B(new_n627), .C1(new_n619), .C2(new_n620), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n542), .B1(new_n578), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n577), .A2(KEYINPUT103), .A3(new_n629), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G230gat), .A2(G233gat), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n562), .B1(new_n604), .B2(new_n603), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT104), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n637), .A2(new_n638), .A3(new_n607), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n610), .A2(new_n562), .A3(new_n605), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n561), .A2(new_n559), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n607), .A2(new_n641), .A3(new_n558), .A4(new_n609), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT104), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT10), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n639), .A2(new_n640), .A3(new_n643), .A4(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n613), .A2(KEYINPUT10), .A3(new_n558), .A4(new_n641), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n636), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT105), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI211_X1 g448(.A(KEYINPUT105), .B(new_n636), .C1(new_n645), .C2(new_n646), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n639), .A2(new_n640), .A3(new_n643), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n636), .ZN(new_n653));
  OR2_X1    g452(.A1(new_n653), .A2(KEYINPUT106), .ZN(new_n654));
  XNOR2_X1  g453(.A(G120gat), .B(G148gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n653), .A2(KEYINPUT106), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n654), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n651), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n653), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n657), .B1(new_n662), .B2(new_n647), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n612), .A2(new_n550), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n595), .A2(new_n548), .A3(new_n549), .A4(new_n590), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(G229gat), .A2(G233gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT13), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT98), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n548), .A2(new_n549), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n675), .A2(new_n596), .A3(new_n593), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n676), .A2(new_n669), .A3(new_n666), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT18), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n676), .A2(KEYINPUT18), .A3(new_n669), .A4(new_n666), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n668), .A2(KEYINPUT98), .A3(new_n671), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n674), .A2(new_n679), .A3(new_n680), .A4(new_n681), .ZN(new_n682));
  XOR2_X1   g481(.A(G113gat), .B(G141gat), .Z(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT96), .B(G197gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT11), .B(G169gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n687), .B(KEYINPUT12), .Z(new_n688));
  NAND2_X1  g487(.A1(new_n682), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT98), .B1(new_n668), .B2(new_n671), .ZN(new_n690));
  AOI211_X1 g489(.A(new_n673), .B(new_n670), .C1(new_n666), .C2(new_n667), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n688), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n692), .A2(new_n693), .A3(new_n680), .A4(new_n679), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n634), .A2(new_n665), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n202), .B1(new_n541), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n537), .A2(KEYINPUT94), .ZN(new_n698));
  INV_X1    g497(.A(new_n496), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n698), .A2(new_n540), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n479), .A2(new_n483), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n696), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n702), .A2(KEYINPUT107), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n697), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(new_n512), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(G1gat), .ZN(G1324gat));
  INV_X1    g506(.A(KEYINPUT42), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT16), .B(G8gat), .Z(new_n709));
  NAND4_X1  g508(.A1(new_n705), .A2(new_n708), .A3(new_n535), .A4(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT107), .B1(new_n702), .B2(new_n703), .ZN(new_n711));
  AOI211_X1 g510(.A(new_n202), .B(new_n696), .C1(new_n700), .C2(new_n701), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n535), .B(new_n709), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT42), .ZN(new_n714));
  INV_X1    g513(.A(G8gat), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n715), .B1(new_n705), .B2(new_n535), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n710), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(KEYINPUT108), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n719));
  OAI211_X1 g518(.A(new_n719), .B(new_n710), .C1(new_n714), .C2(new_n716), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(G1325gat));
  AOI21_X1  g520(.A(G15gat), .B1(new_n705), .B2(new_n480), .ZN(new_n722));
  INV_X1    g521(.A(new_n485), .ZN(new_n723));
  INV_X1    g522(.A(new_n487), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n726), .A2(G15gat), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n722), .B1(new_n705), .B2(new_n727), .ZN(G1326gat));
  AND2_X1   g527(.A1(new_n493), .A2(new_n494), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n465), .B1(new_n705), .B2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n705), .A2(new_n465), .A3(new_n729), .ZN(new_n732));
  XNOR2_X1  g531(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n733), .B1(new_n731), .B2(new_n732), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(G1327gat));
  NOR2_X1   g535(.A1(new_n664), .A2(new_n577), .ZN(new_n737));
  AND4_X1   g536(.A1(new_n702), .A2(new_n630), .A3(new_n695), .A4(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(G29gat), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n738), .A2(new_n739), .A3(new_n512), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT45), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT44), .B1(new_n541), .B2(new_n629), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n702), .A2(new_n743), .A3(new_n630), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT110), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n695), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n689), .A2(new_n694), .A3(KEYINPUT110), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n737), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n745), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n512), .ZN(new_n754));
  OAI21_X1  g553(.A(G29gat), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n741), .A2(new_n755), .ZN(G1328gat));
  INV_X1    g555(.A(new_n588), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n738), .A2(new_n535), .A3(new_n757), .ZN(new_n758));
  XOR2_X1   g557(.A(new_n758), .B(KEYINPUT46), .Z(new_n759));
  NAND2_X1  g558(.A1(new_n366), .A2(new_n367), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n588), .B1(new_n753), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(G1329gat));
  NAND3_X1  g561(.A1(new_n745), .A2(new_n726), .A3(new_n752), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G43gat), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT47), .ZN(new_n765));
  OR2_X1    g564(.A1(new_n765), .A2(KEYINPUT111), .ZN(new_n766));
  INV_X1    g565(.A(new_n480), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n767), .A2(G43gat), .ZN(new_n768));
  AOI22_X1  g567(.A1(new_n738), .A2(new_n768), .B1(KEYINPUT111), .B2(new_n765), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n764), .A2(new_n766), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n766), .B1(new_n764), .B2(new_n769), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n770), .A2(new_n771), .ZN(G1330gat));
  OAI21_X1  g571(.A(G50gat), .B1(new_n753), .B2(new_n477), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n495), .A2(G50gat), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n738), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n773), .A2(KEYINPUT48), .A3(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n745), .A2(new_n729), .A3(new_n752), .ZN(new_n777));
  AOI22_X1  g576(.A1(new_n777), .A2(G50gat), .B1(new_n738), .B2(new_n774), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n776), .B1(new_n778), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g578(.A1(new_n633), .A2(new_n750), .A3(new_n665), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n702), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(new_n754), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(new_n554), .ZN(G1332gat));
  NOR2_X1   g582(.A1(new_n781), .A2(new_n760), .ZN(new_n784));
  NOR2_X1   g583(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n785));
  AND2_X1   g584(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(new_n784), .B2(new_n785), .ZN(G1333gat));
  INV_X1    g587(.A(new_n781), .ZN(new_n789));
  AOI21_X1  g588(.A(G71gat), .B1(new_n789), .B2(new_n480), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n726), .A2(G71gat), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n790), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n792), .B(new_n793), .ZN(G1334gat));
  NAND2_X1  g593(.A1(new_n789), .A2(new_n729), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g595(.A1(new_n750), .A2(new_n577), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n664), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n798), .B1(new_n742), .B2(new_n744), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(G85gat), .B1(new_n800), .B2(new_n754), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n702), .A2(new_n630), .A3(new_n797), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n802), .B(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n512), .A2(new_n664), .A3(new_n435), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n801), .B1(new_n805), .B2(new_n806), .ZN(G1336gat));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n665), .A2(new_n760), .A3(G92gat), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n541), .A2(new_n629), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT51), .B1(new_n810), .B2(new_n797), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n802), .A2(new_n803), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n809), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n808), .B1(new_n813), .B2(KEYINPUT112), .ZN(new_n814));
  AOI211_X1 g613(.A(new_n760), .B(new_n798), .C1(new_n742), .C2(new_n744), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n813), .B1(new_n815), .B2(new_n598), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  OAI221_X1 g616(.A(new_n813), .B1(KEYINPUT112), .B2(new_n808), .C1(new_n815), .C2(new_n598), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(G1337gat));
  OAI21_X1  g618(.A(G99gat), .B1(new_n800), .B2(new_n725), .ZN(new_n820));
  OR3_X1    g619(.A1(new_n767), .A2(G99gat), .A3(new_n665), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n820), .B1(new_n805), .B2(new_n821), .ZN(G1338gat));
  INV_X1    g621(.A(G106gat), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(new_n799), .B2(new_n729), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n665), .A2(new_n477), .A3(G106gat), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n824), .B1(new_n804), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n804), .A2(new_n825), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n827), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n823), .B1(new_n799), .B2(new_n516), .ZN(new_n830));
  OAI22_X1  g629(.A1(new_n826), .A2(new_n827), .B1(new_n829), .B2(new_n830), .ZN(G1339gat));
  NOR3_X1   g630(.A1(new_n633), .A2(new_n750), .A3(new_n664), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n668), .A2(new_n671), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n669), .B1(new_n676), .B2(new_n666), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n687), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n694), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n664), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n645), .A2(new_n646), .ZN(new_n840));
  OAI21_X1  g639(.A(KEYINPUT54), .B1(new_n840), .B2(new_n635), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n635), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT105), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n647), .A2(new_n648), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n841), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n658), .B1(new_n647), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n839), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  OAI211_X1 g648(.A(KEYINPUT55), .B(new_n847), .C1(new_n651), .C2(new_n841), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n849), .A2(new_n661), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n838), .B1(new_n749), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n629), .ZN(new_n853));
  OR3_X1    g652(.A1(new_n851), .A2(new_n629), .A3(new_n836), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n832), .B1(new_n855), .B2(new_n578), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n729), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n754), .A2(new_n535), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(new_n480), .A3(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n860), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n695), .ZN(new_n864));
  OAI21_X1  g663(.A(G113gat), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n634), .A2(new_n665), .A3(new_n749), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n851), .A2(new_n629), .A3(new_n836), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n867), .B1(new_n852), .B2(new_n629), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n866), .B1(new_n868), .B2(new_n577), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n315), .A2(new_n477), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n870), .A2(new_n754), .A3(new_n535), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n267), .A3(new_n750), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n865), .A2(new_n873), .ZN(G1340gat));
  OAI21_X1  g673(.A(G120gat), .B1(new_n863), .B2(new_n665), .ZN(new_n875));
  INV_X1    g674(.A(new_n872), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n665), .A2(new_n276), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(G1341gat));
  INV_X1    g677(.A(new_n265), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n578), .A2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(KEYINPUT114), .B1(new_n863), .B2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT114), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n861), .A2(new_n883), .A3(new_n862), .A4(new_n880), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n879), .B1(new_n876), .B2(new_n578), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n882), .A2(new_n884), .A3(new_n885), .ZN(G1342gat));
  OAI21_X1  g685(.A(G134gat), .B1(new_n863), .B2(new_n629), .ZN(new_n887));
  INV_X1    g686(.A(G134gat), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n872), .A2(new_n888), .A3(new_n630), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT56), .ZN(new_n890));
  XOR2_X1   g689(.A(new_n890), .B(KEYINPUT115), .Z(new_n891));
  OAI211_X1 g690(.A(new_n887), .B(new_n891), .C1(KEYINPUT56), .C2(new_n889), .ZN(G1343gat));
  NOR2_X1   g691(.A1(new_n856), .A2(new_n477), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n725), .A2(new_n858), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n895), .A2(G141gat), .A3(new_n864), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n849), .A2(new_n850), .A3(new_n661), .A4(new_n695), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n630), .B1(new_n838), .B2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT116), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n854), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n898), .A2(new_n899), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n578), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n866), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(KEYINPUT57), .A3(new_n729), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT57), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n905), .B1(new_n856), .B2(new_n477), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n907), .A2(new_n894), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n750), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n896), .B1(new_n909), .B2(G141gat), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT58), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n370), .B1(new_n908), .B2(new_n695), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n896), .A2(KEYINPUT58), .ZN(new_n913));
  OAI22_X1  g712(.A1(new_n910), .A2(new_n911), .B1(new_n912), .B2(new_n913), .ZN(G1344gat));
  NAND4_X1  g713(.A1(new_n893), .A2(new_n373), .A3(new_n664), .A4(new_n894), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT59), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n869), .A2(KEYINPUT57), .A3(new_n516), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT117), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n869), .A2(KEYINPUT117), .A3(KEYINPUT57), .A4(new_n516), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n634), .A2(new_n665), .A3(new_n864), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n578), .B1(new_n898), .B2(new_n867), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n905), .B1(new_n923), .B2(new_n495), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n919), .A2(new_n920), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(new_n664), .A3(new_n894), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n373), .B1(new_n926), .B2(KEYINPUT118), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT118), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n925), .A2(new_n928), .A3(new_n664), .A4(new_n894), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n916), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  AOI211_X1 g729(.A(KEYINPUT59), .B(new_n373), .C1(new_n908), .C2(new_n664), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n915), .B1(new_n930), .B2(new_n931), .ZN(G1345gat));
  OAI21_X1  g731(.A(new_n391), .B1(new_n895), .B2(new_n578), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n907), .A2(new_n894), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n577), .A2(G155gat), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  XOR2_X1   g735(.A(new_n936), .B(KEYINPUT119), .Z(G1346gat));
  OAI21_X1  g736(.A(G162gat), .B1(new_n934), .B2(new_n629), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n893), .A2(new_n392), .A3(new_n630), .A4(new_n894), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT120), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(KEYINPUT121), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT121), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n938), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n945), .ZN(G1347gat));
  NAND2_X1  g745(.A1(new_n754), .A2(new_n535), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n947), .A2(new_n767), .ZN(new_n948));
  XOR2_X1   g747(.A(new_n948), .B(KEYINPUT122), .Z(new_n949));
  NAND2_X1  g748(.A1(new_n857), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(G169gat), .B1(new_n950), .B2(new_n864), .ZN(new_n951));
  XOR2_X1   g750(.A(new_n951), .B(KEYINPUT123), .Z(new_n952));
  NOR2_X1   g751(.A1(new_n870), .A2(new_n947), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n869), .A2(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(G169gat), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n954), .A2(new_n955), .A3(new_n750), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n952), .A2(new_n956), .ZN(G1348gat));
  OR3_X1    g756(.A1(new_n950), .A2(new_n233), .A3(new_n665), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT124), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n958), .A2(new_n959), .ZN(new_n961));
  AOI21_X1  g760(.A(G176gat), .B1(new_n954), .B2(new_n664), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(G1349gat));
  NAND3_X1  g762(.A1(new_n954), .A2(new_n252), .A3(new_n577), .ZN(new_n964));
  XOR2_X1   g763(.A(new_n964), .B(KEYINPUT125), .Z(new_n965));
  OAI21_X1  g764(.A(G183gat), .B1(new_n950), .B2(new_n578), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(KEYINPUT60), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT60), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n965), .A2(new_n969), .A3(new_n966), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n968), .A2(new_n970), .ZN(G1350gat));
  OAI21_X1  g770(.A(G190gat), .B1(new_n950), .B2(new_n629), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT61), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n954), .A2(new_n251), .A3(new_n630), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(G1351gat));
  NAND3_X1  g774(.A1(new_n725), .A2(new_n535), .A3(new_n516), .ZN(new_n976));
  OR2_X1    g775(.A1(new_n976), .A2(KEYINPUT126), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n512), .B1(new_n976), .B2(KEYINPUT126), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n977), .A2(new_n869), .A3(new_n978), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n980), .A2(new_n329), .A3(new_n750), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n726), .A2(new_n947), .ZN(new_n982));
  AND2_X1   g781(.A1(new_n925), .A2(new_n982), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n983), .A2(new_n695), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n981), .B1(new_n984), .B2(new_n329), .ZN(G1352gat));
  NOR3_X1   g784(.A1(new_n979), .A2(G204gat), .A3(new_n665), .ZN(new_n986));
  XNOR2_X1  g785(.A(new_n986), .B(KEYINPUT62), .ZN(new_n987));
  AND3_X1   g786(.A1(new_n925), .A2(new_n664), .A3(new_n982), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n987), .B1(new_n330), .B2(new_n988), .ZN(G1353gat));
  NOR3_X1   g788(.A1(new_n979), .A2(G211gat), .A3(new_n578), .ZN(new_n990));
  XNOR2_X1  g789(.A(new_n990), .B(KEYINPUT127), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n983), .A2(new_n577), .ZN(new_n992));
  AOI21_X1  g791(.A(KEYINPUT63), .B1(new_n992), .B2(G211gat), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT63), .ZN(new_n994));
  AOI211_X1 g793(.A(new_n994), .B(new_n323), .C1(new_n983), .C2(new_n577), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n991), .B1(new_n993), .B2(new_n995), .ZN(G1354gat));
  AOI21_X1  g795(.A(G218gat), .B1(new_n980), .B2(new_n630), .ZN(new_n997));
  NOR2_X1   g796(.A1(new_n629), .A2(new_n324), .ZN(new_n998));
  AOI21_X1  g797(.A(new_n997), .B1(new_n983), .B2(new_n998), .ZN(G1355gat));
endmodule


