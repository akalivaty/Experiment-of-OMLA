

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763;

  BUF_X1 U375 ( .A(G953), .Z(n403) );
  NOR2_X1 U376 ( .A1(n403), .A2(G237), .ZN(n514) );
  XNOR2_X1 U377 ( .A(n379), .B(n382), .ZN(n743) );
  OR2_X1 U378 ( .A1(n593), .A2(n361), .ZN(n353) );
  NAND2_X2 U379 ( .A1(n417), .A2(n423), .ZN(n540) );
  XNOR2_X1 U380 ( .A(n372), .B(KEYINPUT40), .ZN(n646) );
  NOR2_X2 U381 ( .A1(n638), .A2(n736), .ZN(n639) );
  NOR2_X2 U382 ( .A1(n626), .A2(n736), .ZN(n627) );
  XNOR2_X1 U383 ( .A(n535), .B(n534), .ZN(n557) );
  XNOR2_X2 U384 ( .A(n467), .B(G134), .ZN(n504) );
  NOR2_X1 U385 ( .A1(n636), .A2(G902), .ZN(n535) );
  XNOR2_X2 U386 ( .A(n598), .B(KEYINPUT102), .ZN(n563) );
  XNOR2_X2 U387 ( .A(n540), .B(KEYINPUT38), .ZN(n705) );
  XNOR2_X1 U388 ( .A(n588), .B(n587), .ZN(n398) );
  AND2_X1 U389 ( .A1(n370), .A2(n368), .ZN(n367) );
  XNOR2_X1 U390 ( .A(n499), .B(n498), .ZN(n559) );
  XNOR2_X1 U391 ( .A(n411), .B(KEYINPUT100), .ZN(n673) );
  NAND2_X1 U392 ( .A1(n418), .A2(n423), .ZN(n572) );
  XNOR2_X1 U393 ( .A(KEYINPUT66), .B(G101), .ZN(n505) );
  INV_X1 U394 ( .A(KEYINPUT80), .ZN(n376) );
  INV_X1 U395 ( .A(G128), .ZN(n440) );
  BUF_X1 U396 ( .A(KEYINPUT44), .Z(n361) );
  INV_X1 U397 ( .A(KEYINPUT86), .ZN(n373) );
  INV_X1 U398 ( .A(KEYINPUT39), .ZN(n366) );
  INV_X1 U399 ( .A(G146), .ZN(n485) );
  XNOR2_X1 U400 ( .A(n377), .B(n376), .ZN(n409) );
  NAND2_X1 U401 ( .A1(n398), .A2(n437), .ZN(n753) );
  NAND2_X1 U402 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U403 ( .A1(n362), .A2(n356), .ZN(n359) );
  NOR2_X1 U404 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U405 ( .A1(n399), .A2(n670), .ZN(n372) );
  NAND2_X1 U406 ( .A1(n367), .A2(n363), .ZN(n399) );
  XNOR2_X1 U407 ( .A(n402), .B(n569), .ZN(n762) );
  NAND2_X1 U408 ( .A1(n559), .A2(n374), .ZN(n416) );
  NOR2_X1 U409 ( .A1(n412), .A2(n673), .ZN(n574) );
  NOR2_X1 U410 ( .A1(n410), .A2(n689), .ZN(n553) );
  AND2_X1 U411 ( .A1(n433), .A2(n366), .ZN(n365) );
  NOR2_X1 U412 ( .A1(n707), .A2(n709), .ZN(n561) );
  OR2_X1 U413 ( .A1(n609), .A2(n690), .ZN(n410) );
  AND2_X1 U414 ( .A1(n705), .A2(n434), .ZN(n433) );
  XNOR2_X1 U415 ( .A(n400), .B(n435), .ZN(n432) );
  BUF_X1 U416 ( .A(n689), .Z(n374) );
  XNOR2_X1 U417 ( .A(n566), .B(n513), .ZN(n689) );
  XNOR2_X1 U418 ( .A(n598), .B(KEYINPUT6), .ZN(n609) );
  XOR2_X1 U419 ( .A(n641), .B(n640), .Z(n394) );
  OR2_X1 U420 ( .A1(n649), .A2(G902), .ZN(n427) );
  OR2_X2 U421 ( .A1(n641), .A2(G902), .ZN(n385) );
  XNOR2_X1 U422 ( .A(n622), .B(KEYINPUT59), .ZN(n623) );
  XNOR2_X1 U423 ( .A(n386), .B(n752), .ZN(n641) );
  XNOR2_X1 U424 ( .A(n743), .B(n448), .ZN(n630) );
  XNOR2_X1 U425 ( .A(n388), .B(n375), .ZN(n649) );
  XNOR2_X1 U426 ( .A(n517), .B(n378), .ZN(n386) );
  XNOR2_X1 U427 ( .A(n510), .B(n505), .ZN(n375) );
  XNOR2_X1 U428 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U429 ( .A(n504), .B(n503), .ZN(n752) );
  XNOR2_X1 U430 ( .A(n518), .B(KEYINPUT16), .ZN(n379) );
  XNOR2_X1 U431 ( .A(n518), .B(n505), .ZN(n378) );
  NOR2_X1 U432 ( .A1(n492), .A2(n620), .ZN(n621) );
  XNOR2_X1 U433 ( .A(KEYINPUT18), .B(G125), .ZN(n442) );
  XOR2_X1 U434 ( .A(G122), .B(G113), .Z(n476) );
  XOR2_X1 U435 ( .A(G125), .B(KEYINPUT10), .Z(n484) );
  XNOR2_X1 U436 ( .A(G137), .B(G128), .ZN(n520) );
  NAND2_X1 U437 ( .A1(n497), .A2(n601), .ZN(n499) );
  XNOR2_X2 U438 ( .A(n459), .B(n458), .ZN(n601) );
  NAND2_X1 U439 ( .A1(n371), .A2(KEYINPUT39), .ZN(n370) );
  BUF_X1 U440 ( .A(n636), .Z(n354) );
  AND2_X2 U441 ( .A1(n438), .A2(n355), .ZN(n389) );
  XNOR2_X2 U442 ( .A(n616), .B(n395), .ZN(n355) );
  INV_X1 U443 ( .A(n355), .ZN(n737) );
  NAND2_X1 U444 ( .A1(n355), .A2(n409), .ZN(n408) );
  XNOR2_X2 U445 ( .A(n594), .B(KEYINPUT81), .ZN(n362) );
  NOR2_X1 U446 ( .A1(n595), .A2(n353), .ZN(n356) );
  NOR2_X1 U447 ( .A1(n595), .A2(n361), .ZN(n357) );
  NAND2_X1 U448 ( .A1(n357), .A2(n362), .ZN(n358) );
  NAND2_X1 U449 ( .A1(n358), .A2(n593), .ZN(n360) );
  NAND2_X1 U450 ( .A1(n360), .A2(n359), .ZN(n615) );
  NAND2_X2 U451 ( .A1(n591), .A2(n592), .ZN(n594) );
  XNOR2_X2 U452 ( .A(n424), .B(KEYINPUT35), .ZN(n595) );
  NAND2_X1 U453 ( .A1(n432), .A2(n364), .ZN(n363) );
  AND2_X1 U454 ( .A1(n578), .A2(n365), .ZN(n364) );
  NAND2_X1 U455 ( .A1(n369), .A2(KEYINPUT39), .ZN(n368) );
  NAND2_X1 U456 ( .A1(n578), .A2(n433), .ZN(n369) );
  INV_X1 U457 ( .A(n432), .ZN(n371) );
  XNOR2_X1 U458 ( .A(n601), .B(n373), .ZN(n604) );
  AND2_X2 U459 ( .A1(n419), .A2(n391), .ZN(n418) );
  NAND2_X1 U460 ( .A1(n398), .A2(n429), .ZN(n377) );
  XNOR2_X2 U461 ( .A(n381), .B(n380), .ZN(n518) );
  XNOR2_X2 U462 ( .A(KEYINPUT72), .B(KEYINPUT3), .ZN(n380) );
  XNOR2_X2 U463 ( .A(G119), .B(G113), .ZN(n381) );
  XNOR2_X2 U464 ( .A(n465), .B(n509), .ZN(n382) );
  XNOR2_X2 U465 ( .A(n383), .B(G104), .ZN(n509) );
  XNOR2_X2 U466 ( .A(KEYINPUT85), .B(G110), .ZN(n383) );
  XNOR2_X2 U467 ( .A(n384), .B(n439), .ZN(n465) );
  XNOR2_X2 U468 ( .A(G116), .B(G122), .ZN(n384) );
  XNOR2_X2 U469 ( .A(n385), .B(G472), .ZN(n598) );
  XNOR2_X1 U470 ( .A(n406), .B(KEYINPUT64), .ZN(n387) );
  XNOR2_X1 U471 ( .A(n406), .B(KEYINPUT64), .ZN(n731) );
  BUF_X1 U472 ( .A(n752), .Z(n388) );
  NOR2_X2 U473 ( .A1(n389), .A2(n621), .ZN(n407) );
  INV_X1 U474 ( .A(G237), .ZN(n449) );
  XNOR2_X1 U475 ( .A(G140), .B(KEYINPUT68), .ZN(n483) );
  NAND2_X1 U476 ( .A1(n492), .A2(n421), .ZN(n420) );
  INV_X1 U477 ( .A(n450), .ZN(n421) );
  INV_X1 U478 ( .A(KEYINPUT73), .ZN(n593) );
  XNOR2_X1 U479 ( .A(G119), .B(G110), .ZN(n519) );
  XOR2_X1 U480 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n522) );
  INV_X1 U481 ( .A(KEYINPUT48), .ZN(n587) );
  NOR2_X1 U482 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U483 ( .A1(n430), .A2(n620), .ZN(n429) );
  INV_X1 U484 ( .A(n437), .ZN(n430) );
  XNOR2_X1 U485 ( .A(n414), .B(n413), .ZN(n412) );
  INV_X1 U486 ( .A(KEYINPUT104), .ZN(n413) );
  NOR2_X1 U487 ( .A1(n707), .A2(n545), .ZN(n497) );
  XNOR2_X1 U488 ( .A(n539), .B(KEYINPUT67), .ZN(n552) );
  INV_X1 U489 ( .A(KEYINPUT69), .ZN(n472) );
  NAND2_X1 U490 ( .A1(n619), .A2(n450), .ZN(n422) );
  INV_X1 U491 ( .A(G107), .ZN(n439) );
  XOR2_X1 U492 ( .A(KEYINPUT96), .B(KEYINPUT9), .Z(n461) );
  XNOR2_X1 U493 ( .A(KEYINPUT7), .B(KEYINPUT97), .ZN(n460) );
  XNOR2_X1 U494 ( .A(G143), .B(G104), .ZN(n475) );
  XOR2_X1 U495 ( .A(KEYINPUT12), .B(KEYINPUT90), .Z(n478) );
  BUF_X1 U496 ( .A(n703), .Z(n722) );
  INV_X1 U497 ( .A(KEYINPUT30), .ZN(n435) );
  INV_X1 U498 ( .A(n544), .ZN(n434) );
  XNOR2_X1 U499 ( .A(n469), .B(n405), .ZN(n555) );
  XNOR2_X1 U500 ( .A(n470), .B(n471), .ZN(n405) );
  XNOR2_X1 U501 ( .A(n528), .B(n527), .ZN(n636) );
  XNOR2_X1 U502 ( .A(G107), .B(G140), .ZN(n507) );
  XNOR2_X1 U503 ( .A(n408), .B(KEYINPUT75), .ZN(n684) );
  NAND2_X1 U504 ( .A1(n577), .A2(n576), .ZN(n679) );
  XNOR2_X1 U505 ( .A(n404), .B(KEYINPUT32), .ZN(n592) );
  XNOR2_X1 U506 ( .A(n416), .B(KEYINPUT103), .ZN(n537) );
  NAND2_X1 U507 ( .A1(n415), .A2(n610), .ZN(n653) );
  XOR2_X1 U508 ( .A(n482), .B(n481), .Z(n390) );
  INV_X1 U509 ( .A(n396), .ZN(n397) );
  BUF_X1 U510 ( .A(n552), .Z(n690) );
  INV_X1 U511 ( .A(n552), .ZN(n431) );
  AND2_X1 U512 ( .A1(n422), .A2(n704), .ZN(n391) );
  AND2_X1 U513 ( .A1(n432), .A2(n434), .ZN(n392) );
  XOR2_X1 U514 ( .A(n630), .B(n629), .Z(n393) );
  XOR2_X1 U515 ( .A(KEYINPUT79), .B(KEYINPUT45), .Z(n395) );
  AND2_X1 U516 ( .A1(n625), .A2(n403), .ZN(n736) );
  INV_X1 U517 ( .A(n557), .ZN(n396) );
  NOR2_X1 U518 ( .A1(n609), .A2(n548), .ZN(n414) );
  BUF_X1 U519 ( .A(n753), .Z(n428) );
  NAND2_X1 U520 ( .A1(n563), .A2(n704), .ZN(n400) );
  NAND2_X1 U521 ( .A1(n399), .A2(n662), .ZN(n589) );
  XNOR2_X2 U522 ( .A(n605), .B(KEYINPUT105), .ZN(n578) );
  NAND2_X1 U523 ( .A1(n646), .A2(n401), .ZN(n571) );
  INV_X1 U524 ( .A(n762), .ZN(n401) );
  NAND2_X1 U525 ( .A1(n660), .A2(n721), .ZN(n402) );
  NAND2_X1 U526 ( .A1(n559), .A2(n436), .ZN(n404) );
  NOR2_X2 U527 ( .A1(n684), .A2(n407), .ZN(n406) );
  NOR2_X2 U528 ( .A1(n557), .A2(n545), .ZN(n539) );
  NAND2_X1 U529 ( .A1(n555), .A2(n543), .ZN(n411) );
  INV_X1 U530 ( .A(n416), .ZN(n415) );
  OR2_X2 U531 ( .A1(n630), .A2(n420), .ZN(n419) );
  AND2_X1 U532 ( .A1(n419), .A2(n422), .ZN(n417) );
  NAND2_X1 U533 ( .A1(n630), .A2(n450), .ZN(n423) );
  NOR2_X1 U534 ( .A1(n703), .A2(n604), .ZN(n426) );
  OR2_X1 U535 ( .A1(n428), .A2(n737), .ZN(n682) );
  NAND2_X1 U536 ( .A1(n425), .A2(n556), .ZN(n424) );
  XNOR2_X1 U537 ( .A(n426), .B(KEYINPUT34), .ZN(n425) );
  XNOR2_X2 U538 ( .A(n427), .B(n512), .ZN(n566) );
  XNOR2_X1 U539 ( .A(n753), .B(n617), .ZN(n618) );
  NAND2_X2 U540 ( .A1(n431), .A2(n566), .ZN(n605) );
  AND2_X1 U541 ( .A1(n558), .A2(n609), .ZN(n436) );
  AND2_X1 U542 ( .A1(n590), .A2(n589), .ZN(n437) );
  AND2_X1 U543 ( .A1(n618), .A2(n619), .ZN(n438) );
  INV_X1 U544 ( .A(KEYINPUT74), .ZN(n617) );
  XNOR2_X1 U545 ( .A(n531), .B(n530), .ZN(n532) );
  INV_X1 U546 ( .A(n736), .ZN(n632) );
  BUF_X1 U547 ( .A(n646), .Z(n647) );
  XNOR2_X2 U548 ( .A(G143), .B(KEYINPUT77), .ZN(n441) );
  XNOR2_X2 U549 ( .A(n441), .B(n440), .ZN(n467) );
  XNOR2_X2 U550 ( .A(G146), .B(KEYINPUT4), .ZN(n500) );
  XNOR2_X1 U551 ( .A(n500), .B(n442), .ZN(n443) );
  XNOR2_X1 U552 ( .A(n467), .B(n443), .ZN(n447) );
  INV_X2 U553 ( .A(G953), .ZN(n745) );
  NAND2_X1 U554 ( .A1(n745), .A2(G224), .ZN(n444) );
  XNOR2_X1 U555 ( .A(n444), .B(KEYINPUT17), .ZN(n445) );
  XNOR2_X1 U556 ( .A(n445), .B(n505), .ZN(n446) );
  XNOR2_X1 U557 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U558 ( .A(G902), .B(KEYINPUT15), .ZN(n492) );
  INV_X1 U559 ( .A(n492), .ZN(n619) );
  INV_X1 U560 ( .A(G902), .ZN(n486) );
  NAND2_X1 U561 ( .A1(n486), .A2(n449), .ZN(n451) );
  NAND2_X1 U562 ( .A1(n451), .A2(G210), .ZN(n450) );
  NAND2_X1 U563 ( .A1(n451), .A2(G214), .ZN(n704) );
  XNOR2_X2 U564 ( .A(n572), .B(KEYINPUT19), .ZN(n661) );
  NAND2_X1 U565 ( .A1(G237), .A2(G234), .ZN(n452) );
  XNOR2_X1 U566 ( .A(n452), .B(KEYINPUT14), .ZN(n685) );
  NOR2_X1 U567 ( .A1(G902), .A2(n745), .ZN(n454) );
  NOR2_X1 U568 ( .A1(n403), .A2(G952), .ZN(n453) );
  NOR2_X1 U569 ( .A1(n454), .A2(n453), .ZN(n455) );
  AND2_X1 U570 ( .A1(n685), .A2(n455), .ZN(n542) );
  NAND2_X1 U571 ( .A1(n403), .A2(G898), .ZN(n456) );
  AND2_X1 U572 ( .A1(n542), .A2(n456), .ZN(n457) );
  NAND2_X1 U573 ( .A1(n661), .A2(n457), .ZN(n459) );
  XNOR2_X1 U574 ( .A(KEYINPUT83), .B(KEYINPUT0), .ZN(n458) );
  XNOR2_X1 U575 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n470) );
  XNOR2_X1 U576 ( .A(n461), .B(n460), .ZN(n464) );
  NAND2_X1 U577 ( .A1(G234), .A2(n745), .ZN(n462) );
  XOR2_X1 U578 ( .A(KEYINPUT8), .B(n462), .Z(n524) );
  NAND2_X1 U579 ( .A1(G217), .A2(n524), .ZN(n463) );
  XOR2_X1 U580 ( .A(n464), .B(n463), .Z(n466) );
  XNOR2_X1 U581 ( .A(n466), .B(n465), .ZN(n468) );
  XNOR2_X1 U582 ( .A(n504), .B(n468), .ZN(n733) );
  NOR2_X1 U583 ( .A1(G902), .A2(n733), .ZN(n469) );
  INV_X1 U584 ( .A(G478), .ZN(n471) );
  XNOR2_X1 U585 ( .A(n472), .B(G131), .ZN(n501) );
  XOR2_X1 U586 ( .A(n501), .B(KEYINPUT91), .Z(n474) );
  NAND2_X1 U587 ( .A1(n514), .A2(G214), .ZN(n473) );
  XNOR2_X1 U588 ( .A(n474), .B(n473), .ZN(n482) );
  XNOR2_X1 U589 ( .A(n476), .B(n475), .ZN(n480) );
  XNOR2_X1 U590 ( .A(KEYINPUT11), .B(KEYINPUT92), .ZN(n477) );
  XNOR2_X1 U591 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U592 ( .A(n480), .B(n479), .Z(n481) );
  XNOR2_X1 U593 ( .A(n484), .B(n483), .ZN(n751) );
  XNOR2_X1 U594 ( .A(n751), .B(n485), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n390), .B(n527), .ZN(n622) );
  NAND2_X1 U596 ( .A1(n622), .A2(n486), .ZN(n491) );
  XOR2_X1 U597 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n488) );
  XNOR2_X1 U598 ( .A(KEYINPUT95), .B(KEYINPUT13), .ZN(n487) );
  XNOR2_X1 U599 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U600 ( .A(G475), .B(n489), .ZN(n490) );
  XNOR2_X1 U601 ( .A(n491), .B(n490), .ZN(n543) );
  INV_X1 U602 ( .A(n543), .ZN(n554) );
  NAND2_X1 U603 ( .A1(n555), .A2(n554), .ZN(n707) );
  NAND2_X1 U604 ( .A1(n492), .A2(G234), .ZN(n494) );
  XNOR2_X1 U605 ( .A(KEYINPUT88), .B(KEYINPUT20), .ZN(n493) );
  XNOR2_X1 U606 ( .A(n494), .B(n493), .ZN(n529) );
  NAND2_X1 U607 ( .A1(n529), .A2(G221), .ZN(n496) );
  INV_X1 U608 ( .A(KEYINPUT21), .ZN(n495) );
  XNOR2_X1 U609 ( .A(n496), .B(n495), .ZN(n686) );
  INV_X1 U610 ( .A(n686), .ZN(n545) );
  INV_X1 U611 ( .A(KEYINPUT22), .ZN(n498) );
  XNOR2_X1 U612 ( .A(n500), .B(G137), .ZN(n502) );
  XNOR2_X1 U613 ( .A(n502), .B(n501), .ZN(n503) );
  NAND2_X1 U614 ( .A1(n745), .A2(G227), .ZN(n506) );
  XNOR2_X1 U615 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U616 ( .A(n509), .B(n508), .ZN(n510) );
  INV_X1 U617 ( .A(KEYINPUT71), .ZN(n511) );
  XNOR2_X1 U618 ( .A(n511), .B(G469), .ZN(n512) );
  XNOR2_X1 U619 ( .A(KEYINPUT65), .B(KEYINPUT1), .ZN(n513) );
  XNOR2_X1 U620 ( .A(G116), .B(KEYINPUT5), .ZN(n516) );
  NAND2_X1 U621 ( .A1(G210), .A2(n514), .ZN(n515) );
  XNOR2_X1 U622 ( .A(n516), .B(n515), .ZN(n517) );
  INV_X1 U623 ( .A(n519), .ZN(n521) );
  XNOR2_X1 U624 ( .A(n521), .B(n520), .ZN(n523) );
  XNOR2_X1 U625 ( .A(n523), .B(n522), .ZN(n526) );
  NAND2_X1 U626 ( .A1(G221), .A2(n524), .ZN(n525) );
  XNOR2_X1 U627 ( .A(n526), .B(n525), .ZN(n528) );
  AND2_X1 U628 ( .A1(G217), .A2(n529), .ZN(n533) );
  XNOR2_X1 U629 ( .A(KEYINPUT25), .B(KEYINPUT87), .ZN(n531) );
  INV_X1 U630 ( .A(KEYINPUT76), .ZN(n530) );
  NOR2_X1 U631 ( .A1(n563), .A2(n396), .ZN(n536) );
  NAND2_X1 U632 ( .A1(n537), .A2(n536), .ZN(n591) );
  XOR2_X1 U633 ( .A(G110), .B(KEYINPUT109), .Z(n538) );
  XNOR2_X1 U634 ( .A(n591), .B(n538), .ZN(G12) );
  NAND2_X1 U635 ( .A1(n403), .A2(G900), .ZN(n541) );
  NAND2_X1 U636 ( .A1(n542), .A2(n541), .ZN(n544) );
  OR2_X1 U637 ( .A1(n555), .A2(n543), .ZN(n677) );
  INV_X1 U638 ( .A(n677), .ZN(n662) );
  XNOR2_X1 U639 ( .A(n589), .B(G134), .ZN(G36) );
  NOR2_X1 U640 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U641 ( .A(n546), .B(KEYINPUT70), .ZN(n547) );
  AND2_X1 U642 ( .A1(n397), .A2(n547), .ZN(n562) );
  INV_X1 U643 ( .A(n562), .ZN(n548) );
  NAND2_X1 U644 ( .A1(n574), .A2(n704), .ZN(n549) );
  INV_X1 U645 ( .A(n374), .ZN(n576) );
  NOR2_X1 U646 ( .A1(n549), .A2(n576), .ZN(n550) );
  XOR2_X1 U647 ( .A(KEYINPUT43), .B(n550), .Z(n551) );
  NAND2_X1 U648 ( .A1(n551), .A2(n540), .ZN(n590) );
  XNOR2_X1 U649 ( .A(n590), .B(G140), .ZN(G42) );
  XNOR2_X1 U650 ( .A(n553), .B(KEYINPUT33), .ZN(n703) );
  OR2_X1 U651 ( .A1(n555), .A2(n554), .ZN(n579) );
  INV_X1 U652 ( .A(n579), .ZN(n556) );
  XOR2_X1 U653 ( .A(n595), .B(G122), .Z(G24) );
  XNOR2_X1 U654 ( .A(n397), .B(KEYINPUT101), .ZN(n687) );
  NOR2_X1 U655 ( .A1(n687), .A2(n689), .ZN(n558) );
  XNOR2_X1 U656 ( .A(n592), .B(G119), .ZN(G21) );
  INV_X1 U657 ( .A(n673), .ZN(n670) );
  NAND2_X1 U658 ( .A1(n705), .A2(n704), .ZN(n709) );
  XNOR2_X1 U659 ( .A(KEYINPUT41), .B(KEYINPUT107), .ZN(n560) );
  XNOR2_X1 U660 ( .A(n561), .B(n560), .ZN(n721) );
  NAND2_X1 U661 ( .A1(n563), .A2(n562), .ZN(n565) );
  INV_X1 U662 ( .A(KEYINPUT28), .ZN(n564) );
  XNOR2_X1 U663 ( .A(n565), .B(n564), .ZN(n568) );
  XNOR2_X1 U664 ( .A(n566), .B(KEYINPUT106), .ZN(n567) );
  AND2_X1 U665 ( .A1(n568), .A2(n567), .ZN(n660) );
  INV_X1 U666 ( .A(KEYINPUT42), .ZN(n569) );
  INV_X1 U667 ( .A(KEYINPUT46), .ZN(n570) );
  XNOR2_X1 U668 ( .A(n571), .B(n570), .ZN(n586) );
  INV_X1 U669 ( .A(n572), .ZN(n573) );
  NAND2_X1 U670 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U671 ( .A(KEYINPUT36), .B(n575), .Z(n577) );
  AND2_X1 U672 ( .A1(n578), .A2(n392), .ZN(n581) );
  NOR2_X1 U673 ( .A1(n579), .A2(n540), .ZN(n580) );
  NAND2_X1 U674 ( .A1(n581), .A2(n580), .ZN(n669) );
  NAND2_X1 U675 ( .A1(n679), .A2(n669), .ZN(n584) );
  AND2_X1 U676 ( .A1(n661), .A2(n660), .ZN(n671) );
  NAND2_X1 U677 ( .A1(n673), .A2(n677), .ZN(n708) );
  NAND2_X1 U678 ( .A1(n671), .A2(n708), .ZN(n582) );
  XNOR2_X1 U679 ( .A(n582), .B(KEYINPUT47), .ZN(n583) );
  NAND2_X1 U680 ( .A1(n586), .A2(n585), .ZN(n588) );
  INV_X1 U681 ( .A(KEYINPUT2), .ZN(n620) );
  INV_X1 U682 ( .A(KEYINPUT44), .ZN(n596) );
  NOR2_X1 U683 ( .A1(n597), .A2(n596), .ZN(n613) );
  BUF_X1 U684 ( .A(n598), .Z(n599) );
  NAND2_X1 U685 ( .A1(n431), .A2(n599), .ZN(n600) );
  NOR2_X1 U686 ( .A1(n600), .A2(n374), .ZN(n696) );
  NAND2_X1 U687 ( .A1(n696), .A2(n601), .ZN(n603) );
  XNOR2_X1 U688 ( .A(KEYINPUT89), .B(KEYINPUT31), .ZN(n602) );
  XNOR2_X1 U689 ( .A(n603), .B(n602), .ZN(n676) );
  INV_X1 U690 ( .A(n604), .ZN(n607) );
  NOR2_X1 U691 ( .A1(n605), .A2(n599), .ZN(n606) );
  NAND2_X1 U692 ( .A1(n607), .A2(n606), .ZN(n657) );
  NAND2_X1 U693 ( .A1(n676), .A2(n657), .ZN(n608) );
  NAND2_X1 U694 ( .A1(n608), .A2(n708), .ZN(n611) );
  AND2_X1 U695 ( .A1(n609), .A2(n687), .ZN(n610) );
  NAND2_X1 U696 ( .A1(n611), .A2(n653), .ZN(n612) );
  NOR2_X1 U697 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U698 ( .A1(n731), .A2(G475), .ZN(n624) );
  XNOR2_X1 U699 ( .A(n624), .B(n623), .ZN(n626) );
  INV_X1 U700 ( .A(G952), .ZN(n625) );
  XNOR2_X1 U701 ( .A(n627), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U702 ( .A1(n387), .A2(G210), .ZN(n631) );
  XOR2_X1 U703 ( .A(KEYINPUT78), .B(KEYINPUT54), .Z(n628) );
  XNOR2_X1 U704 ( .A(n628), .B(KEYINPUT55), .ZN(n629) );
  XNOR2_X1 U705 ( .A(n631), .B(n393), .ZN(n633) );
  AND2_X2 U706 ( .A1(n633), .A2(n632), .ZN(n635) );
  XOR2_X1 U707 ( .A(KEYINPUT121), .B(KEYINPUT56), .Z(n634) );
  XNOR2_X1 U708 ( .A(n635), .B(n634), .ZN(G51) );
  NAND2_X1 U709 ( .A1(n731), .A2(G217), .ZN(n637) );
  XNOR2_X1 U710 ( .A(n637), .B(n354), .ZN(n638) );
  XNOR2_X1 U711 ( .A(n639), .B(KEYINPUT122), .ZN(G66) );
  NAND2_X1 U712 ( .A1(n387), .A2(G472), .ZN(n642) );
  XNOR2_X1 U713 ( .A(KEYINPUT84), .B(KEYINPUT62), .ZN(n640) );
  XNOR2_X1 U714 ( .A(n642), .B(n394), .ZN(n643) );
  AND2_X2 U715 ( .A1(n643), .A2(n632), .ZN(n645) );
  XOR2_X1 U716 ( .A(KEYINPUT82), .B(KEYINPUT63), .Z(n644) );
  XNOR2_X1 U717 ( .A(n645), .B(n644), .ZN(G57) );
  XNOR2_X1 U718 ( .A(n647), .B(G131), .ZN(G33) );
  NAND2_X1 U719 ( .A1(n732), .A2(G469), .ZN(n651) );
  XOR2_X1 U720 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n648) );
  XNOR2_X1 U721 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U722 ( .A(n651), .B(n650), .ZN(n652) );
  NOR2_X1 U723 ( .A1(n652), .A2(n736), .ZN(G54) );
  XNOR2_X1 U724 ( .A(G101), .B(n653), .ZN(G3) );
  NOR2_X1 U725 ( .A1(n657), .A2(n673), .ZN(n654) );
  XOR2_X1 U726 ( .A(G104), .B(n654), .Z(G6) );
  XOR2_X1 U727 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n656) );
  XNOR2_X1 U728 ( .A(G107), .B(KEYINPUT108), .ZN(n655) );
  XNOR2_X1 U729 ( .A(n656), .B(n655), .ZN(n659) );
  NOR2_X1 U730 ( .A1(n657), .A2(n677), .ZN(n658) );
  XOR2_X1 U731 ( .A(n659), .B(n658), .Z(G9) );
  INV_X1 U732 ( .A(n660), .ZN(n664) );
  NAND2_X1 U733 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U734 ( .A1(n664), .A2(n663), .ZN(n668) );
  XOR2_X1 U735 ( .A(KEYINPUT111), .B(KEYINPUT29), .Z(n666) );
  XNOR2_X1 U736 ( .A(G128), .B(KEYINPUT110), .ZN(n665) );
  XNOR2_X1 U737 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U738 ( .A(n668), .B(n667), .ZN(G30) );
  XNOR2_X1 U739 ( .A(G143), .B(n669), .ZN(G45) );
  AND2_X1 U740 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U741 ( .A(G146), .B(n672), .Z(G48) );
  NOR2_X1 U742 ( .A1(n673), .A2(n676), .ZN(n674) );
  XOR2_X1 U743 ( .A(KEYINPUT112), .B(n674), .Z(n675) );
  XNOR2_X1 U744 ( .A(G113), .B(n675), .ZN(G15) );
  NOR2_X1 U745 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U746 ( .A(G116), .B(n678), .Z(G18) );
  XOR2_X1 U747 ( .A(KEYINPUT113), .B(KEYINPUT37), .Z(n681) );
  XOR2_X1 U748 ( .A(G125), .B(n679), .Z(n680) );
  XNOR2_X1 U749 ( .A(n681), .B(n680), .ZN(G27) );
  XOR2_X1 U750 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n730) );
  AND2_X1 U751 ( .A1(n682), .A2(n620), .ZN(n683) );
  NOR2_X1 U752 ( .A1(n684), .A2(n683), .ZN(n728) );
  NAND2_X1 U753 ( .A1(G952), .A2(n685), .ZN(n719) );
  XOR2_X1 U754 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n700) );
  NOR2_X1 U755 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U756 ( .A(KEYINPUT49), .B(n688), .ZN(n694) );
  NAND2_X1 U757 ( .A1(n690), .A2(n374), .ZN(n691) );
  XNOR2_X1 U758 ( .A(n691), .B(KEYINPUT114), .ZN(n692) );
  XNOR2_X1 U759 ( .A(KEYINPUT50), .B(n692), .ZN(n693) );
  NAND2_X1 U760 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U761 ( .A1(n695), .A2(n599), .ZN(n697) );
  NOR2_X1 U762 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U763 ( .A(n698), .B(KEYINPUT115), .ZN(n699) );
  XNOR2_X1 U764 ( .A(n700), .B(n699), .ZN(n701) );
  NAND2_X1 U765 ( .A1(n721), .A2(n701), .ZN(n702) );
  XNOR2_X1 U766 ( .A(KEYINPUT117), .B(n702), .ZN(n716) );
  NOR2_X1 U767 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U768 ( .A1(n707), .A2(n706), .ZN(n712) );
  INV_X1 U769 ( .A(n708), .ZN(n710) );
  NOR2_X1 U770 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U771 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U772 ( .A1(n722), .A2(n713), .ZN(n714) );
  XNOR2_X1 U773 ( .A(n714), .B(KEYINPUT118), .ZN(n715) );
  NOR2_X1 U774 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U775 ( .A(n717), .B(KEYINPUT52), .ZN(n718) );
  NOR2_X1 U776 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U777 ( .A(n720), .B(KEYINPUT119), .ZN(n726) );
  INV_X1 U778 ( .A(n721), .ZN(n723) );
  NOR2_X1 U779 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U780 ( .A1(n724), .A2(n403), .ZN(n725) );
  NAND2_X1 U781 ( .A1(n726), .A2(n725), .ZN(n727) );
  OR2_X1 U782 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U783 ( .A(n730), .B(n729), .ZN(G75) );
  BUF_X1 U784 ( .A(n387), .Z(n732) );
  NAND2_X1 U785 ( .A1(n732), .A2(G478), .ZN(n734) );
  XNOR2_X1 U786 ( .A(n734), .B(n733), .ZN(n735) );
  NOR2_X1 U787 ( .A1(n736), .A2(n735), .ZN(G63) );
  NOR2_X1 U788 ( .A1(n737), .A2(n403), .ZN(n742) );
  NAND2_X1 U789 ( .A1(n403), .A2(G224), .ZN(n738) );
  XNOR2_X1 U790 ( .A(KEYINPUT61), .B(n738), .ZN(n739) );
  NAND2_X1 U791 ( .A1(n739), .A2(G898), .ZN(n740) );
  XNOR2_X1 U792 ( .A(n740), .B(KEYINPUT123), .ZN(n741) );
  NOR2_X1 U793 ( .A1(n742), .A2(n741), .ZN(n750) );
  BUF_X1 U794 ( .A(n743), .Z(n744) );
  XNOR2_X1 U795 ( .A(n744), .B(G101), .ZN(n747) );
  NOR2_X1 U796 ( .A1(G898), .A2(n745), .ZN(n746) );
  NOR2_X1 U797 ( .A1(n747), .A2(n746), .ZN(n748) );
  XOR2_X1 U798 ( .A(KEYINPUT124), .B(n748), .Z(n749) );
  XNOR2_X1 U799 ( .A(n750), .B(n749), .ZN(G69) );
  XOR2_X1 U800 ( .A(n388), .B(n751), .Z(n756) );
  XNOR2_X1 U801 ( .A(n428), .B(n756), .ZN(n754) );
  NOR2_X1 U802 ( .A1(n754), .A2(n403), .ZN(n755) );
  XNOR2_X1 U803 ( .A(KEYINPUT125), .B(n755), .ZN(n760) );
  XOR2_X1 U804 ( .A(G227), .B(n756), .Z(n757) );
  NAND2_X1 U805 ( .A1(n757), .A2(G900), .ZN(n758) );
  NAND2_X1 U806 ( .A1(n758), .A2(n403), .ZN(n759) );
  NAND2_X1 U807 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U808 ( .A(KEYINPUT126), .B(n761), .ZN(G72) );
  XNOR2_X1 U809 ( .A(G137), .B(KEYINPUT127), .ZN(n763) );
  XNOR2_X1 U810 ( .A(n763), .B(n762), .ZN(G39) );
endmodule

