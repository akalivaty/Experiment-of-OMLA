//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n566, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n580, new_n581, new_n582,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n628, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1164;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT67), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT68), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G237), .A2(G236), .A3(G235), .A4(G238), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT69), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n456), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(new_n453), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  INV_X1    g041(.A(G113), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  OAI22_X1  g043(.A1(new_n465), .A2(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n468), .A2(G2105), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n469), .A2(G2105), .B1(G101), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n473), .B1(new_n463), .B2(new_n464), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT70), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n477), .A2(KEYINPUT70), .A3(new_n473), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n471), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n477), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n465), .A2(G2105), .ZN(new_n484));
  AOI22_X1  g059(.A1(new_n483), .A2(G124), .B1(new_n484), .B2(G136), .ZN(new_n485));
  INV_X1    g060(.A(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(KEYINPUT71), .B1(G100), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NOR3_X1   g063(.A1(KEYINPUT71), .A2(G100), .A3(G2105), .ZN(new_n489));
  OAI221_X1 g064(.A(G2104), .B1(G112), .B2(new_n486), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n485), .A2(new_n490), .ZN(G162));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(KEYINPUT73), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n493), .B(new_n495), .C1(new_n464), .C2(new_n463), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n497), .B(G2104), .C1(G114), .C2(new_n486), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT73), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n494), .A2(KEYINPUT73), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n503), .B1(new_n477), .B2(new_n493), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  AND2_X1   g080(.A1(G126), .A2(G2105), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n477), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g084(.A(KEYINPUT72), .B(new_n506), .C1(new_n463), .C2(new_n464), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  OR2_X1    g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT74), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n520), .B1(new_n518), .B2(KEYINPUT6), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n522), .A2(KEYINPUT74), .A3(G651), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n521), .A2(new_n523), .B1(KEYINPUT6), .B2(new_n518), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n524), .A2(G88), .A3(new_n516), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n521), .A2(new_n523), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n518), .A2(KEYINPUT6), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n526), .A2(G50), .A3(G543), .A4(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT75), .ZN(new_n529));
  AND3_X1   g104(.A1(new_n525), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n529), .B1(new_n525), .B2(new_n528), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n519), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(G166));
  NAND2_X1  g108(.A1(new_n524), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G51), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n526), .A2(new_n527), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n514), .A2(new_n515), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G89), .ZN(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(KEYINPUT7), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(KEYINPUT7), .ZN(new_n543));
  AND2_X1   g118(.A1(G63), .A2(G651), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n542), .A2(new_n543), .B1(new_n516), .B2(new_n544), .ZN(new_n545));
  AND3_X1   g120(.A1(new_n536), .A2(new_n540), .A3(new_n545), .ZN(G168));
  XOR2_X1   g121(.A(KEYINPUT76), .B(G52), .Z(new_n547));
  NAND2_X1  g122(.A1(new_n535), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n539), .A2(G90), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n518), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G56), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n538), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G651), .ZN(new_n557));
  XOR2_X1   g132(.A(KEYINPUT77), .B(G43), .Z(new_n558));
  NAND3_X1  g133(.A1(new_n524), .A2(G543), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n524), .A2(G81), .A3(new_n516), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n557), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(new_n563));
  XOR2_X1   g138(.A(new_n563), .B(KEYINPUT78), .Z(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g140(.A(KEYINPUT79), .B(KEYINPUT8), .Z(new_n566));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n566), .B(new_n567), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  XOR2_X1   g144(.A(KEYINPUT80), .B(KEYINPUT9), .Z(new_n570));
  NAND3_X1  g145(.A1(new_n535), .A2(G53), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n539), .A2(G91), .ZN(new_n572));
  NOR2_X1   g147(.A1(KEYINPUT80), .A2(KEYINPUT9), .ZN(new_n573));
  INV_X1    g148(.A(G53), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n534), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n516), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n576), .A2(new_n518), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n571), .A2(new_n572), .A3(new_n575), .A4(new_n577), .ZN(G299));
  INV_X1    g153(.A(G168), .ZN(G286));
  NAND2_X1  g154(.A1(new_n532), .A2(KEYINPUT81), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT81), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n581), .B(new_n519), .C1(new_n530), .C2(new_n531), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n580), .A2(new_n582), .ZN(G303));
  NAND4_X1  g158(.A1(new_n526), .A2(G87), .A3(new_n516), .A4(new_n527), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT82), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n524), .A2(KEYINPUT82), .A3(G87), .A4(new_n516), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n526), .A2(G49), .A3(G543), .A4(new_n527), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n586), .A2(new_n587), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(KEYINPUT83), .ZN(new_n591));
  AND2_X1   g166(.A1(new_n588), .A2(new_n589), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT83), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n592), .A2(new_n593), .A3(new_n587), .A4(new_n586), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G288));
  NAND3_X1  g171(.A1(new_n524), .A2(G86), .A3(new_n516), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n524), .A2(G48), .A3(G543), .ZN(new_n598));
  INV_X1    g173(.A(G61), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n599), .B1(new_n514), .B2(new_n515), .ZN(new_n600));
  AND2_X1   g175(.A1(G73), .A2(G543), .ZN(new_n601));
  OAI21_X1  g176(.A(G651), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n597), .A2(new_n598), .A3(new_n602), .ZN(G305));
  NAND2_X1  g178(.A1(new_n535), .A2(G47), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n539), .A2(G85), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n606));
  OAI211_X1 g181(.A(new_n604), .B(new_n605), .C1(new_n518), .C2(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(G301), .A2(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(G79), .A2(G543), .ZN(new_n609));
  INV_X1    g184(.A(G66), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n538), .B2(new_n610), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n535), .A2(G54), .B1(new_n611), .B2(G651), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  NAND4_X1  g188(.A1(new_n526), .A2(G92), .A3(new_n516), .A4(new_n527), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n614), .A2(KEYINPUT84), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(KEYINPUT84), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(KEYINPUT10), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT10), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n615), .A2(new_n619), .A3(new_n616), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n613), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n608), .B1(new_n621), .B2(G868), .ZN(G284));
  OAI21_X1  g197(.A(new_n608), .B1(new_n621), .B2(G868), .ZN(G321));
  NAND2_X1  g198(.A1(G286), .A2(G868), .ZN(new_n624));
  INV_X1    g199(.A(G299), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(G297));
  OAI21_X1  g201(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(G280));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n621), .B1(new_n628), .B2(G860), .ZN(G148));
  NAND2_X1  g204(.A1(new_n621), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G868), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(G868), .B2(new_n562), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n483), .A2(G123), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n484), .A2(G135), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n486), .A2(G111), .ZN(new_n636));
  OAI21_X1  g211(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n634), .B(new_n635), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT86), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n640), .A2(G2096), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n477), .A2(new_n470), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT12), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2100), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT85), .B(KEYINPUT13), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n640), .A2(G2096), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n641), .A2(new_n646), .A3(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(G2427), .B(G2430), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT88), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT87), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n652), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(KEYINPUT14), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  XOR2_X1   g234(.A(G1341), .B(G1348), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2443), .B(G2446), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n657), .A2(new_n661), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(G14), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n663), .B1(new_n662), .B2(new_n664), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(G401));
  XOR2_X1   g243(.A(KEYINPUT89), .B(KEYINPUT17), .Z(new_n669));
  XNOR2_X1  g244(.A(G2072), .B(G2078), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2067), .B(G2678), .ZN(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n671), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n674), .B1(new_n672), .B2(new_n670), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n671), .B2(new_n672), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n673), .A2(new_n672), .A3(new_n670), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT18), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n675), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G2096), .B(G2100), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G227));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT19), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1956), .B(G2474), .Z(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  AND2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT90), .B(KEYINPUT20), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n686), .A2(new_n687), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  MUX2_X1   g268(.A(new_n693), .B(new_n692), .S(new_n685), .Z(new_n694));
  NOR2_X1   g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1991), .B(G1996), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1981), .B(G1986), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(G229));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G21), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G168), .B2(new_n703), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n705), .A2(G1966), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT102), .Z(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(G1966), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT100), .ZN(new_n709));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  OR3_X1    g285(.A1(new_n640), .A2(KEYINPUT101), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(KEYINPUT101), .B1(new_n640), .B2(new_n710), .ZN(new_n712));
  INV_X1    g287(.A(G28), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n713), .A2(KEYINPUT30), .ZN(new_n714));
  AOI21_X1  g289(.A(G29), .B1(new_n713), .B2(KEYINPUT30), .ZN(new_n715));
  OR2_X1    g290(.A1(KEYINPUT31), .A2(G11), .ZN(new_n716));
  NAND2_X1  g291(.A1(KEYINPUT31), .A2(G11), .ZN(new_n717));
  AOI22_X1  g292(.A1(new_n714), .A2(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n711), .A2(new_n712), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(G5), .A2(G16), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT103), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G301), .B2(new_n703), .ZN(new_n722));
  INV_X1    g297(.A(G1961), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OR4_X1    g299(.A1(new_n707), .A2(new_n709), .A3(new_n719), .A4(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(KEYINPUT104), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n710), .A2(G32), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n484), .A2(G141), .B1(G105), .B2(new_n470), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n483), .A2(G129), .ZN(new_n729));
  NAND3_X1  g304(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT26), .Z(new_n731));
  NAND3_X1  g306(.A1(new_n728), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n727), .B1(new_n733), .B2(new_n710), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT27), .ZN(new_n735));
  INV_X1    g310(.A(G1996), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n484), .A2(G140), .ZN(new_n738));
  OR2_X1    g313(.A1(G104), .A2(G2105), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n739), .B(G2104), .C1(G116), .C2(new_n486), .ZN(new_n740));
  INV_X1    g315(.A(G128), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n738), .B(new_n740), .C1(new_n741), .C2(new_n482), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G29), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n710), .A2(G26), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT28), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G2067), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n710), .A2(G35), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G162), .B2(new_n710), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT29), .B(G2090), .Z(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G27), .A2(G29), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G164), .B2(G29), .ZN(new_n754));
  INV_X1    g329(.A(G2078), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n748), .A2(new_n752), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n703), .A2(G19), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT98), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n562), .B2(new_n703), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1341), .ZN(new_n761));
  NOR3_X1   g336(.A1(new_n737), .A2(new_n757), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n710), .A2(G33), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n486), .A2(G103), .A3(G2104), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT25), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n484), .A2(G139), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n486), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT99), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n763), .B1(new_n771), .B2(new_n710), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G2072), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT24), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(G34), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(G34), .ZN(new_n776));
  AOI21_X1  g351(.A(G29), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n480), .B2(G29), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G2084), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n773), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n772), .A2(G2072), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n703), .A2(G20), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT23), .Z(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G299), .B2(G16), .ZN(new_n784));
  INV_X1    g359(.A(G1956), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n722), .A2(new_n723), .ZN(new_n787));
  NOR4_X1   g362(.A1(new_n780), .A2(new_n781), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n703), .A2(G4), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n621), .B2(new_n703), .ZN(new_n790));
  INV_X1    g365(.A(G1348), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n726), .A2(new_n762), .A3(new_n788), .A4(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n725), .A2(KEYINPUT104), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT36), .ZN(new_n796));
  INV_X1    g371(.A(G25), .ZN(new_n797));
  OR3_X1    g372(.A1(new_n797), .A2(KEYINPUT91), .A3(G29), .ZN(new_n798));
  OAI21_X1  g373(.A(KEYINPUT91), .B1(new_n797), .B2(G29), .ZN(new_n799));
  OAI21_X1  g374(.A(KEYINPUT93), .B1(G95), .B2(G2105), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  NOR3_X1   g376(.A1(KEYINPUT93), .A2(G95), .A3(G2105), .ZN(new_n802));
  OAI221_X1 g377(.A(G2104), .B1(G107), .B2(new_n486), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT94), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n484), .A2(G131), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT92), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n483), .A2(G119), .ZN(new_n807));
  AND3_X1   g382(.A1(new_n804), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n798), .B(new_n799), .C1(new_n808), .C2(new_n710), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT35), .B(G1991), .Z(new_n810));
  XOR2_X1   g385(.A(new_n809), .B(new_n810), .Z(new_n811));
  MUX2_X1   g386(.A(G24), .B(G290), .S(G16), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1986), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT95), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n592), .A2(KEYINPUT95), .A3(new_n587), .A4(new_n586), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  MUX2_X1   g393(.A(G23), .B(new_n818), .S(G16), .Z(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT33), .B(G1976), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  OR2_X1    g396(.A1(G6), .A2(G16), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G305), .B2(new_n703), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT32), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(G1981), .ZN(new_n825));
  NOR2_X1   g400(.A1(G16), .A2(G22), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(G166), .B2(G16), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT96), .B(G1971), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n821), .A2(new_n825), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n814), .B1(new_n830), .B2(KEYINPUT34), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(KEYINPUT97), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT97), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n814), .B(new_n833), .C1(KEYINPUT34), .C2(new_n830), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n830), .A2(KEYINPUT34), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n796), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n835), .A2(new_n796), .A3(new_n836), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n795), .B1(new_n838), .B2(new_n839), .ZN(G311));
  NOR2_X1   g415(.A1(new_n793), .A2(new_n794), .ZN(new_n841));
  INV_X1    g416(.A(new_n839), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n842), .B2(new_n837), .ZN(G150));
  NAND2_X1  g418(.A1(new_n621), .A2(G559), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT38), .Z(new_n845));
  NAND2_X1  g420(.A1(G80), .A2(G543), .ZN(new_n846));
  INV_X1    g421(.A(G67), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n846), .B1(new_n538), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G651), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n524), .A2(G93), .A3(new_n516), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n524), .A2(G55), .A3(G543), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n561), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n561), .A2(new_n852), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n845), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT39), .ZN(new_n858));
  AOI21_X1  g433(.A(G860), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n859), .B1(new_n858), .B2(new_n857), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n852), .A2(G860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT37), .Z(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(G145));
  XNOR2_X1  g438(.A(new_n512), .B(new_n742), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n732), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(new_n770), .ZN(new_n866));
  INV_X1    g441(.A(new_n771), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n866), .B1(new_n867), .B2(new_n865), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n484), .A2(G142), .ZN(new_n869));
  OAI21_X1  g444(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT105), .ZN(new_n871));
  INV_X1    g446(.A(G118), .ZN(new_n872));
  AOI22_X1  g447(.A1(new_n870), .A2(new_n871), .B1(new_n872), .B2(G2105), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n871), .B2(new_n870), .ZN(new_n874));
  INV_X1    g449(.A(G130), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n869), .B(new_n874), .C1(new_n875), .C2(new_n482), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT106), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n643), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n808), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n868), .B(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n640), .B(G162), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(G160), .ZN(new_n882));
  AOI21_X1  g457(.A(G37), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(new_n882), .B2(new_n880), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT40), .ZN(G395));
  AND3_X1   g460(.A1(new_n615), .A2(new_n619), .A3(new_n616), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n619), .B1(new_n615), .B2(new_n616), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n612), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT107), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(new_n889), .A3(new_n625), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n621), .A2(G299), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n889), .B1(new_n888), .B2(new_n625), .ZN(new_n893));
  OAI21_X1  g468(.A(KEYINPUT41), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n630), .B(new_n856), .ZN(new_n895));
  OAI21_X1  g470(.A(KEYINPUT107), .B1(new_n621), .B2(G299), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n896), .A2(new_n897), .A3(new_n891), .A4(new_n890), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n894), .A2(new_n895), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n896), .A2(new_n891), .A3(new_n890), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n899), .B1(new_n895), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT108), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT42), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n818), .B(G166), .ZN(new_n907));
  XOR2_X1   g482(.A(G290), .B(G305), .Z(new_n908));
  XNOR2_X1  g483(.A(new_n907), .B(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n910), .B1(new_n903), .B2(new_n904), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n902), .A2(new_n905), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n906), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n911), .B1(new_n906), .B2(new_n912), .ZN(new_n914));
  OAI21_X1  g489(.A(G868), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n915), .B1(G868), .B2(new_n916), .ZN(G295));
  OAI21_X1  g492(.A(new_n915), .B1(G868), .B2(new_n916), .ZN(G331));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT43), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n854), .A2(new_n855), .A3(G171), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n562), .A2(new_n916), .ZN(new_n922));
  AOI21_X1  g497(.A(G301), .B1(new_n922), .B2(new_n853), .ZN(new_n923));
  OAI21_X1  g498(.A(G286), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(G171), .B1(new_n854), .B2(new_n855), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n922), .A2(G301), .A3(new_n853), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(G168), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n900), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n921), .A2(new_n923), .A3(G286), .ZN(new_n932));
  AOI21_X1  g507(.A(G168), .B1(new_n925), .B2(new_n926), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n934), .A2(new_n894), .A3(new_n898), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n928), .A2(KEYINPUT109), .A3(new_n900), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n931), .A2(new_n935), .A3(new_n909), .A4(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(G37), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n931), .A2(new_n935), .A3(new_n936), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n910), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n920), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n935), .A2(new_n929), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n910), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n944), .A2(new_n937), .A3(new_n938), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n919), .B1(new_n942), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n941), .A2(new_n920), .A3(new_n938), .A4(new_n937), .ZN(new_n949));
  AND4_X1   g524(.A1(KEYINPUT110), .A2(new_n948), .A3(KEYINPUT44), .A4(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n919), .B1(new_n945), .B2(KEYINPUT43), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT110), .B1(new_n951), .B2(new_n949), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n947), .B1(new_n950), .B2(new_n952), .ZN(G397));
  OR2_X1    g528(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n954));
  NAND2_X1  g529(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n466), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n467), .A2(new_n468), .ZN(new_n957));
  OAI21_X1  g532(.A(G2105), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n470), .A2(G101), .ZN(new_n959));
  XOR2_X1   g534(.A(KEYINPUT111), .B(G40), .Z(new_n960));
  NAND4_X1  g535(.A1(new_n479), .A2(new_n958), .A3(new_n959), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT112), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n471), .A2(new_n963), .A3(new_n479), .A4(new_n960), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(G1384), .B1(new_n505), .B2(new_n511), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n965), .A2(KEYINPUT45), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n967), .A2(G1996), .A3(new_n732), .ZN(new_n968));
  XOR2_X1   g543(.A(new_n968), .B(KEYINPUT113), .Z(new_n969));
  INV_X1    g544(.A(G2067), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n742), .B(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n971), .B1(G1996), .B2(new_n732), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n967), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n808), .B(new_n810), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n974), .B1(new_n967), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(G290), .A2(G1986), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n967), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT48), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  AND4_X1   g555(.A1(new_n810), .A2(new_n969), .A3(new_n808), .A4(new_n973), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n742), .A2(G2067), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n967), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n967), .A2(new_n736), .ZN(new_n984));
  XOR2_X1   g559(.A(new_n984), .B(KEYINPUT46), .Z(new_n985));
  NAND2_X1  g560(.A1(new_n971), .A2(new_n733), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n967), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT125), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n989), .B(new_n990), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n980), .A2(new_n983), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT50), .ZN(new_n993));
  AOI22_X1  g568(.A1(new_n962), .A2(new_n964), .B1(new_n966), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT115), .B1(new_n966), .B2(new_n993), .ZN(new_n995));
  INV_X1    g570(.A(G1384), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT72), .B1(new_n477), .B2(new_n506), .ZN(new_n997));
  INV_X1    g572(.A(new_n510), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n486), .A2(G138), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n1000), .B1(new_n954), .B2(new_n955), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n496), .B(new_n498), .C1(new_n1001), .C2(new_n503), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n996), .B1(new_n999), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT115), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(new_n1004), .A3(KEYINPUT50), .ZN(new_n1005));
  XNOR2_X1  g580(.A(KEYINPUT117), .B(G2084), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n994), .A2(new_n995), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1966), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1009), .A2(G1384), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(new_n999), .B2(new_n1002), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1011), .B1(new_n966), .B2(KEYINPUT45), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1008), .B1(new_n965), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1007), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(G8), .B1(new_n1014), .B2(G286), .ZN(new_n1015));
  AOI21_X1  g590(.A(G168), .B1(new_n1007), .B2(new_n1013), .ZN(new_n1016));
  OAI21_X1  g591(.A(KEYINPUT51), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1018), .B(G8), .C1(new_n1014), .C2(G286), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT62), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n962), .A2(new_n964), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n966), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n816), .A2(G1976), .A3(new_n817), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1023), .A2(G8), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G305), .A2(G1981), .ZN(new_n1026));
  INV_X1    g601(.A(G1981), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n598), .A2(new_n597), .A3(new_n1027), .A4(new_n602), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n1026), .A2(KEYINPUT49), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT49), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G8), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1032), .B1(new_n1022), .B2(new_n966), .ZN(new_n1033));
  AOI22_X1  g608(.A1(new_n1025), .A2(KEYINPUT52), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n1035));
  INV_X1    g610(.A(G1976), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n591), .A2(new_n1036), .A3(new_n594), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1035), .B1(new_n1025), .B2(new_n1039), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1041), .A2(KEYINPUT116), .A3(new_n1033), .A4(new_n1024), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n1034), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n1011), .A2(KEYINPUT114), .B1(new_n1003), .B2(new_n1009), .ZN(new_n1044));
  OR2_X1    g619(.A1(new_n1011), .A2(KEYINPUT114), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(new_n1022), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G1971), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G2090), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n994), .A2(new_n1049), .A3(new_n995), .A4(new_n1005), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1032), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n580), .A2(G8), .A3(new_n582), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n580), .A2(KEYINPUT55), .A3(G8), .A4(new_n582), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1051), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n966), .A2(new_n993), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1003), .A2(KEYINPUT50), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1022), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1049), .A2(new_n1060), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1054), .B(new_n1055), .C1(new_n1061), .C2(new_n1032), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1043), .A2(new_n1057), .A3(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n995), .A2(new_n1022), .A3(new_n1058), .A4(new_n1005), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT120), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n994), .A2(KEYINPUT120), .A3(new_n995), .A4(new_n1005), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1066), .A2(new_n723), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(new_n1046), .B2(G2078), .ZN(new_n1070));
  OR4_X1    g645(.A1(new_n1069), .A2(new_n965), .A3(new_n1012), .A4(G2078), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(G171), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1063), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT62), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1017), .A2(new_n1075), .A3(new_n1019), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1021), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  AOI211_X1 g652(.A(new_n1032), .B(G286), .C1(new_n1007), .C2(new_n1013), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1043), .A2(new_n1078), .A3(new_n1062), .A4(new_n1057), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT63), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1051), .A2(new_n1056), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1034), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT118), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1057), .A2(KEYINPUT63), .A3(new_n1078), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n1082), .A2(new_n1083), .A3(KEYINPUT118), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1081), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1083), .A2(new_n1057), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1090), .A2(new_n1036), .A3(new_n595), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n1028), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1089), .B1(new_n1033), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1077), .A2(new_n1088), .A3(new_n1093), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n755), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1044), .A2(new_n1045), .A3(G160), .A4(new_n1095), .ZN(new_n1096));
  AND4_X1   g671(.A1(G301), .A2(new_n1068), .A3(new_n1070), .A4(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT123), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT54), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1068), .A2(G301), .A3(new_n1070), .A4(new_n1096), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1073), .A2(KEYINPUT123), .A3(new_n1100), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1099), .A2(KEYINPUT124), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT124), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1068), .A2(new_n1071), .A3(G301), .A4(new_n1070), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1068), .A2(new_n1070), .A3(new_n1096), .ZN(new_n1105));
  OAI211_X1 g680(.A(KEYINPUT54), .B(new_n1104), .C1(new_n1105), .C2(G301), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1043), .A2(new_n1057), .A3(new_n1062), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(new_n1107), .A3(new_n1020), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1102), .A2(new_n1103), .A3(new_n1108), .ZN(new_n1109));
  XOR2_X1   g684(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1110));
  XOR2_X1   g685(.A(KEYINPUT58), .B(G1341), .Z(new_n1111));
  NAND2_X1  g686(.A1(new_n1023), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1044), .A2(new_n1045), .A3(new_n1022), .A4(new_n736), .ZN(new_n1113));
  AOI211_X1 g688(.A(new_n561), .B(new_n1110), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n562), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1117), .A2(KEYINPUT59), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1114), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1022), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n785), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT56), .B(G2072), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1044), .A2(new_n1045), .A3(new_n1022), .A4(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1125));
  XNOR2_X1  g700(.A(G299), .B(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT61), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1121), .A2(new_n1126), .A3(new_n1123), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1129), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1119), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(KEYINPUT122), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1066), .A2(new_n791), .A3(new_n1067), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1022), .A2(new_n970), .A3(new_n966), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT60), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n621), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1135), .A2(KEYINPUT60), .A3(new_n888), .A4(new_n1136), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1119), .B(new_n1144), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1134), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1130), .A2(new_n621), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1147), .A2(new_n1137), .B1(new_n1127), .B2(new_n1124), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1094), .B1(new_n1109), .B2(new_n1149), .ZN(new_n1150));
  AND2_X1   g725(.A1(G290), .A2(G1986), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n967), .B1(new_n977), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n976), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n992), .B1(new_n1150), .B2(new_n1153), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g729(.A1(G227), .A2(new_n461), .ZN(new_n1156));
  OAI21_X1  g730(.A(new_n1156), .B1(new_n666), .B2(new_n667), .ZN(new_n1157));
  NAND2_X1  g731(.A1(new_n1157), .A2(KEYINPUT127), .ZN(new_n1158));
  OR2_X1    g732(.A1(new_n1157), .A2(KEYINPUT127), .ZN(new_n1159));
  AND2_X1   g733(.A1(new_n1159), .A2(new_n701), .ZN(new_n1160));
  NAND3_X1  g734(.A1(new_n884), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  NOR2_X1   g735(.A1(new_n942), .A2(new_n946), .ZN(new_n1162));
  NOR2_X1   g736(.A1(new_n1161), .A2(new_n1162), .ZN(G308));
  AND2_X1   g737(.A1(new_n1160), .A2(new_n1158), .ZN(new_n1164));
  OAI211_X1 g738(.A(new_n1164), .B(new_n884), .C1(new_n942), .C2(new_n946), .ZN(G225));
endmodule


