//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 0 0 0 1 0 0 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n187));
  INV_X1    g001(.A(G116), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT68), .A2(G116), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(G119), .A3(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G116), .ZN(new_n193));
  INV_X1    g007(.A(G113), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT2), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G113), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n191), .A2(new_n193), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT69), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n191), .A2(new_n198), .A3(KEYINPUT69), .A4(new_n193), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT67), .ZN(new_n204));
  AND3_X1   g018(.A1(new_n195), .A2(new_n197), .A3(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n204), .B1(new_n195), .B2(new_n197), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n191), .A2(new_n193), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n203), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G104), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT3), .B1(new_n211), .B2(G107), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT3), .ZN(new_n213));
  INV_X1    g027(.A(G107), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(G104), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n211), .A2(G107), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n212), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G101), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT82), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G101), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n212), .A2(new_n215), .A3(new_n221), .A4(new_n216), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n222), .A2(KEYINPUT4), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n217), .A2(KEYINPUT82), .A3(G101), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n220), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT4), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n217), .A2(new_n226), .A3(G101), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n210), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n191), .A2(KEYINPUT5), .A3(new_n193), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n193), .A2(KEYINPUT5), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(new_n194), .ZN(new_n231));
  AOI22_X1  g045(.A1(new_n201), .A2(new_n202), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT83), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n211), .A2(G107), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n214), .A2(G104), .ZN(new_n235));
  OAI21_X1  g049(.A(G101), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n233), .B1(new_n222), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n222), .A2(new_n236), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(KEYINPUT83), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n232), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n228), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(G110), .B(G122), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n228), .A2(new_n242), .A3(new_n240), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(KEYINPUT6), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G146), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G143), .ZN(new_n248));
  INV_X1    g062(.A(G143), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G146), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  AND2_X1   g065(.A1(KEYINPUT65), .A2(G128), .ZN(new_n252));
  NOR2_X1   g066(.A1(KEYINPUT65), .A2(G128), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n255), .B1(G143), .B2(new_n247), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n251), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G125), .ZN(new_n258));
  XNOR2_X1  g072(.A(G143), .B(G146), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(new_n255), .A3(G128), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(KEYINPUT0), .A2(G128), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  XOR2_X1   g077(.A(KEYINPUT0), .B(G128), .Z(new_n264));
  OAI21_X1  g078(.A(new_n263), .B1(new_n259), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n261), .B1(new_n258), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT86), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT86), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n268), .B1(new_n265), .B2(new_n258), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G224), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n271), .A2(G953), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n272), .B(KEYINPUT87), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n270), .B(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n241), .A2(new_n275), .A3(new_n243), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n246), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT7), .B1(new_n271), .B2(G953), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n267), .A2(new_n269), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n266), .A2(new_n278), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n232), .A2(new_n238), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n242), .B(KEYINPUT8), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n284), .B1(new_n232), .B2(new_n238), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(G902), .B1(new_n287), .B2(new_n245), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n277), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(G210), .B1(G237), .B2(G902), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n277), .A2(new_n290), .A3(new_n288), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(KEYINPUT88), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n290), .B1(new_n277), .B2(new_n288), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT88), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G953), .ZN(new_n298));
  INV_X1    g112(.A(G952), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n299), .A2(KEYINPUT94), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n299), .A2(KEYINPUT94), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n302), .B1(G234), .B2(G237), .ZN(new_n303));
  AND2_X1   g117(.A1(KEYINPUT70), .A2(G953), .ZN(new_n304));
  NOR2_X1   g118(.A1(KEYINPUT70), .A2(G953), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G902), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n308), .B1(G234), .B2(G237), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n310), .B(KEYINPUT95), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT21), .B(G898), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n303), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n313), .B(KEYINPUT96), .ZN(new_n314));
  OAI21_X1  g128(.A(G214), .B1(G237), .B2(G902), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n294), .A2(new_n297), .A3(new_n314), .A4(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n306), .A2(G227), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(KEYINPUT81), .ZN(new_n318));
  XOR2_X1   g132(.A(G110), .B(G140), .Z(new_n319));
  XNOR2_X1  g133(.A(new_n318), .B(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n265), .A2(new_n227), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n225), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT10), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n324), .B1(new_n257), .B2(new_n260), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n325), .B1(new_n239), .B2(new_n237), .ZN(new_n326));
  INV_X1    g140(.A(G137), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n327), .A2(G134), .ZN(new_n328));
  INV_X1    g142(.A(G134), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT11), .B1(new_n329), .B2(G137), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT11), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(new_n327), .A3(G134), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n328), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G131), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n333), .B(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n248), .A2(KEYINPUT1), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n259), .B1(G128), .B2(new_n337), .ZN(new_n338));
  AND4_X1   g152(.A1(new_n255), .A2(new_n248), .A3(new_n250), .A4(G128), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n222), .B(new_n236), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n324), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n323), .A2(new_n326), .A3(new_n336), .A4(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  AOI22_X1  g157(.A1(new_n225), .A2(new_n322), .B1(new_n340), .B2(new_n324), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n336), .B1(new_n344), .B2(new_n326), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n321), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT12), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n238), .A2(new_n257), .A3(new_n260), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n340), .A2(new_n348), .A3(KEYINPUT84), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT84), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n238), .A2(new_n350), .A3(new_n257), .A4(new_n260), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n335), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n347), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n335), .A2(new_n351), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n340), .A2(new_n348), .A3(KEYINPUT84), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(KEYINPUT12), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n342), .A2(KEYINPUT85), .A3(new_n320), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT85), .B1(new_n342), .B2(new_n320), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n346), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G469), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n362), .A3(new_n308), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n349), .A2(new_n347), .A3(new_n352), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT12), .B1(new_n354), .B2(new_n355), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n342), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n342), .A2(new_n320), .ZN(new_n367));
  INV_X1    g181(.A(new_n345), .ZN(new_n368));
  AOI22_X1  g182(.A1(new_n366), .A2(new_n321), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G469), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n362), .A2(new_n308), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n363), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT9), .B(G234), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n374), .B(KEYINPUT79), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n308), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G221), .ZN(new_n377));
  XOR2_X1   g191(.A(new_n377), .B(KEYINPUT80), .Z(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n373), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT20), .ZN(new_n381));
  XNOR2_X1  g195(.A(G113), .B(G122), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(new_n211), .ZN(new_n383));
  OR2_X1    g197(.A1(KEYINPUT70), .A2(G953), .ZN(new_n384));
  INV_X1    g198(.A(G237), .ZN(new_n385));
  NAND2_X1  g199(.A1(KEYINPUT70), .A2(G953), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n384), .A2(G214), .A3(new_n385), .A4(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n249), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n306), .A2(G143), .A3(G214), .A4(new_n385), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT18), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n390), .B1(new_n391), .B2(new_n334), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n388), .A2(new_n389), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(KEYINPUT18), .A3(G131), .ZN(new_n394));
  INV_X1    g208(.A(G140), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G125), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n258), .A2(G140), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(G146), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n396), .A2(KEYINPUT76), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT76), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n395), .A3(G125), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n400), .A2(new_n402), .A3(new_n397), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n403), .A2(G146), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n392), .B(new_n394), .C1(new_n399), .C2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(KEYINPUT89), .B1(new_n393), .B2(G131), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT89), .ZN(new_n407));
  AOI211_X1 g221(.A(new_n407), .B(new_n334), .C1(new_n388), .C2(new_n389), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT17), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT92), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI211_X1 g225(.A(KEYINPUT92), .B(KEYINPUT17), .C1(new_n406), .C2(new_n408), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n403), .A2(KEYINPUT16), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT16), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n396), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(new_n247), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT77), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n413), .A2(new_n415), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G146), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n413), .A2(KEYINPUT77), .A3(new_n247), .A4(new_n415), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n418), .A2(new_n420), .A3(KEYINPUT91), .A4(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n411), .A2(new_n412), .A3(new_n422), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n418), .A2(new_n420), .A3(new_n421), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n407), .B1(new_n390), .B2(new_n334), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n393), .A2(KEYINPUT89), .A3(G131), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n390), .A2(new_n334), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  OAI22_X1  g242(.A1(new_n424), .A2(KEYINPUT91), .B1(new_n428), .B2(KEYINPUT17), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n383), .B(new_n405), .C1(new_n423), .C2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(KEYINPUT90), .B1(new_n398), .B2(KEYINPUT19), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n403), .A2(KEYINPUT19), .ZN(new_n432));
  MUX2_X1   g246(.A(KEYINPUT90), .B(new_n431), .S(new_n432), .Z(new_n433));
  OAI21_X1  g247(.A(new_n420), .B1(new_n433), .B2(G146), .ZN(new_n434));
  INV_X1    g248(.A(new_n428), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n405), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n383), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n430), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(G475), .A2(G902), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n381), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n440), .ZN(new_n442));
  AOI211_X1 g256(.A(KEYINPUT20), .B(new_n442), .C1(new_n430), .C2(new_n438), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n405), .B1(new_n423), .B2(new_n429), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n437), .ZN(new_n445));
  AOI21_X1  g259(.A(G902), .B1(new_n445), .B2(new_n430), .ZN(new_n446));
  INV_X1    g260(.A(G475), .ZN(new_n447));
  OAI22_X1  g261(.A1(new_n441), .A2(new_n443), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n253), .ZN(new_n449));
  NAND2_X1  g263(.A1(KEYINPUT65), .A2(G128), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(G143), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n249), .A2(G128), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n329), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(G134), .A3(new_n452), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT13), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n451), .A2(new_n456), .A3(G134), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n451), .A2(new_n456), .A3(G134), .A4(new_n452), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n189), .A2(G122), .A3(new_n190), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT93), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT93), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n189), .A2(new_n462), .A3(G122), .A4(new_n190), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n188), .A2(G122), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n214), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  AOI211_X1 g281(.A(G107), .B(new_n465), .C1(new_n461), .C2(new_n463), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n458), .B(new_n459), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n465), .B1(new_n464), .B2(KEYINPUT14), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT14), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n461), .A2(new_n471), .A3(new_n463), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n214), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n464), .A2(new_n214), .A3(new_n466), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(new_n454), .A3(new_n455), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n469), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n375), .A2(G217), .A3(new_n298), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n477), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n469), .B(new_n479), .C1(new_n473), .C2(new_n475), .ZN(new_n480));
  AOI21_X1  g294(.A(G902), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G478), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(KEYINPUT15), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  OR2_X1    g298(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n481), .A2(new_n484), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NOR4_X1   g301(.A1(new_n316), .A2(new_n380), .A3(new_n448), .A4(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n418), .A2(new_n420), .A3(new_n421), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n254), .A2(KEYINPUT23), .A3(G119), .ZN(new_n490));
  INV_X1    g304(.A(G128), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n491), .A2(G119), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT23), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT75), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n494), .B1(new_n192), .B2(G128), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT75), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n496), .B(KEYINPUT23), .C1(new_n491), .C2(G119), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n490), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n492), .B1(new_n254), .B2(G119), .ZN(new_n500));
  XOR2_X1   g314(.A(KEYINPUT24), .B(G110), .Z(new_n501));
  AOI22_X1  g315(.A1(new_n499), .A2(G110), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n489), .A2(new_n502), .ZN(new_n503));
  OAI22_X1  g317(.A1(new_n499), .A2(G110), .B1(new_n500), .B2(new_n501), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n399), .B1(new_n419), .B2(G146), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(KEYINPUT22), .B(G137), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(KEYINPUT78), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n306), .A2(G221), .A3(G234), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n503), .A2(new_n506), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n511), .B1(new_n503), .B2(new_n506), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(G217), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n515), .B1(G234), .B2(new_n308), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n516), .A2(G902), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n308), .B1(new_n512), .B2(new_n513), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT25), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g336(.A(KEYINPUT25), .B(new_n308), .C1(new_n512), .C2(new_n513), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n519), .B1(new_n524), .B2(new_n516), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  AOI211_X1 g340(.A(G131), .B(new_n328), .C1(new_n330), .C2(new_n332), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n330), .A2(new_n332), .ZN(new_n528));
  INV_X1    g342(.A(new_n328), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n334), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n265), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT64), .B1(new_n327), .B2(G134), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT64), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n329), .A3(G137), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n327), .A2(G134), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(G131), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n528), .A2(new_n334), .A3(new_n529), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT65), .B(G128), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n259), .B1(new_n337), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n537), .B(new_n538), .C1(new_n540), .C2(new_n339), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n531), .A2(KEYINPUT30), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n210), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT30), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT66), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n257), .A2(new_n260), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n547), .A2(KEYINPUT66), .A3(new_n537), .A4(new_n538), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n546), .A2(new_n548), .A3(new_n531), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n543), .B1(new_n544), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n201), .A2(new_n202), .B1(new_n207), .B2(new_n208), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(new_n541), .A3(new_n531), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n306), .A2(G210), .A3(new_n385), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT27), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT27), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n306), .A2(new_n555), .A3(G210), .A4(new_n385), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT26), .B(G101), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n554), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n557), .B1(new_n554), .B2(new_n556), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n552), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(KEYINPUT71), .B1(new_n550), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n549), .A2(new_n544), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n542), .A2(new_n210), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT71), .ZN(new_n566));
  INV_X1    g380(.A(new_n561), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n562), .A2(KEYINPUT31), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT72), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT72), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n562), .A2(new_n568), .A3(new_n571), .A4(KEYINPUT31), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n550), .A2(KEYINPUT31), .A3(new_n561), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n552), .A2(KEYINPUT28), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT28), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n551), .A2(new_n575), .A3(new_n541), .A4(new_n531), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n549), .A2(new_n210), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OR2_X1    g393(.A1(new_n558), .A2(new_n559), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(KEYINPUT73), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT73), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n574), .A2(new_n576), .B1(new_n549), .B2(new_n210), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n582), .B1(new_n583), .B2(new_n560), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n573), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n570), .A2(new_n572), .A3(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(G472), .A2(G902), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(KEYINPUT74), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(KEYINPUT32), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT32), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n586), .A2(new_n592), .A3(new_n589), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n531), .A2(new_n541), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n210), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n577), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n560), .A2(KEYINPUT29), .ZN(new_n598));
  INV_X1    g412(.A(new_n552), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n550), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n600), .A2(new_n560), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT29), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n602), .B1(new_n579), .B2(new_n580), .ZN(new_n603));
  OAI221_X1 g417(.A(new_n308), .B1(new_n597), .B2(new_n598), .C1(new_n601), .C2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(G472), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n526), .B1(new_n594), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n488), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT97), .B(G101), .Z(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G3));
  AND3_X1   g423(.A1(new_n525), .A2(new_n373), .A3(new_n379), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT98), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n586), .A2(new_n611), .A3(new_n308), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(G472), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n611), .B1(new_n586), .B2(new_n308), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n610), .B(new_n590), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(KEYINPUT99), .ZN(new_n616));
  INV_X1    g430(.A(new_n614), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n617), .A2(G472), .A3(new_n612), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT99), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n618), .A2(new_n619), .A3(new_n590), .A4(new_n610), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n482), .A2(new_n308), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n481), .B2(new_n482), .ZN(new_n622));
  INV_X1    g436(.A(new_n480), .ZN(new_n623));
  AND2_X1   g437(.A1(KEYINPUT68), .A2(G116), .ZN(new_n624));
  NOR2_X1   g438(.A1(KEYINPUT68), .A2(G116), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n462), .B1(new_n626), .B2(G122), .ZN(new_n627));
  INV_X1    g441(.A(new_n463), .ZN(new_n628));
  OAI21_X1  g442(.A(KEYINPUT14), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n629), .A2(new_n466), .A3(new_n472), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(G107), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n454), .A2(new_n455), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n468), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n479), .B1(new_n634), .B2(new_n469), .ZN(new_n635));
  OAI21_X1  g449(.A(KEYINPUT33), .B1(new_n623), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n478), .A2(new_n637), .A3(new_n480), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n636), .A2(G478), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n622), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT100), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT100), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n622), .A2(new_n639), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n448), .A2(new_n644), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n277), .A2(new_n290), .A3(new_n288), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n314), .B(new_n315), .C1(new_n646), .C2(new_n295), .ZN(new_n647));
  OAI21_X1  g461(.A(KEYINPUT101), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n647), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT101), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n649), .A2(new_n650), .A3(new_n448), .A4(new_n644), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n616), .A2(new_n620), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT34), .B(G104), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G6));
  NAND2_X1  g469(.A1(new_n616), .A2(new_n620), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n487), .B1(new_n446), .B2(new_n447), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n439), .A2(new_n440), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(KEYINPUT20), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n439), .A2(new_n381), .A3(new_n440), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n659), .A2(KEYINPUT102), .A3(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n662), .B1(new_n441), .B2(new_n443), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n657), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n664), .A2(new_n665), .A3(new_n649), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n665), .B1(new_n664), .B2(new_n649), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n656), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT35), .B(G107), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G9));
  NAND2_X1  g485(.A1(new_n503), .A2(new_n506), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n511), .A2(KEYINPUT36), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n674), .A2(new_n518), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(new_n524), .B2(new_n516), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n590), .B(new_n677), .C1(new_n613), .C2(new_n614), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT104), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n618), .A2(KEYINPUT104), .A3(new_n590), .A4(new_n677), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n680), .A2(new_n681), .A3(new_n488), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT37), .B(G110), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G12));
  AND3_X1   g498(.A1(new_n586), .A2(new_n592), .A3(new_n589), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n592), .B1(new_n586), .B2(new_n589), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n605), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(G900), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n303), .B1(new_n311), .B2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n315), .B1(new_n646), .B2(new_n295), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n380), .A2(new_n691), .A3(new_n676), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n687), .A2(new_n664), .A3(new_n690), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G128), .ZN(G30));
  NAND2_X1  g508(.A1(new_n342), .A2(new_n320), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT85), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(new_n357), .A3(new_n358), .ZN(new_n698));
  AOI21_X1  g512(.A(G902), .B1(new_n698), .B2(new_n346), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n371), .B1(new_n699), .B2(new_n362), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n378), .B1(new_n700), .B2(new_n370), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n689), .B(KEYINPUT39), .Z(new_n702));
  AND2_X1   g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(KEYINPUT40), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n685), .A2(new_n686), .ZN(new_n705));
  INV_X1    g519(.A(G472), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n562), .A2(new_n568), .ZN(new_n707));
  INV_X1    g521(.A(new_n596), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n580), .B1(new_n708), .B2(new_n599), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n706), .B1(new_n710), .B2(new_n308), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n705), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n294), .A2(new_n297), .ZN(new_n713));
  XOR2_X1   g527(.A(new_n713), .B(KEYINPUT38), .Z(new_n714));
  NAND2_X1  g528(.A1(new_n448), .A2(new_n487), .ZN(new_n715));
  INV_X1    g529(.A(new_n315), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n715), .A2(new_n716), .A3(new_n677), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n704), .A2(new_n712), .A3(new_n714), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G143), .ZN(G45));
  AND3_X1   g533(.A1(new_n448), .A2(new_n644), .A3(new_n690), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n687), .A2(new_n720), .A3(new_n692), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT105), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n687), .A2(new_n720), .A3(KEYINPUT105), .A4(new_n692), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G146), .ZN(G48));
  NAND2_X1  g540(.A1(new_n361), .A2(new_n308), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(G469), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n363), .A3(new_n377), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n687), .A2(new_n525), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n652), .ZN(new_n732));
  XNOR2_X1  g546(.A(KEYINPUT41), .B(G113), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G15));
  OAI21_X1  g548(.A(new_n731), .B1(new_n666), .B2(new_n667), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G116), .ZN(G18));
  INV_X1    g550(.A(new_n314), .ZN(new_n737));
  NOR4_X1   g551(.A1(new_n691), .A2(new_n729), .A3(new_n676), .A4(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n448), .ZN(new_n739));
  INV_X1    g553(.A(new_n486), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n481), .A2(new_n484), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n738), .A2(new_n687), .A3(new_n739), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G119), .ZN(G21));
  NOR2_X1   g558(.A1(new_n691), .A2(new_n729), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n745), .A2(new_n314), .A3(new_n448), .A4(new_n487), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n573), .B1(new_n580), .B2(new_n597), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n588), .B1(new_n747), .B2(new_n569), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n586), .A2(new_n308), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n748), .B1(new_n749), .B2(G472), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n525), .ZN(new_n751));
  OAI21_X1  g565(.A(KEYINPUT106), .B1(new_n746), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n706), .B1(new_n586), .B2(new_n308), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n526), .A2(new_n753), .A3(new_n748), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT106), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n448), .A2(new_n314), .A3(new_n487), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n754), .A2(new_n755), .A3(new_n756), .A4(new_n745), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n752), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g572(.A(KEYINPUT107), .B(G122), .Z(new_n759));
  XNOR2_X1  g573(.A(new_n758), .B(new_n759), .ZN(G24));
  NOR3_X1   g574(.A1(new_n753), .A2(new_n676), .A3(new_n748), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n720), .A2(new_n761), .A3(new_n745), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G125), .ZN(G27));
  INV_X1    g577(.A(new_n377), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT108), .B1(new_n369), .B2(G469), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n320), .B1(new_n357), .B2(new_n342), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n695), .A2(new_n345), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT108), .ZN(new_n768));
  NOR4_X1   g582(.A1(new_n766), .A2(new_n767), .A3(new_n768), .A4(new_n362), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n764), .B1(new_n770), .B2(new_n700), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n713), .A2(new_n315), .A3(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n772), .A2(new_n687), .A3(new_n525), .A4(new_n720), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT42), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n606), .A2(KEYINPUT42), .A3(new_n720), .A4(new_n772), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G131), .ZN(G33));
  AOI211_X1 g592(.A(new_n689), .B(new_n657), .C1(new_n661), .C2(new_n663), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n779), .A2(new_n772), .A3(new_n687), .A4(new_n525), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G134), .ZN(G36));
  AOI21_X1  g595(.A(new_n676), .B1(new_n618), .B2(new_n590), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n739), .A2(new_n644), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(KEYINPUT43), .ZN(new_n784));
  INV_X1    g598(.A(new_n644), .ZN(new_n785));
  OR3_X1    g599(.A1(new_n785), .A2(KEYINPUT43), .A3(new_n448), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n782), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT44), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n786), .A2(new_n784), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n790), .A2(KEYINPUT44), .A3(new_n782), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n369), .A2(KEYINPUT45), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n369), .A2(KEYINPUT45), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(G469), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n372), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT46), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n794), .A2(KEYINPUT46), .A3(new_n372), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n797), .A2(new_n363), .A3(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n799), .A2(new_n377), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n716), .B1(new_n294), .B2(new_n297), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n800), .A2(new_n702), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n789), .A2(new_n791), .A3(new_n802), .ZN(new_n803));
  XOR2_X1   g617(.A(KEYINPUT109), .B(G137), .Z(new_n804));
  XNOR2_X1  g618(.A(new_n803), .B(new_n804), .ZN(G39));
  AND2_X1   g619(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n806));
  NOR2_X1   g620(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n799), .B(new_n377), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n808), .B1(new_n800), .B2(new_n807), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n591), .A2(new_n593), .B1(G472), .B2(new_n604), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n810), .A2(new_n526), .A3(new_n720), .A4(new_n801), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(new_n395), .ZN(G42));
  NOR3_X1   g627(.A1(new_n526), .A2(new_n716), .A3(new_n378), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n728), .A2(new_n363), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n815), .A2(KEYINPUT49), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(KEYINPUT49), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n814), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  OR4_X1    g632(.A1(new_n712), .A2(new_n714), .A3(new_n783), .A4(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n790), .A2(new_n303), .A3(new_n754), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n315), .B1(KEYINPUT113), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n730), .A2(new_n822), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n820), .A2(new_n714), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n821), .A2(KEYINPUT113), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n824), .B(new_n825), .Z(new_n826));
  INV_X1    g640(.A(KEYINPUT51), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n809), .B1(new_n379), .B2(new_n815), .ZN(new_n828));
  INV_X1    g642(.A(new_n820), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(new_n829), .A3(new_n801), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n801), .A2(new_n730), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n790), .A2(new_n303), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n761), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n525), .A2(new_n303), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n712), .A2(new_n831), .A3(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n739), .A3(new_n785), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n830), .A2(new_n835), .A3(new_n838), .ZN(new_n839));
  OR3_X1    g653(.A1(new_n826), .A2(new_n827), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n827), .B1(new_n826), .B2(new_n839), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n834), .A2(new_n842), .A3(KEYINPUT48), .A4(new_n606), .ZN(new_n843));
  XNOR2_X1  g657(.A(KEYINPUT114), .B(KEYINPUT48), .ZN(new_n844));
  INV_X1    g658(.A(new_n606), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n844), .B1(new_n833), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n829), .A2(new_n745), .ZN(new_n847));
  INV_X1    g661(.A(new_n645), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n302), .B1(new_n837), .B2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n843), .A2(new_n846), .A3(new_n847), .A4(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT115), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n840), .B(new_n841), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n735), .A2(new_n758), .A3(new_n732), .A4(new_n743), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n713), .A2(new_n771), .A3(new_n315), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n810), .A2(new_n526), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n661), .A2(new_n663), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n801), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT111), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n862), .B1(new_n740), .B2(new_n741), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT111), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n863), .A2(new_n690), .A3(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n446), .A2(new_n447), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n865), .A2(new_n677), .A3(new_n701), .A4(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n861), .A2(new_n868), .ZN(new_n869));
  AOI22_X1  g683(.A1(new_n859), .A2(new_n779), .B1(new_n869), .B2(new_n687), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n720), .A2(new_n761), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT112), .B1(new_n871), .B2(new_n858), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT112), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n772), .A2(new_n873), .A3(new_n720), .A4(new_n761), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n863), .A2(new_n864), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n739), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n316), .B1(new_n878), .B2(new_n645), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n616), .A2(new_n620), .A3(new_n879), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n880), .A2(new_n682), .A3(new_n607), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n857), .A2(new_n876), .A3(new_n777), .A4(new_n881), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n693), .A2(new_n762), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n715), .A2(new_n691), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n677), .A2(new_n689), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n712), .A2(new_n771), .A3(new_n884), .A4(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n725), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT52), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n693), .A2(new_n762), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n889), .B1(new_n723), .B2(new_n724), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT52), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n890), .A2(new_n891), .A3(new_n886), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n855), .B1(new_n882), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n891), .B1(new_n890), .B2(new_n886), .ZN(new_n895));
  AND4_X1   g709(.A1(new_n891), .A2(new_n725), .A3(new_n883), .A4(new_n886), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n777), .A2(new_n875), .A3(new_n870), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n880), .A2(new_n682), .A3(new_n607), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n898), .A2(new_n856), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n889), .A2(KEYINPUT52), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n855), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n897), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n894), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT54), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n897), .A2(new_n900), .A3(KEYINPUT53), .A4(new_n901), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n906), .A2(new_n894), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n854), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(G952), .A2(G953), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n819), .B1(new_n910), .B2(new_n911), .ZN(G75));
  NAND2_X1  g726(.A1(new_n906), .A2(new_n894), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n913), .A2(G210), .A3(G902), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n914), .A2(KEYINPUT56), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n246), .A2(new_n276), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(new_n274), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT55), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n306), .A2(G952), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  XNOR2_X1  g735(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n921), .B1(new_n914), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n919), .A2(new_n924), .ZN(G51));
  NAND2_X1  g739(.A1(new_n901), .A2(KEYINPUT53), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n882), .A2(new_n893), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(KEYINPUT53), .B1(new_n897), .B2(new_n900), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n929), .A2(new_n308), .A3(new_n794), .ZN(new_n930));
  INV_X1    g744(.A(new_n361), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT54), .B1(new_n927), .B2(new_n928), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n908), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n371), .B(KEYINPUT57), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT117), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n930), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n934), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n938), .B1(new_n932), .B2(new_n908), .ZN(new_n939));
  OAI21_X1  g753(.A(KEYINPUT117), .B1(new_n939), .B2(new_n931), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n920), .B1(new_n937), .B2(new_n940), .ZN(G54));
  NAND4_X1  g755(.A1(new_n913), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n942));
  INV_X1    g756(.A(new_n439), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n944), .A2(new_n945), .A3(new_n920), .ZN(G60));
  NAND2_X1  g760(.A1(new_n636), .A2(new_n638), .ZN(new_n947));
  XOR2_X1   g761(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(new_n621), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n933), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n947), .B1(new_n909), .B2(new_n949), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n950), .A2(new_n951), .A3(new_n920), .ZN(G63));
  XNOR2_X1  g766(.A(KEYINPUT119), .B(KEYINPUT60), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n515), .A2(new_n308), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n514), .B1(new_n929), .B2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n674), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n913), .A2(new_n958), .A3(new_n955), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n957), .A2(new_n921), .A3(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT61), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(G66));
  OAI21_X1  g776(.A(G953), .B1(new_n312), .B2(new_n271), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n856), .A2(new_n899), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n963), .B1(new_n964), .B2(new_n307), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n916), .B1(G898), .B2(new_n306), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(G69));
  NAND2_X1  g781(.A1(new_n563), .A2(new_n542), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(new_n433), .Z(new_n969));
  XNOR2_X1  g783(.A(KEYINPUT120), .B(KEYINPUT121), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n969), .B(new_n970), .Z(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT122), .Z(new_n972));
  INV_X1    g786(.A(KEYINPUT62), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n890), .A2(new_n973), .A3(new_n718), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT123), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n812), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n803), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n973), .B1(new_n890), .B2(new_n718), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n703), .A2(new_n801), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(new_n645), .B2(new_n878), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n980), .B1(new_n606), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n976), .A2(new_n979), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n972), .B1(new_n984), .B2(new_n306), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n800), .A2(new_n606), .A3(new_n702), .A4(new_n884), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n777), .A2(new_n780), .A3(new_n986), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n979), .A2(KEYINPUT124), .A3(new_n890), .A4(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT124), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n987), .A2(new_n890), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n989), .B1(new_n990), .B2(new_n978), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n988), .A2(new_n991), .A3(new_n306), .ZN(new_n992));
  INV_X1    g806(.A(new_n971), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n993), .B1(G900), .B2(new_n307), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n985), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n972), .A2(KEYINPUT125), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n306), .B1(G227), .B2(G900), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n995), .B(new_n998), .ZN(G72));
  XNOR2_X1  g813(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n706), .A2(new_n308), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1000), .B(new_n1001), .Z(new_n1002));
  INV_X1    g816(.A(new_n964), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1002), .B1(new_n984), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(new_n600), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1004), .A2(new_n560), .A3(new_n1005), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n1005), .A2(new_n560), .ZN(new_n1007));
  AND3_X1   g821(.A1(new_n988), .A2(new_n991), .A3(new_n964), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1002), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(new_n601), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1009), .B1(new_n1011), .B2(new_n707), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n920), .B1(new_n904), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1006), .A2(new_n1010), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(KEYINPUT127), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT127), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n1006), .A2(new_n1010), .A3(new_n1016), .A4(new_n1013), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1015), .A2(new_n1017), .ZN(G57));
endmodule


