

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738;

  NOR2_X1 U380 ( .A1(n684), .A2(n581), .ZN(n573) );
  AND2_X1 U381 ( .A1(n713), .A2(n614), .ZN(n690) );
  INV_X1 U382 ( .A(G953), .ZN(n727) );
  NOR2_X1 U383 ( .A1(n581), .A2(n580), .ZN(n640) );
  XNOR2_X2 U384 ( .A(G128), .B(KEYINPUT65), .ZN(n439) );
  NOR2_X1 U385 ( .A1(n529), .A2(KEYINPUT71), .ZN(n528) );
  INV_X1 U386 ( .A(n605), .ZN(n668) );
  NOR2_X1 U387 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U388 ( .A1(n735), .A2(n632), .ZN(n527) );
  XNOR2_X1 U389 ( .A(n570), .B(n469), .ZN(n605) );
  XNOR2_X1 U390 ( .A(n480), .B(n479), .ZN(n720) );
  XNOR2_X1 U391 ( .A(n443), .B(n442), .ZN(n477) );
  XOR2_X1 U392 ( .A(KEYINPUT3), .B(G116), .Z(n443) );
  XNOR2_X1 U393 ( .A(G119), .B(G101), .ZN(n442) );
  XNOR2_X2 U394 ( .A(n428), .B(n361), .ZN(n569) );
  XNOR2_X1 U395 ( .A(n371), .B(KEYINPUT115), .ZN(n658) );
  OR2_X1 U396 ( .A1(n656), .A2(n657), .ZN(n371) );
  XNOR2_X1 U397 ( .A(n444), .B(n458), .ZN(n724) );
  XNOR2_X1 U398 ( .A(n384), .B(n450), .ZN(n622) );
  XNOR2_X1 U399 ( .A(n444), .B(n477), .ZN(n384) );
  XNOR2_X1 U400 ( .A(G137), .B(G113), .ZN(n448) );
  XNOR2_X1 U401 ( .A(n720), .B(n481), .ZN(n700) );
  XNOR2_X1 U402 ( .A(n405), .B(n404), .ZN(n476) );
  XNOR2_X1 U403 ( .A(n474), .B(n473), .ZN(n404) );
  NOR2_X1 U404 ( .A1(n634), .A2(n639), .ZN(n538) );
  NOR2_X1 U405 ( .A1(G953), .A2(G237), .ZN(n507) );
  NAND2_X1 U406 ( .A1(G237), .A2(G234), .ZN(n487) );
  XNOR2_X1 U407 ( .A(G131), .B(G134), .ZN(n440) );
  XNOR2_X1 U408 ( .A(n452), .B(n451), .ZN(n495) );
  INV_X1 U409 ( .A(KEYINPUT8), .ZN(n451) );
  XNOR2_X1 U410 ( .A(G110), .B(G104), .ZN(n434) );
  XOR2_X1 U411 ( .A(G101), .B(G107), .Z(n435) );
  XNOR2_X1 U412 ( .A(KEYINPUT38), .B(KEYINPUT73), .ZN(n368) );
  OR2_X1 U413 ( .A1(G902), .A2(G237), .ZN(n484) );
  XNOR2_X1 U414 ( .A(n383), .B(n382), .ZN(n540) );
  INV_X1 U415 ( .A(G472), .ZN(n382) );
  OR2_X1 U416 ( .A1(n622), .A2(G902), .ZN(n383) );
  AND2_X1 U417 ( .A1(n594), .A2(n592), .ZN(n393) );
  INV_X1 U418 ( .A(n540), .ZN(n673) );
  XOR2_X1 U419 ( .A(KEYINPUT6), .B(n540), .Z(n595) );
  NOR2_X1 U420 ( .A1(G902), .A2(n466), .ZN(n467) );
  XOR2_X1 U421 ( .A(G104), .B(G113), .Z(n511) );
  XOR2_X1 U422 ( .A(G137), .B(G140), .Z(n458) );
  XNOR2_X1 U423 ( .A(G116), .B(KEYINPUT9), .ZN(n498) );
  INV_X1 U424 ( .A(G143), .ZN(n429) );
  NAND2_X1 U425 ( .A1(n432), .A2(n431), .ZN(n430) );
  INV_X1 U426 ( .A(n613), .ZN(n431) );
  XNOR2_X1 U427 ( .A(n421), .B(n419), .ZN(n536) );
  XNOR2_X1 U428 ( .A(n420), .B(KEYINPUT98), .ZN(n419) );
  OR2_X1 U429 ( .A1(n705), .A2(G902), .ZN(n421) );
  INV_X1 U430 ( .A(G478), .ZN(n420) );
  BUF_X1 U431 ( .A(n668), .Z(n378) );
  BUF_X1 U432 ( .A(n673), .Z(n367) );
  OR2_X1 U433 ( .A1(n711), .A2(G902), .ZN(n428) );
  XNOR2_X1 U434 ( .A(KEYINPUT67), .B(KEYINPUT22), .ZN(n525) );
  NAND2_X1 U435 ( .A1(n541), .A2(n524), .ZN(n526) );
  AND2_X1 U436 ( .A1(n523), .A2(n592), .ZN(n524) );
  XNOR2_X1 U437 ( .A(n622), .B(n621), .ZN(n418) );
  XNOR2_X1 U438 ( .A(n415), .B(n413), .ZN(n711) );
  XNOR2_X1 U439 ( .A(n455), .B(n414), .ZN(n413) );
  XNOR2_X1 U440 ( .A(n725), .B(n433), .ZN(n415) );
  XNOR2_X1 U441 ( .A(n458), .B(n459), .ZN(n414) );
  NAND2_X1 U442 ( .A1(n710), .A2(G217), .ZN(n388) );
  XNOR2_X1 U443 ( .A(n700), .B(n698), .ZN(n408) );
  XOR2_X1 U444 ( .A(KEYINPUT86), .B(n616), .Z(n712) );
  XNOR2_X1 U445 ( .A(n650), .B(n598), .ZN(n599) );
  INV_X1 U446 ( .A(KEYINPUT116), .ZN(n373) );
  XOR2_X1 U447 ( .A(G146), .B(KEYINPUT5), .Z(n446) );
  XNOR2_X1 U448 ( .A(G143), .B(G131), .ZN(n504) );
  XOR2_X1 U449 ( .A(KEYINPUT96), .B(G122), .Z(n505) );
  XOR2_X1 U450 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n509) );
  XNOR2_X1 U451 ( .A(n456), .B(G146), .ZN(n474) );
  INV_X1 U452 ( .A(G125), .ZN(n456) );
  XNOR2_X1 U453 ( .A(KEYINPUT87), .B(KEYINPUT85), .ZN(n473) );
  XNOR2_X1 U454 ( .A(n363), .B(n358), .ZN(n405) );
  NAND2_X1 U455 ( .A1(n369), .A2(n713), .ZN(n432) );
  XNOR2_X1 U456 ( .A(n390), .B(KEYINPUT81), .ZN(n369) );
  INV_X1 U457 ( .A(n576), .ZN(n561) );
  XNOR2_X1 U458 ( .A(G902), .B(KEYINPUT15), .ZN(n613) );
  OR2_X1 U459 ( .A1(n359), .A2(n399), .ZN(n398) );
  XNOR2_X1 U460 ( .A(G110), .B(G119), .ZN(n459) );
  XNOR2_X1 U461 ( .A(n457), .B(KEYINPUT68), .ZN(n725) );
  XNOR2_X1 U462 ( .A(n474), .B(KEYINPUT10), .ZN(n457) );
  XNOR2_X1 U463 ( .A(n724), .B(n441), .ZN(n466) );
  XNOR2_X1 U464 ( .A(n680), .B(n374), .ZN(n681) );
  XNOR2_X1 U465 ( .A(KEYINPUT118), .B(KEYINPUT52), .ZN(n374) );
  NOR2_X1 U466 ( .A1(n655), .A2(n656), .ZN(n568) );
  NOR2_X1 U467 ( .A1(n642), .A2(n422), .ZN(n604) );
  AND2_X1 U468 ( .A1(n661), .A2(n541), .ZN(n493) );
  XNOR2_X1 U469 ( .A(n380), .B(KEYINPUT93), .ZN(n675) );
  OR2_X1 U470 ( .A1(n539), .A2(n540), .ZN(n380) );
  XNOR2_X1 U471 ( .A(n392), .B(n391), .ZN(n571) );
  INV_X1 U472 ( .A(KEYINPUT28), .ZN(n391) );
  NAND2_X1 U473 ( .A1(n367), .A2(n393), .ZN(n392) );
  XNOR2_X1 U474 ( .A(n426), .B(n427), .ZN(n556) );
  INV_X1 U475 ( .A(KEYINPUT90), .ZN(n427) );
  AND2_X1 U476 ( .A1(n569), .A2(n592), .ZN(n370) );
  AND2_X2 U477 ( .A1(n397), .A2(n394), .ZN(n541) );
  NAND2_X1 U478 ( .A1(n396), .A2(n395), .ZN(n394) );
  AND2_X1 U479 ( .A1(n400), .A2(n398), .ZN(n397) );
  AND2_X1 U480 ( .A1(n359), .A2(n399), .ZN(n395) );
  XOR2_X1 U481 ( .A(KEYINPUT16), .B(n477), .Z(n480) );
  XNOR2_X1 U482 ( .A(n503), .B(n502), .ZN(n705) );
  XNOR2_X1 U483 ( .A(n566), .B(n565), .ZN(n737) );
  NOR2_X1 U484 ( .A1(n642), .A2(n610), .ZN(n566) );
  XNOR2_X1 U485 ( .A(n402), .B(n365), .ZN(n735) );
  XNOR2_X1 U486 ( .A(n537), .B(KEYINPUT99), .ZN(n639) );
  NOR2_X1 U487 ( .A1(n378), .A2(n367), .ZN(n401) );
  NAND2_X1 U488 ( .A1(n417), .A2(n712), .ZN(n416) );
  XNOR2_X1 U489 ( .A(n620), .B(n418), .ZN(n417) );
  NAND2_X1 U490 ( .A1(n386), .A2(n712), .ZN(n385) );
  XNOR2_X1 U491 ( .A(n388), .B(n387), .ZN(n386) );
  INV_X1 U492 ( .A(n711), .ZN(n387) );
  XNOR2_X1 U493 ( .A(KEYINPUT123), .B(KEYINPUT60), .ZN(n410) );
  NAND2_X1 U494 ( .A1(n412), .A2(n712), .ZN(n411) );
  XNOR2_X1 U495 ( .A(n703), .B(n704), .ZN(n412) );
  NAND2_X1 U496 ( .A1(n407), .A2(n712), .ZN(n406) );
  XNOR2_X1 U497 ( .A(n699), .B(n408), .ZN(n407) );
  XNOR2_X1 U498 ( .A(n696), .B(n375), .ZN(G75) );
  XNOR2_X1 U499 ( .A(n697), .B(n376), .ZN(n375) );
  INV_X1 U500 ( .A(KEYINPUT121), .ZN(n376) );
  XOR2_X1 U501 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n358) );
  OR2_X1 U502 ( .A1(n560), .A2(n491), .ZN(n359) );
  AND2_X1 U503 ( .A1(n521), .A2(n378), .ZN(n360) );
  XOR2_X1 U504 ( .A(n463), .B(n462), .Z(n361) );
  AND2_X1 U505 ( .A1(n360), .A2(n663), .ZN(n362) );
  AND2_X1 U506 ( .A1(G224), .A2(n727), .ZN(n363) );
  AND2_X1 U507 ( .A1(n612), .A2(KEYINPUT2), .ZN(n364) );
  XOR2_X1 U508 ( .A(KEYINPUT66), .B(KEYINPUT32), .Z(n365) );
  XOR2_X1 U509 ( .A(n552), .B(KEYINPUT45), .Z(n366) );
  NOR2_X1 U510 ( .A1(n595), .A2(n593), .ZN(n423) );
  INV_X1 U511 ( .A(n541), .ZN(n544) );
  INV_X1 U512 ( .A(n575), .ZN(n381) );
  NAND2_X1 U513 ( .A1(n555), .A2(n556), .ZN(n575) );
  XNOR2_X1 U514 ( .A(n557), .B(n368), .ZN(n653) );
  NAND2_X1 U515 ( .A1(n570), .A2(n370), .ZN(n426) );
  NAND2_X1 U516 ( .A1(n372), .A2(n685), .ZN(n662) );
  XNOR2_X1 U517 ( .A(n660), .B(n373), .ZN(n372) );
  NOR2_X4 U518 ( .A1(n377), .A2(n430), .ZN(n710) );
  NOR2_X2 U519 ( .A1(n690), .A2(KEYINPUT2), .ZN(n377) );
  XNOR2_X1 U520 ( .A(n379), .B(KEYINPUT95), .ZN(n547) );
  NAND2_X1 U521 ( .A1(n646), .A2(n627), .ZN(n379) );
  NAND2_X1 U522 ( .A1(n381), .A2(n562), .ZN(n563) );
  XNOR2_X2 U523 ( .A(n475), .B(n440), .ZN(n444) );
  XNOR2_X1 U524 ( .A(n385), .B(KEYINPUT125), .ZN(G66) );
  XNOR2_X2 U525 ( .A(n520), .B(n519), .ZN(n734) );
  XNOR2_X1 U526 ( .A(n411), .B(n410), .ZN(G60) );
  XNOR2_X1 U527 ( .A(n416), .B(n623), .ZN(G57) );
  XNOR2_X1 U528 ( .A(n603), .B(KEYINPUT48), .ZN(n389) );
  AND2_X1 U529 ( .A1(n389), .A2(n612), .ZN(n614) );
  NAND2_X1 U530 ( .A1(n389), .A2(n364), .ZN(n390) );
  INV_X1 U531 ( .A(n580), .ZN(n396) );
  INV_X1 U532 ( .A(KEYINPUT0), .ZN(n399) );
  NAND2_X1 U533 ( .A1(n580), .A2(KEYINPUT0), .ZN(n400) );
  XNOR2_X2 U534 ( .A(n485), .B(n486), .ZN(n580) );
  NAND2_X1 U535 ( .A1(n362), .A2(n530), .ZN(n402) );
  AND2_X1 U536 ( .A1(n530), .A2(n663), .ZN(n403) );
  AND2_X1 U537 ( .A1(n403), .A2(n401), .ZN(n632) );
  XNOR2_X1 U538 ( .A(n406), .B(n701), .ZN(G51) );
  INV_X1 U539 ( .A(n432), .ZN(n692) );
  XNOR2_X2 U540 ( .A(n409), .B(n366), .ZN(n713) );
  NAND2_X1 U541 ( .A1(n550), .A2(n551), .ZN(n409) );
  AND2_X1 U542 ( .A1(n557), .A2(n604), .ZN(n596) );
  NAND2_X1 U543 ( .A1(n423), .A2(n594), .ZN(n422) );
  XNOR2_X1 U544 ( .A(n425), .B(n424), .ZN(n617) );
  XNOR2_X1 U545 ( .A(n615), .B(KEYINPUT57), .ZN(n424) );
  NAND2_X1 U546 ( .A1(n710), .A2(G469), .ZN(n425) );
  XNOR2_X2 U547 ( .A(n467), .B(n468), .ZN(n570) );
  XNOR2_X2 U548 ( .A(n501), .B(KEYINPUT4), .ZN(n475) );
  XNOR2_X2 U549 ( .A(n439), .B(n429), .ZN(n501) );
  XNOR2_X1 U550 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U551 ( .A(n454), .B(n453), .Z(n433) );
  INV_X1 U552 ( .A(KEYINPUT83), .ZN(n598) );
  NAND2_X1 U553 ( .A1(n727), .A2(G234), .ZN(n452) );
  XNOR2_X1 U554 ( .A(n470), .B(KEYINPUT101), .ZN(n471) );
  XNOR2_X1 U555 ( .A(n472), .B(n471), .ZN(n661) );
  AND2_X1 U556 ( .A1(n653), .A2(n561), .ZN(n562) );
  INV_X1 U557 ( .A(KEYINPUT122), .ZN(n619) );
  XNOR2_X1 U558 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U559 ( .A(G146), .B(n436), .Z(n438) );
  NAND2_X1 U560 ( .A1(G227), .A2(n727), .ZN(n437) );
  XNOR2_X1 U561 ( .A(n438), .B(n437), .ZN(n441) );
  XNOR2_X1 U562 ( .A(n466), .B(KEYINPUT58), .ZN(n615) );
  NAND2_X1 U563 ( .A1(G210), .A2(n507), .ZN(n445) );
  XNOR2_X1 U564 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U565 ( .A(n447), .B(KEYINPUT91), .Z(n449) );
  XNOR2_X1 U566 ( .A(n449), .B(n448), .ZN(n450) );
  NAND2_X1 U567 ( .A1(G221), .A2(n495), .ZN(n455) );
  XOR2_X1 U568 ( .A(KEYINPUT24), .B(KEYINPUT88), .Z(n454) );
  XNOR2_X1 U569 ( .A(G128), .B(KEYINPUT23), .ZN(n453) );
  XOR2_X1 U570 ( .A(KEYINPUT20), .B(KEYINPUT89), .Z(n461) );
  NAND2_X1 U571 ( .A1(G234), .A2(n613), .ZN(n460) );
  XNOR2_X1 U572 ( .A(n461), .B(n460), .ZN(n464) );
  AND2_X1 U573 ( .A1(G217), .A2(n464), .ZN(n463) );
  XNOR2_X1 U574 ( .A(KEYINPUT25), .B(KEYINPUT75), .ZN(n462) );
  NAND2_X1 U575 ( .A1(n464), .A2(G221), .ZN(n465) );
  XNOR2_X1 U576 ( .A(n465), .B(KEYINPUT21), .ZN(n664) );
  INV_X1 U577 ( .A(n664), .ZN(n592) );
  AND2_X1 U578 ( .A1(n569), .A2(n592), .ZN(n667) );
  XNOR2_X1 U579 ( .A(KEYINPUT69), .B(G469), .ZN(n468) );
  INV_X1 U580 ( .A(KEYINPUT1), .ZN(n469) );
  NAND2_X1 U581 ( .A1(n667), .A2(n668), .ZN(n539) );
  NOR2_X1 U582 ( .A1(n595), .A2(n539), .ZN(n472) );
  XNOR2_X1 U583 ( .A(KEYINPUT33), .B(KEYINPUT70), .ZN(n470) );
  XOR2_X1 U584 ( .A(KEYINPUT74), .B(KEYINPUT19), .Z(n486) );
  XNOR2_X1 U585 ( .A(n475), .B(n476), .ZN(n481) );
  XOR2_X1 U586 ( .A(G107), .B(G122), .Z(n494) );
  XNOR2_X1 U587 ( .A(G110), .B(n494), .ZN(n478) );
  XNOR2_X1 U588 ( .A(n478), .B(n511), .ZN(n479) );
  NAND2_X1 U589 ( .A1(n700), .A2(n613), .ZN(n483) );
  AND2_X1 U590 ( .A1(G210), .A2(n484), .ZN(n482) );
  XNOR2_X2 U591 ( .A(n483), .B(n482), .ZN(n557) );
  NAND2_X1 U592 ( .A1(G214), .A2(n484), .ZN(n652) );
  NAND2_X1 U593 ( .A1(n557), .A2(n652), .ZN(n485) );
  XNOR2_X1 U594 ( .A(n487), .B(KEYINPUT14), .ZN(n488) );
  XNOR2_X1 U595 ( .A(KEYINPUT72), .B(n488), .ZN(n489) );
  NAND2_X1 U596 ( .A1(G952), .A2(n489), .ZN(n682) );
  NOR2_X1 U597 ( .A1(G953), .A2(n682), .ZN(n560) );
  AND2_X1 U598 ( .A1(n489), .A2(G953), .ZN(n490) );
  NAND2_X1 U599 ( .A1(G902), .A2(n490), .ZN(n558) );
  NOR2_X1 U600 ( .A1(G898), .A2(n558), .ZN(n491) );
  XNOR2_X1 U601 ( .A(KEYINPUT76), .B(KEYINPUT34), .ZN(n492) );
  XNOR2_X1 U602 ( .A(n493), .B(n492), .ZN(n518) );
  XOR2_X1 U603 ( .A(G134), .B(n494), .Z(n497) );
  NAND2_X1 U604 ( .A1(G217), .A2(n495), .ZN(n496) );
  XNOR2_X1 U605 ( .A(n497), .B(n496), .ZN(n503) );
  XOR2_X1 U606 ( .A(KEYINPUT97), .B(KEYINPUT7), .Z(n499) );
  XNOR2_X1 U607 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U608 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U609 ( .A(n725), .B(n506), .ZN(n515) );
  NAND2_X1 U610 ( .A1(n507), .A2(G214), .ZN(n508) );
  XNOR2_X1 U611 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U612 ( .A(G140), .B(n510), .ZN(n513) );
  INV_X1 U613 ( .A(n511), .ZN(n512) );
  XNOR2_X1 U614 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U615 ( .A(n515), .B(n514), .ZN(n702) );
  NOR2_X1 U616 ( .A1(G902), .A2(n702), .ZN(n517) );
  XNOR2_X1 U617 ( .A(KEYINPUT13), .B(G475), .ZN(n516) );
  XNOR2_X1 U618 ( .A(n517), .B(n516), .ZN(n535) );
  INV_X1 U619 ( .A(n535), .ZN(n522) );
  NOR2_X1 U620 ( .A1(n536), .A2(n522), .ZN(n578) );
  NAND2_X1 U621 ( .A1(n518), .A2(n578), .ZN(n520) );
  INV_X1 U622 ( .A(KEYINPUT35), .ZN(n519) );
  INV_X1 U623 ( .A(n595), .ZN(n532) );
  XNOR2_X1 U624 ( .A(KEYINPUT77), .B(n532), .ZN(n521) );
  INV_X1 U625 ( .A(n569), .ZN(n663) );
  NAND2_X1 U626 ( .A1(n522), .A2(n536), .ZN(n655) );
  INV_X1 U627 ( .A(n655), .ZN(n523) );
  XNOR2_X1 U628 ( .A(n526), .B(n525), .ZN(n530) );
  NAND2_X1 U629 ( .A1(n734), .A2(n527), .ZN(n529) );
  XNOR2_X1 U630 ( .A(n528), .B(KEYINPUT44), .ZN(n551) );
  NAND2_X1 U631 ( .A1(n529), .A2(KEYINPUT71), .ZN(n534) );
  NAND2_X1 U632 ( .A1(n605), .A2(n530), .ZN(n531) );
  NOR2_X1 U633 ( .A1(n532), .A2(n531), .ZN(n533) );
  NAND2_X1 U634 ( .A1(n533), .A2(n569), .ZN(n624) );
  NAND2_X1 U635 ( .A1(n534), .A2(n624), .ZN(n549) );
  NOR2_X1 U636 ( .A1(n535), .A2(n536), .ZN(n634) );
  NAND2_X1 U637 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U638 ( .A(n538), .B(KEYINPUT100), .ZN(n657) );
  XOR2_X1 U639 ( .A(KEYINPUT94), .B(KEYINPUT31), .Z(n543) );
  NAND2_X1 U640 ( .A1(n675), .A2(n541), .ZN(n542) );
  XNOR2_X1 U641 ( .A(n543), .B(n542), .ZN(n646) );
  NOR2_X1 U642 ( .A1(n544), .A2(n367), .ZN(n545) );
  NAND2_X1 U643 ( .A1(n556), .A2(n545), .ZN(n546) );
  XNOR2_X1 U644 ( .A(KEYINPUT92), .B(n546), .ZN(n627) );
  NOR2_X1 U645 ( .A1(n657), .A2(n547), .ZN(n548) );
  NOR2_X1 U646 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U647 ( .A(KEYINPUT80), .B(KEYINPUT64), .Z(n552) );
  INV_X1 U648 ( .A(n639), .ZN(n642) );
  XOR2_X1 U649 ( .A(KEYINPUT84), .B(KEYINPUT39), .Z(n564) );
  NAND2_X1 U650 ( .A1(n652), .A2(n673), .ZN(n554) );
  XNOR2_X1 U651 ( .A(KEYINPUT30), .B(KEYINPUT103), .ZN(n553) );
  XNOR2_X1 U652 ( .A(n554), .B(n553), .ZN(n555) );
  NOR2_X1 U653 ( .A1(G900), .A2(n558), .ZN(n559) );
  NOR2_X1 U654 ( .A1(n560), .A2(n559), .ZN(n576) );
  XNOR2_X1 U655 ( .A(n564), .B(n563), .ZN(n610) );
  INV_X1 U656 ( .A(KEYINPUT40), .ZN(n565) );
  NAND2_X1 U657 ( .A1(n653), .A2(n652), .ZN(n656) );
  XNOR2_X1 U658 ( .A(KEYINPUT41), .B(KEYINPUT104), .ZN(n567) );
  XNOR2_X1 U659 ( .A(n568), .B(n567), .ZN(n684) );
  NOR2_X1 U660 ( .A1(n576), .A2(n569), .ZN(n594) );
  NAND2_X1 U661 ( .A1(n571), .A2(n570), .ZN(n581) );
  XNOR2_X1 U662 ( .A(KEYINPUT42), .B(KEYINPUT105), .ZN(n572) );
  XNOR2_X1 U663 ( .A(n573), .B(n572), .ZN(n738) );
  NAND2_X1 U664 ( .A1(n737), .A2(n738), .ZN(n574) );
  XNOR2_X1 U665 ( .A(KEYINPUT46), .B(n574), .ZN(n602) );
  INV_X1 U666 ( .A(n557), .ZN(n607) );
  NOR2_X1 U667 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U668 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U669 ( .A1(n607), .A2(n579), .ZN(n638) );
  INV_X1 U670 ( .A(n657), .ZN(n587) );
  OR2_X1 U671 ( .A1(n587), .A2(KEYINPUT79), .ZN(n582) );
  NAND2_X1 U672 ( .A1(n640), .A2(n582), .ZN(n583) );
  NAND2_X1 U673 ( .A1(n583), .A2(KEYINPUT47), .ZN(n585) );
  NAND2_X1 U674 ( .A1(n587), .A2(KEYINPUT79), .ZN(n584) );
  NAND2_X1 U675 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U676 ( .A1(n638), .A2(n586), .ZN(n591) );
  AND2_X1 U677 ( .A1(n587), .A2(n640), .ZN(n588) );
  NOR2_X1 U678 ( .A1(n588), .A2(KEYINPUT79), .ZN(n589) );
  OR2_X1 U679 ( .A1(KEYINPUT47), .A2(n589), .ZN(n590) );
  AND2_X1 U680 ( .A1(n591), .A2(n590), .ZN(n600) );
  NAND2_X1 U681 ( .A1(n592), .A2(n652), .ZN(n593) );
  XNOR2_X1 U682 ( .A(n596), .B(KEYINPUT36), .ZN(n597) );
  NAND2_X1 U683 ( .A1(n597), .A2(n378), .ZN(n650) );
  NAND2_X1 U684 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U685 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U686 ( .A(n606), .B(KEYINPUT43), .ZN(n608) );
  NAND2_X1 U687 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U688 ( .A(KEYINPUT102), .B(n609), .ZN(n736) );
  INV_X1 U689 ( .A(n634), .ZN(n645) );
  NOR2_X1 U690 ( .A1(n610), .A2(n645), .ZN(n651) );
  INV_X1 U691 ( .A(n651), .ZN(n611) );
  AND2_X1 U692 ( .A1(n736), .A2(n611), .ZN(n612) );
  NOR2_X1 U693 ( .A1(G952), .A2(n727), .ZN(n616) );
  NAND2_X1 U694 ( .A1(n617), .A2(n712), .ZN(n618) );
  XNOR2_X1 U695 ( .A(n619), .B(n618), .ZN(G54) );
  XOR2_X1 U696 ( .A(KEYINPUT62), .B(KEYINPUT106), .Z(n621) );
  NAND2_X1 U697 ( .A1(n710), .A2(G472), .ZN(n620) );
  XOR2_X1 U698 ( .A(KEYINPUT63), .B(KEYINPUT107), .Z(n623) );
  XNOR2_X1 U699 ( .A(G101), .B(n624), .ZN(G3) );
  NOR2_X1 U700 ( .A1(n627), .A2(n642), .ZN(n625) );
  XOR2_X1 U701 ( .A(KEYINPUT108), .B(n625), .Z(n626) );
  XNOR2_X1 U702 ( .A(G104), .B(n626), .ZN(G6) );
  NOR2_X1 U703 ( .A1(n645), .A2(n627), .ZN(n631) );
  XOR2_X1 U704 ( .A(KEYINPUT109), .B(KEYINPUT26), .Z(n629) );
  XNOR2_X1 U705 ( .A(G107), .B(KEYINPUT27), .ZN(n628) );
  XNOR2_X1 U706 ( .A(n629), .B(n628), .ZN(n630) );
  XNOR2_X1 U707 ( .A(n631), .B(n630), .ZN(G9) );
  XOR2_X1 U708 ( .A(G110), .B(n632), .Z(n633) );
  XNOR2_X1 U709 ( .A(KEYINPUT110), .B(n633), .ZN(G12) );
  XOR2_X1 U710 ( .A(KEYINPUT111), .B(KEYINPUT29), .Z(n636) );
  NAND2_X1 U711 ( .A1(n640), .A2(n634), .ZN(n635) );
  XNOR2_X1 U712 ( .A(n636), .B(n635), .ZN(n637) );
  XOR2_X1 U713 ( .A(G128), .B(n637), .Z(G30) );
  XOR2_X1 U714 ( .A(G143), .B(n638), .Z(G45) );
  NAND2_X1 U715 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U716 ( .A(n641), .B(G146), .ZN(G48) );
  NOR2_X1 U717 ( .A1(n646), .A2(n642), .ZN(n643) );
  XOR2_X1 U718 ( .A(KEYINPUT112), .B(n643), .Z(n644) );
  XNOR2_X1 U719 ( .A(G113), .B(n644), .ZN(G15) );
  NOR2_X1 U720 ( .A1(n646), .A2(n645), .ZN(n648) );
  XNOR2_X1 U721 ( .A(G116), .B(KEYINPUT113), .ZN(n647) );
  XNOR2_X1 U722 ( .A(n648), .B(n647), .ZN(G18) );
  XOR2_X1 U723 ( .A(G125), .B(KEYINPUT37), .Z(n649) );
  XNOR2_X1 U724 ( .A(n650), .B(n649), .ZN(G27) );
  XOR2_X1 U725 ( .A(G134), .B(n651), .Z(G36) );
  XOR2_X1 U726 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n697) );
  NOR2_X1 U727 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U728 ( .A1(n655), .A2(n654), .ZN(n659) );
  NOR2_X1 U729 ( .A1(n659), .A2(n658), .ZN(n660) );
  BUF_X1 U730 ( .A(n661), .Z(n685) );
  XNOR2_X1 U731 ( .A(n662), .B(KEYINPUT117), .ZN(n679) );
  XOR2_X1 U732 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n666) );
  NAND2_X1 U733 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U734 ( .A(n666), .B(n665), .ZN(n671) );
  NOR2_X1 U735 ( .A1(n667), .A2(n378), .ZN(n669) );
  XOR2_X1 U736 ( .A(KEYINPUT50), .B(n669), .Z(n670) );
  NAND2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U738 ( .A1(n367), .A2(n672), .ZN(n674) );
  NOR2_X1 U739 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U740 ( .A(KEYINPUT51), .B(n676), .Z(n677) );
  NOR2_X1 U741 ( .A1(n677), .A2(n684), .ZN(n678) );
  NOR2_X1 U742 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U743 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U744 ( .A(n683), .B(KEYINPUT119), .ZN(n688) );
  INV_X1 U745 ( .A(n684), .ZN(n686) );
  NAND2_X1 U746 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U747 ( .A1(n688), .A2(n687), .ZN(n694) );
  XNOR2_X1 U748 ( .A(KEYINPUT2), .B(KEYINPUT78), .ZN(n689) );
  NOR2_X1 U749 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U750 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U751 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U752 ( .A1(n695), .A2(n727), .ZN(n696) );
  NAND2_X1 U753 ( .A1(n710), .A2(G210), .ZN(n699) );
  XOR2_X1 U754 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n698) );
  XOR2_X1 U755 ( .A(KEYINPUT82), .B(KEYINPUT56), .Z(n701) );
  XNOR2_X1 U756 ( .A(n702), .B(KEYINPUT59), .ZN(n704) );
  NAND2_X1 U757 ( .A1(G475), .A2(n710), .ZN(n703) );
  XNOR2_X1 U758 ( .A(n705), .B(KEYINPUT124), .ZN(n707) );
  NAND2_X1 U759 ( .A1(G478), .A2(n710), .ZN(n706) );
  XNOR2_X1 U760 ( .A(n707), .B(n706), .ZN(n709) );
  INV_X1 U761 ( .A(n712), .ZN(n708) );
  NOR2_X1 U762 ( .A1(n709), .A2(n708), .ZN(G63) );
  NAND2_X1 U763 ( .A1(n727), .A2(n713), .ZN(n718) );
  NAND2_X1 U764 ( .A1(G224), .A2(G953), .ZN(n714) );
  XNOR2_X1 U765 ( .A(n714), .B(KEYINPUT61), .ZN(n715) );
  XNOR2_X1 U766 ( .A(KEYINPUT126), .B(n715), .ZN(n716) );
  NAND2_X1 U767 ( .A1(n716), .A2(G898), .ZN(n717) );
  NAND2_X1 U768 ( .A1(n718), .A2(n717), .ZN(n722) );
  NOR2_X1 U769 ( .A1(G898), .A2(n727), .ZN(n719) );
  NOR2_X1 U770 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U771 ( .A(n722), .B(n721), .ZN(n723) );
  XOR2_X1 U772 ( .A(KEYINPUT127), .B(n723), .Z(G69) );
  XOR2_X1 U773 ( .A(n725), .B(n724), .Z(n729) );
  INV_X1 U774 ( .A(n729), .ZN(n726) );
  XNOR2_X1 U775 ( .A(n726), .B(n614), .ZN(n728) );
  NAND2_X1 U776 ( .A1(n728), .A2(n727), .ZN(n733) );
  XNOR2_X1 U777 ( .A(G227), .B(n729), .ZN(n730) );
  NAND2_X1 U778 ( .A1(n730), .A2(G900), .ZN(n731) );
  NAND2_X1 U779 ( .A1(n731), .A2(G953), .ZN(n732) );
  NAND2_X1 U780 ( .A1(n733), .A2(n732), .ZN(G72) );
  XNOR2_X1 U781 ( .A(n734), .B(G122), .ZN(G24) );
  XOR2_X1 U782 ( .A(n735), .B(G119), .Z(G21) );
  XNOR2_X1 U783 ( .A(G140), .B(n736), .ZN(G42) );
  XNOR2_X1 U784 ( .A(G131), .B(n737), .ZN(G33) );
  XNOR2_X1 U785 ( .A(G137), .B(n738), .ZN(G39) );
endmodule

