//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1299, new_n1300, new_n1301, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1378, new_n1379, new_n1380, new_n1381;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n210), .ZN(new_n217));
  INV_X1    g0017(.A(new_n201), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(new_n215), .A2(KEYINPUT0), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n221), .B1(KEYINPUT0), .B2(new_n215), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT64), .Z(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n212), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT1), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n223), .A2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT65), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n202), .A2(G68), .ZN(new_n246));
  INV_X1    g0046(.A(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n245), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(G58), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(new_n247), .ZN(new_n254));
  OR2_X1    g0054(.A1(new_n254), .A2(new_n201), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n255), .A2(G20), .B1(G159), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT3), .B(G33), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT7), .ZN(new_n259));
  NOR3_X1   g0059(.A1(new_n258), .A2(new_n259), .A3(G20), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT71), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT3), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n261), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n262), .A2(G33), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(new_n268), .A3(KEYINPUT71), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n266), .A2(new_n210), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n260), .B1(new_n270), .B2(new_n259), .ZN(new_n271));
  OAI211_X1 g0071(.A(KEYINPUT16), .B(new_n257), .C1(new_n271), .C2(new_n247), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n216), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT16), .ZN(new_n275));
  INV_X1    g0075(.A(new_n257), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n259), .B1(new_n258), .B2(G20), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n267), .A2(new_n268), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n247), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n275), .B1(new_n276), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n272), .A2(new_n274), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT8), .B(G58), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n210), .A2(G1), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  AOI211_X1 g0089(.A(new_n284), .B(new_n274), .C1(new_n289), .C2(KEYINPUT72), .ZN(new_n290));
  OR2_X1    g0090(.A1(new_n289), .A2(KEYINPUT72), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n290), .A2(new_n291), .B1(new_n284), .B2(new_n285), .ZN(new_n292));
  AND2_X1   g0092(.A1(new_n282), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G223), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(G1698), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(new_n267), .A3(new_n268), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT73), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G87), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n267), .A2(new_n268), .A3(G226), .A4(G1698), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n295), .A2(new_n267), .A3(new_n268), .A4(KEYINPUT73), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n298), .A2(new_n299), .A3(new_n300), .A4(new_n301), .ZN(new_n302));
  AND2_X1   g0102(.A1(G33), .A2(G41), .ZN(new_n303));
  NOR3_X1   g0103(.A1(new_n303), .A2(KEYINPUT68), .A3(new_n216), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT68), .ZN(new_n305));
  AND2_X1   g0105(.A1(G1), .A2(G13), .ZN(new_n306));
  NAND2_X1  g0106(.A1(G33), .A2(G41), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n302), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G179), .ZN(new_n311));
  INV_X1    g0111(.A(G274), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n312), .B1(new_n306), .B2(new_n307), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n307), .A2(G1), .A3(G13), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n314), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n316), .B1(new_n234), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n310), .A2(new_n311), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT74), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n310), .A2(new_n320), .ZN(new_n323));
  INV_X1    g0123(.A(G169), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n319), .B1(new_n302), .B2(new_n309), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT74), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n327), .A3(new_n311), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n322), .A2(new_n325), .A3(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(KEYINPUT18), .B1(new_n293), .B2(new_n329), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n322), .A2(new_n325), .A3(new_n328), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT18), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n282), .A2(new_n292), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G190), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n335), .A2(KEYINPUT75), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n335), .A2(KEYINPUT75), .ZN(new_n337));
  OR2_X1    g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n326), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(G200), .B2(new_n326), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n341), .A2(new_n282), .A3(new_n292), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT17), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n341), .A2(new_n282), .A3(KEYINPUT17), .A4(new_n292), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n330), .A2(new_n334), .A3(new_n344), .A4(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n316), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n318), .A2(KEYINPUT66), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT66), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n317), .A2(new_n350), .A3(new_n314), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n348), .B1(new_n352), .B2(G238), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT13), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n267), .A2(new_n268), .A3(G232), .A4(G1698), .ZN(new_n355));
  INV_X1    g0155(.A(G1698), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n267), .A2(new_n268), .A3(G226), .A4(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G33), .A2(G97), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n355), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n309), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n353), .A2(new_n354), .A3(new_n360), .ZN(new_n361));
  AND3_X1   g0161(.A1(new_n317), .A2(new_n350), .A3(new_n314), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n350), .B1(new_n317), .B2(new_n314), .ZN(new_n363));
  OAI21_X1  g0163(.A(G238), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n360), .A2(new_n364), .A3(new_n316), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(KEYINPUT13), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n361), .A2(new_n366), .A3(G190), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n284), .A2(new_n247), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n368), .B(KEYINPUT12), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n256), .A2(G50), .B1(G20), .B2(new_n247), .ZN(new_n370));
  INV_X1    g0170(.A(G77), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n210), .A2(G33), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n373), .A2(KEYINPUT11), .A3(new_n274), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n284), .A2(new_n274), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n375), .A2(G68), .A3(new_n288), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n369), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT11), .B1(new_n373), .B2(new_n274), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n367), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G200), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n381), .B1(new_n361), .B2(new_n366), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n354), .B1(new_n353), .B2(new_n360), .ZN(new_n384));
  AND4_X1   g0184(.A1(new_n354), .A2(new_n360), .A3(new_n364), .A4(new_n316), .ZN(new_n385));
  OAI21_X1  g0185(.A(G169), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT14), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n361), .A2(new_n366), .A3(G179), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT14), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n389), .B(G169), .C1(new_n384), .C2(new_n385), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n387), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n379), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n383), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT67), .ZN(new_n394));
  INV_X1    g0194(.A(G226), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n395), .B1(new_n349), .B2(new_n351), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n394), .B1(new_n396), .B2(new_n348), .ZN(new_n397));
  OAI21_X1  g0197(.A(G226), .B1(new_n362), .B2(new_n363), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n398), .A2(KEYINPUT67), .A3(new_n316), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n258), .A2(G222), .A3(new_n356), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n258), .A2(G223), .A3(G1698), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n400), .B(new_n401), .C1(new_n371), .C2(new_n258), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n309), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n397), .A2(new_n399), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT70), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n405), .A3(G200), .ZN(new_n406));
  INV_X1    g0206(.A(new_n274), .ZN(new_n407));
  INV_X1    g0207(.A(new_n256), .ZN(new_n408));
  INV_X1    g0208(.A(G150), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n372), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n410), .B1(new_n286), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n210), .B1(new_n201), .B2(new_n202), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n407), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n287), .A2(new_n202), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n375), .A2(new_n416), .B1(new_n202), .B2(new_n284), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT9), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT9), .ZN(new_n420));
  AOI211_X1 g0220(.A(new_n413), .B(new_n410), .C1(new_n286), .C2(new_n411), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n420), .B(new_n417), .C1(new_n421), .C2(new_n407), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n397), .A2(G190), .A3(new_n399), .A4(new_n403), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n406), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n405), .B1(new_n404), .B2(G200), .ZN(new_n426));
  OAI21_X1  g0226(.A(KEYINPUT10), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n423), .A2(new_n424), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n404), .A2(G200), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT70), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT10), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n428), .A2(new_n430), .A3(new_n431), .A4(new_n406), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n427), .A2(new_n432), .ZN(new_n433));
  OR2_X1    g0233(.A1(new_n404), .A2(G179), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n417), .B1(new_n421), .B2(new_n407), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n404), .A2(new_n324), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  OAI22_X1  g0237(.A1(new_n285), .A2(new_n408), .B1(new_n210), .B2(new_n371), .ZN(new_n438));
  XNOR2_X1  g0238(.A(KEYINPUT15), .B(G87), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n439), .A2(new_n372), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n274), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n287), .A2(new_n371), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n375), .A2(new_n442), .B1(new_n371), .B2(new_n284), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n267), .A2(new_n268), .A3(G232), .A4(new_n356), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n267), .A2(new_n268), .A3(G238), .A4(G1698), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n445), .B(new_n446), .C1(new_n206), .C2(new_n258), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n309), .ZN(new_n448));
  OAI21_X1  g0248(.A(G244), .B1(new_n362), .B2(new_n363), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(new_n316), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n444), .B1(new_n450), .B2(G200), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT69), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n348), .B1(new_n352), .B2(G244), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n381), .B1(new_n454), .B2(new_n448), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT69), .B1(new_n455), .B2(new_n444), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n454), .A2(G190), .A3(new_n448), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n453), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n450), .A2(new_n324), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n454), .A2(new_n311), .A3(new_n448), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(new_n444), .A3(new_n460), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n437), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n347), .A2(new_n393), .A3(new_n433), .A4(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(G13), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(G1), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n210), .A2(G107), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT85), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT25), .ZN(new_n469));
  OR2_X1    g0269(.A1(new_n468), .A2(KEYINPUT25), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(KEYINPUT25), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n470), .A2(new_n465), .A3(new_n471), .A4(new_n466), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n209), .A2(G33), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n283), .A2(new_n473), .A3(new_n216), .A4(new_n273), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n469), .B(new_n472), .C1(new_n206), .C2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT86), .ZN(new_n476));
  OR2_X1    g0276(.A1(new_n474), .A2(new_n206), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT86), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n477), .A2(new_n478), .A3(new_n469), .A4(new_n472), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT23), .B1(new_n206), .B2(G20), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G116), .ZN(new_n483));
  OAI22_X1  g0283(.A1(new_n481), .A2(new_n482), .B1(G20), .B2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n267), .A2(new_n268), .A3(new_n210), .A4(G87), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT22), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT22), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n258), .A2(new_n487), .A3(new_n210), .A4(G87), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n484), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT24), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n274), .B1(new_n489), .B2(KEYINPUT24), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n480), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n267), .A2(new_n268), .A3(G250), .A4(new_n356), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT87), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n258), .A2(KEYINPUT87), .A3(G250), .A4(new_n356), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n267), .A2(new_n268), .A3(G257), .A4(G1698), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G33), .A2(G294), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n309), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G45), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(G1), .ZN(new_n504));
  NAND2_X1  g0304(.A1(KEYINPUT5), .A2(G41), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(KEYINPUT5), .A2(G41), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(G274), .B1(new_n303), .B2(new_n216), .ZN(new_n509));
  OAI21_X1  g0309(.A(KEYINPUT77), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n209), .A2(G45), .ZN(new_n511));
  OR2_X1    g0311(.A1(KEYINPUT5), .A2(G41), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n511), .B1(new_n512), .B2(new_n505), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT77), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n513), .A2(new_n514), .A3(new_n313), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n508), .A2(new_n317), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G264), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n502), .A2(new_n311), .A3(new_n516), .A4(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n501), .B1(new_n496), .B2(new_n497), .ZN(new_n520));
  INV_X1    g0320(.A(new_n309), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n516), .B(new_n518), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n324), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n493), .A2(new_n519), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n258), .A2(G264), .A3(G1698), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n278), .A2(G303), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n267), .A2(new_n268), .A3(G257), .A4(new_n356), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n309), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n517), .A2(G270), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n529), .A2(new_n530), .A3(new_n516), .ZN(new_n531));
  INV_X1    g0331(.A(G116), .ZN(new_n532));
  OR2_X1    g0332(.A1(new_n474), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G283), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n534), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n532), .A2(G20), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n535), .A2(new_n274), .A3(new_n536), .ZN(new_n537));
  XOR2_X1   g0337(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n284), .A2(new_n532), .ZN(new_n540));
  NOR2_X1   g0340(.A1(KEYINPUT84), .A2(KEYINPUT20), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n535), .A2(new_n274), .A3(new_n536), .A4(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n533), .A2(new_n539), .A3(new_n540), .A4(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n531), .A2(KEYINPUT21), .A3(G169), .A4(new_n543), .ZN(new_n544));
  AOI22_X1  g0344(.A1(G270), .A2(new_n517), .B1(new_n510), .B2(new_n515), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n545), .A2(new_n543), .A3(G179), .A4(new_n529), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n531), .A2(G169), .A3(new_n543), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT21), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n524), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n258), .A2(G244), .A3(G1698), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n267), .A2(new_n268), .A3(G238), .A4(new_n356), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(new_n483), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n309), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT81), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n504), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n511), .A2(KEYINPUT81), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n557), .A2(new_n558), .A3(G250), .A4(new_n317), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n313), .A2(new_n504), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n563), .A2(new_n335), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT19), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n210), .B1(new_n358), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(G87), .B2(new_n207), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n267), .A2(new_n268), .A3(new_n210), .A4(G68), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n565), .B1(new_n372), .B2(new_n205), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n274), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n439), .A2(new_n284), .ZN(new_n572));
  INV_X1    g0372(.A(G87), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n571), .B(new_n572), .C1(new_n573), .C2(new_n474), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n381), .B1(new_n555), .B2(new_n562), .ZN(new_n575));
  NOR3_X1   g0375(.A1(new_n564), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  OR2_X1    g0376(.A1(new_n474), .A2(new_n439), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n571), .A2(new_n572), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT82), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT82), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n571), .A2(new_n580), .A3(new_n572), .A4(new_n577), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n563), .A2(G169), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n555), .A2(G179), .A3(new_n562), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n582), .A2(KEYINPUT83), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT83), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n579), .A2(new_n586), .A3(new_n581), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n576), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n267), .A2(new_n268), .A3(G244), .A4(new_n356), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT4), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n534), .ZN(new_n592));
  NAND2_X1  g0392(.A1(G250), .A2(G1698), .ZN(new_n593));
  NAND2_X1  g0393(.A1(KEYINPUT4), .A2(G244), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n593), .B1(new_n594), .B2(G1698), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n592), .B1(new_n258), .B2(new_n595), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n591), .A2(new_n596), .A3(KEYINPUT76), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT76), .B1(new_n591), .B2(new_n596), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n309), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n517), .A2(G257), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n600), .A2(new_n516), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n599), .A2(KEYINPUT78), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(KEYINPUT78), .B1(new_n599), .B2(new_n601), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n324), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n284), .A2(new_n205), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n474), .B2(new_n205), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n206), .B1(new_n277), .B2(new_n279), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  XNOR2_X1  g0408(.A(G97), .B(G107), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT6), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n610), .A2(new_n205), .A3(G107), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n614), .A2(G20), .B1(G77), .B2(new_n256), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n608), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n606), .B1(new_n616), .B2(new_n274), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT79), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n591), .A2(new_n596), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT76), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n591), .A2(new_n596), .A3(KEYINPUT76), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n521), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n600), .A2(new_n516), .A3(new_n311), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n618), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n599), .A2(new_n601), .A3(KEYINPUT79), .A4(new_n311), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n617), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n604), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT80), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT78), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n600), .A2(new_n516), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n630), .B1(new_n623), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n599), .A2(new_n601), .A3(KEYINPUT78), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(G190), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n612), .B1(new_n610), .B2(new_n609), .ZN(new_n635));
  OAI22_X1  g0435(.A1(new_n635), .A2(new_n210), .B1(new_n371), .B2(new_n408), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n274), .B1(new_n636), .B2(new_n607), .ZN(new_n637));
  INV_X1    g0437(.A(new_n606), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n599), .A2(new_n601), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n639), .B1(G200), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n634), .A2(new_n641), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n628), .A2(new_n629), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n629), .B1(new_n628), .B2(new_n642), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n588), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n489), .A2(KEYINPUT24), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n646), .A2(new_n274), .A3(new_n490), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n502), .A2(G190), .A3(new_n516), .A4(new_n518), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n522), .A2(G200), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n647), .A2(new_n648), .A3(new_n649), .A4(new_n480), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n531), .A2(G200), .ZN(new_n651));
  INV_X1    g0451(.A(new_n543), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n651), .B(new_n652), .C1(new_n339), .C2(new_n531), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NOR4_X1   g0454(.A1(new_n463), .A2(new_n551), .A3(new_n645), .A4(new_n654), .ZN(G372));
  NAND2_X1  g0455(.A1(new_n330), .A2(new_n334), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n344), .A2(new_n345), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n390), .A2(new_n388), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n361), .A2(new_n366), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n389), .B1(new_n659), .B2(G169), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n392), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n383), .B2(new_n461), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n657), .B1(new_n662), .B2(KEYINPUT88), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT88), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n661), .B(new_n664), .C1(new_n383), .C2(new_n461), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n656), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT89), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n433), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n427), .A2(KEYINPUT89), .A3(new_n432), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n437), .B1(new_n666), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT90), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI211_X1 g0473(.A(KEYINPUT90), .B(new_n437), .C1(new_n666), .C2(new_n670), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n463), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n583), .A2(new_n584), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n582), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  OR3_X1    g0479(.A1(new_n564), .A2(new_n574), .A3(new_n575), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n650), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n547), .A2(new_n550), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n681), .B1(new_n682), .B2(new_n524), .ZN(new_n683));
  AOI22_X1  g0483(.A1(new_n604), .A2(new_n627), .B1(new_n634), .B2(new_n641), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n679), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n628), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n686), .A2(new_n588), .A3(KEYINPUT26), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT26), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n680), .A2(new_n678), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n688), .B1(new_n628), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n676), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n675), .A2(new_n693), .ZN(G369));
  INV_X1    g0494(.A(KEYINPUT91), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n465), .A2(new_n695), .A3(new_n210), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT91), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT92), .B1(new_n699), .B2(KEYINPUT27), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT92), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT27), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n696), .A2(new_n698), .A3(new_n701), .A4(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT93), .ZN(new_n705));
  INV_X1    g0505(.A(G213), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n706), .B1(new_n699), .B2(KEYINPUT27), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n705), .B1(new_n704), .B2(new_n707), .ZN(new_n710));
  XNOR2_X1  g0510(.A(KEYINPUT94), .B(G343), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n543), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n682), .B(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n714), .A2(G330), .A3(new_n653), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n712), .A2(new_n493), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n650), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n524), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n524), .A2(new_n712), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n716), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n682), .A2(new_n712), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n720), .B1(new_n719), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n724), .A2(new_n726), .ZN(G399));
  INV_X1    g0527(.A(new_n213), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G41), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(G1), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(new_n219), .B2(new_n730), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT28), .ZN(new_n734));
  INV_X1    g0534(.A(new_n712), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n692), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(KEYINPUT29), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT29), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n686), .A2(new_n588), .A3(new_n688), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n680), .A2(new_n650), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n684), .A2(new_n551), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(KEYINPUT26), .B1(new_n628), .B2(new_n689), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n739), .A2(new_n741), .A3(new_n678), .A4(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n738), .B1(new_n743), .B2(new_n735), .ZN(new_n744));
  INV_X1    g0544(.A(G330), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n545), .A2(G179), .A3(new_n529), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n563), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n502), .A2(new_n518), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n747), .A2(new_n632), .A3(new_n749), .A4(new_n633), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT30), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n748), .A2(new_n746), .A3(new_n563), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n753), .A2(KEYINPUT30), .A3(new_n632), .A4(new_n633), .ZN(new_n754));
  AOI21_X1  g0554(.A(G179), .B1(new_n545), .B2(new_n529), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n640), .A2(new_n755), .A3(new_n522), .A4(new_n563), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n752), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  AND3_X1   g0557(.A1(new_n757), .A2(KEYINPUT31), .A3(new_n712), .ZN(new_n758));
  AOI21_X1  g0558(.A(KEYINPUT31), .B1(new_n757), .B2(new_n712), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n551), .A2(new_n654), .A3(new_n712), .ZN(new_n761));
  OAI211_X1 g0561(.A(new_n588), .B(new_n761), .C1(new_n643), .C2(new_n644), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n745), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n737), .A2(new_n744), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n734), .B1(new_n764), .B2(G1), .ZN(G364));
  NAND2_X1  g0565(.A1(new_n714), .A2(new_n653), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(new_n745), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n464), .A2(G20), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n209), .B1(new_n768), .B2(G45), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n729), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n767), .A2(new_n715), .A3(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT95), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n766), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n213), .A2(G355), .A3(new_n258), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n266), .A2(new_n269), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n728), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(G45), .B2(new_n219), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n251), .A2(new_n503), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n779), .B1(G116), .B2(new_n213), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n306), .B1(new_n210), .B2(G169), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n785), .A2(KEYINPUT96), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(KEYINPUT96), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n777), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n772), .B1(new_n784), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n788), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n210), .A2(new_n311), .A3(new_n381), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n338), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n210), .A2(new_n311), .A3(G200), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n335), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n794), .A2(G50), .B1(G77), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n338), .A2(new_n795), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n253), .B2(new_n799), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT97), .Z(new_n801));
  NAND2_X1  g0601(.A1(new_n311), .A2(G200), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT98), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n804), .A2(new_n210), .A3(G190), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G107), .ZN(new_n806));
  NOR2_X1   g0606(.A1(G179), .A2(G200), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G190), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(G20), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G97), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n806), .A2(new_n258), .A3(new_n810), .ZN(new_n811));
  NOR3_X1   g0611(.A1(new_n804), .A2(new_n210), .A3(new_n335), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n573), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n807), .A2(G20), .A3(new_n335), .ZN(new_n815));
  INV_X1    g0615(.A(G159), .ZN(new_n816));
  NOR3_X1   g0616(.A1(new_n815), .A2(KEYINPUT32), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(KEYINPUT32), .B1(new_n815), .B2(new_n816), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n792), .A2(new_n335), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n818), .B1(new_n819), .B2(new_n247), .ZN(new_n820));
  NOR4_X1   g0620(.A1(new_n811), .A2(new_n814), .A3(new_n817), .A4(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G311), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n796), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G326), .ZN(new_n824));
  INV_X1    g0624(.A(G294), .ZN(new_n825));
  INV_X1    g0625(.A(new_n809), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n793), .A2(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n819), .ZN(new_n828));
  XNOR2_X1  g0628(.A(KEYINPUT33), .B(G317), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n823), .B(new_n827), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n799), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(G322), .ZN(new_n832));
  INV_X1    g0632(.A(new_n815), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n258), .B1(new_n833), .B2(G329), .ZN(new_n834));
  INV_X1    g0634(.A(G303), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n832), .B(new_n834), .C1(new_n835), .C2(new_n813), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G283), .B2(new_n805), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n801), .A2(new_n821), .B1(new_n830), .B2(new_n837), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n778), .B(new_n790), .C1(new_n791), .C2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n774), .A2(new_n839), .ZN(G396));
  INV_X1    g0640(.A(new_n461), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n704), .A2(new_n707), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(KEYINPUT93), .ZN(new_n843));
  INV_X1    g0643(.A(new_n711), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n843), .A2(new_n444), .A3(new_n708), .A4(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n841), .B1(new_n458), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n712), .A2(new_n461), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT101), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n457), .B1(new_n451), .B2(new_n452), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n455), .A2(KEYINPUT69), .A3(new_n444), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n845), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n461), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT101), .ZN(new_n853));
  INV_X1    g0653(.A(new_n847), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n848), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n736), .A2(new_n856), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n848), .A2(new_n855), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n692), .A2(new_n735), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n757), .A2(new_n712), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT31), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n757), .A2(KEYINPUT31), .A3(new_n712), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n762), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(G330), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n771), .B1(new_n860), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n866), .B2(new_n860), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n791), .A2(new_n776), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n771), .B1(new_n869), .B2(G77), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT99), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n794), .A2(G303), .B1(G283), .B2(new_n828), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n872), .B1(new_n532), .B2(new_n796), .C1(new_n825), .C2(new_n799), .ZN(new_n873));
  INV_X1    g0673(.A(new_n805), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n874), .A2(new_n573), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n813), .A2(new_n206), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n810), .B(new_n278), .C1(new_n822), .C2(new_n815), .ZN(new_n877));
  NOR4_X1   g0677(.A1(new_n873), .A2(new_n875), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n874), .A2(new_n247), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(G50), .B2(new_n812), .ZN(new_n880));
  INV_X1    g0680(.A(new_n780), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n881), .B1(G132), .B2(new_n833), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n880), .B(new_n882), .C1(new_n253), .C2(new_n826), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT34), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n794), .A2(G137), .B1(G159), .B2(new_n797), .ZN(new_n885));
  XOR2_X1   g0685(.A(KEYINPUT100), .B(G143), .Z(new_n886));
  OAI221_X1 g0686(.A(new_n885), .B1(new_n409), .B2(new_n819), .C1(new_n799), .C2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n883), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n887), .A2(new_n884), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n878), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI221_X1 g0690(.A(new_n871), .B1(new_n791), .B2(new_n890), .C1(new_n858), .C2(new_n776), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n868), .A2(new_n891), .ZN(G384));
  OR2_X1    g0692(.A1(new_n614), .A2(KEYINPUT35), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n614), .A2(KEYINPUT35), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n893), .A2(G116), .A3(new_n217), .A4(new_n894), .ZN(new_n895));
  XOR2_X1   g0695(.A(new_n895), .B(KEYINPUT36), .Z(new_n896));
  OR3_X1    g0696(.A1(new_n219), .A2(new_n371), .A3(new_n254), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n209), .B(G13), .C1(new_n897), .C2(new_n246), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT40), .ZN(new_n900));
  INV_X1    g0700(.A(new_n383), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n712), .A2(new_n392), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n661), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n392), .B(new_n712), .C1(new_n391), .C2(new_n383), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n905), .A2(new_n856), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n331), .A2(new_n333), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT37), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n709), .A2(new_n710), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n333), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n907), .A2(new_n908), .A3(new_n910), .A4(new_n342), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n257), .B1(new_n271), .B2(new_n247), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n275), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(new_n274), .A3(new_n272), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n329), .B1(new_n292), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n843), .A2(new_n708), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n914), .B2(new_n292), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n341), .A2(new_n282), .A3(new_n292), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n915), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n911), .B1(new_n919), .B2(new_n908), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n346), .A2(new_n917), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n920), .A2(KEYINPUT38), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT38), .B1(new_n920), .B2(new_n921), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n865), .B(new_n906), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n865), .A2(new_n906), .A3(KEYINPUT40), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n907), .A2(new_n342), .A3(new_n910), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(KEYINPUT37), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n911), .ZN(new_n928));
  INV_X1    g0728(.A(new_n910), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n346), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  XOR2_X1   g0731(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n920), .A2(new_n921), .A3(KEYINPUT38), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n900), .A2(new_n924), .B1(new_n925), .B2(new_n935), .ZN(new_n936));
  AND3_X1   g0736(.A1(new_n936), .A2(new_n676), .A3(new_n865), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n936), .B1(new_n676), .B2(new_n865), .ZN(new_n938));
  NOR3_X1   g0738(.A1(new_n937), .A2(new_n938), .A3(new_n745), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT104), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n859), .A2(new_n854), .ZN(new_n941));
  INV_X1    g0741(.A(new_n905), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n941), .B(new_n942), .C1(new_n923), .C2(new_n922), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT39), .ZN(new_n944));
  INV_X1    g0744(.A(new_n932), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n928), .B2(new_n930), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n944), .B1(new_n922), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n920), .A2(new_n921), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT38), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n950), .A2(KEYINPUT39), .A3(new_n934), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n391), .A2(new_n392), .A3(new_n735), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT102), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n947), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n656), .A2(new_n916), .ZN(new_n956));
  AND3_X1   g0756(.A1(new_n943), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n676), .B1(new_n737), .B2(new_n744), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n675), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n957), .B(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n940), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(G1), .B1(new_n464), .B2(G20), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n961), .A2(KEYINPUT105), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n940), .B2(new_n960), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT105), .B1(new_n961), .B2(new_n962), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n899), .B1(new_n964), .B2(new_n965), .ZN(G367));
  NAND2_X1  g0766(.A1(new_n712), .A2(new_n574), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n689), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n679), .B2(new_n967), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT106), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(KEYINPUT107), .B1(new_n971), .B2(KEYINPUT43), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT107), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT43), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n970), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n725), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n722), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n684), .B1(new_n617), .B2(new_n735), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n686), .A2(new_n712), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n982), .A2(KEYINPUT42), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n628), .B1(new_n979), .B2(new_n524), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n735), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n982), .A2(KEYINPUT42), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n983), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n976), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n976), .B1(new_n987), .B2(new_n988), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n716), .A2(new_n723), .A3(new_n981), .ZN(new_n992));
  NOR3_X1   g0792(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n992), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n987), .A2(new_n988), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n995), .A2(new_n975), .A3(new_n972), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n994), .B1(new_n996), .B2(new_n989), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n993), .A2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n729), .B(KEYINPUT41), .Z(new_n999));
  NOR2_X1   g0799(.A1(new_n737), .A2(new_n744), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n978), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n722), .A2(new_n977), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n716), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1001), .A2(new_n715), .A3(new_n1002), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1000), .A2(new_n1006), .A3(new_n866), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(KEYINPUT108), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n726), .A2(new_n981), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT45), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT44), .ZN(new_n1012));
  OR3_X1    g0812(.A1(new_n981), .A2(new_n726), .A3(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1012), .B1(new_n726), .B2(new_n981), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AND3_X1   g0815(.A1(new_n1011), .A2(new_n1015), .A3(new_n724), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n724), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT108), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n764), .A2(new_n1019), .A3(new_n1006), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1008), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n999), .B1(new_n1021), .B2(new_n764), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n998), .B1(new_n1022), .B2(new_n770), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n789), .B1(new_n213), .B2(new_n439), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n781), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1025), .A2(new_n240), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n771), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT46), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n813), .B2(new_n532), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n812), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n831), .A2(G303), .B1(G283), .B2(new_n797), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n828), .A2(G294), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n794), .A2(G311), .B1(G107), .B2(new_n809), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n780), .B1(G317), .B2(new_n833), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(new_n205), .C2(new_n874), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n826), .A2(new_n247), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n886), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1037), .B1(new_n794), .B2(new_n1038), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n202), .B2(new_n796), .C1(new_n816), .C2(new_n819), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n805), .A2(G77), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n812), .A2(G58), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n831), .A2(G150), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n278), .B1(new_n833), .B2(G137), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n1033), .A2(new_n1036), .B1(new_n1040), .B2(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT109), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT47), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n791), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1027), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n777), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1051), .B1(new_n971), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1023), .A2(new_n1053), .ZN(G387));
  INV_X1    g0854(.A(new_n731), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1055), .A2(new_n213), .A3(new_n258), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(G107), .B2(new_n213), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n237), .A2(new_n503), .ZN(new_n1058));
  AOI211_X1 g0858(.A(G45), .B(new_n1055), .C1(G68), .C2(G77), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n285), .A2(G50), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT50), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1025), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1057), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n789), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n771), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n874), .A2(new_n205), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n831), .A2(G50), .B1(G68), .B2(new_n797), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1067), .B(new_n780), .C1(new_n409), .C2(new_n815), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n439), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n809), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1070), .B1(new_n285), .B2(new_n819), .C1(new_n793), .C2(new_n816), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n813), .A2(new_n371), .ZN(new_n1072));
  OR4_X1    g0872(.A1(new_n1066), .A2(new_n1068), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(G317), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n799), .A2(new_n1074), .B1(new_n835), .B2(new_n796), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT110), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  OAI221_X1 g0877(.A(KEYINPUT110), .B1(new_n835), .B2(new_n796), .C1(new_n799), .C2(new_n1074), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n794), .A2(G322), .B1(G311), .B2(new_n828), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT48), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n812), .A2(G294), .B1(G283), .B2(new_n809), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT49), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n881), .B1(new_n824), .B2(new_n815), .C1(new_n874), .C2(new_n532), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1073), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1065), .B1(new_n1091), .B2(new_n788), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT111), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1094), .B(new_n1095), .C1(new_n722), .C2(new_n777), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n770), .B2(new_n1006), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n764), .A2(new_n1006), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(KEYINPUT112), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1099), .A2(new_n729), .A3(new_n1007), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1098), .A2(KEYINPUT112), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1097), .B1(new_n1100), .B2(new_n1101), .ZN(G393));
  AND2_X1   g0902(.A1(new_n764), .A2(new_n1006), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1021), .B(new_n729), .C1(new_n1103), .C2(new_n1018), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1018), .A2(new_n770), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1064), .B1(G97), .B2(new_n728), .ZN(new_n1106));
  OR2_X1    g0906(.A1(new_n1025), .A2(new_n244), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n772), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n826), .A2(new_n371), .B1(new_n819), .B2(new_n202), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n881), .B(new_n875), .C1(new_n833), .C2(new_n1038), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n247), .B2(new_n813), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1109), .B(new_n1111), .C1(new_n286), .C2(new_n797), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n409), .A2(new_n793), .B1(new_n799), .B2(new_n816), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT51), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n797), .A2(G294), .B1(G116), .B2(new_n809), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n835), .B2(new_n819), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT113), .Z(new_n1117));
  AOI21_X1  g0917(.A(new_n258), .B1(new_n833), .B2(G322), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n806), .A2(new_n1118), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n822), .A2(new_n799), .B1(new_n793), .B2(new_n1074), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT52), .Z(new_n1121));
  AOI211_X1 g0921(.A(new_n1119), .B(new_n1121), .C1(G283), .C2(new_n812), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1112), .A2(new_n1114), .B1(new_n1117), .B2(new_n1122), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1108), .B1(new_n1052), .B2(new_n981), .C1(new_n1123), .C2(new_n791), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1104), .A2(new_n1105), .A3(new_n1124), .ZN(G390));
  AND4_X1   g0925(.A1(G330), .A2(new_n865), .A3(new_n858), .A4(new_n942), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n858), .A2(new_n743), .A3(new_n735), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n854), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n942), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n954), .B1(new_n933), .B2(new_n934), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n712), .B1(new_n685), .B2(new_n691), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n847), .B1(new_n1131), .B2(new_n858), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n953), .B1(new_n1132), .B2(new_n905), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n947), .A2(new_n951), .ZN(new_n1134));
  AOI221_X4 g0934(.A(new_n1126), .B1(new_n1129), .B2(new_n1130), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n763), .A2(new_n858), .A3(new_n942), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1136), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n770), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n771), .B1(new_n869), .B2(new_n286), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n794), .A2(G283), .B1(G107), .B2(new_n828), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1143), .B1(new_n205), .B2(new_n796), .C1(new_n532), .C2(new_n799), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n278), .B1(new_n815), .B2(new_n825), .C1(new_n826), .C2(new_n371), .ZN(new_n1145));
  NOR4_X1   g0945(.A1(new_n1144), .A2(new_n814), .A3(new_n879), .A4(new_n1145), .ZN(new_n1146));
  OR2_X1    g0946(.A1(new_n1146), .A2(KEYINPUT116), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(KEYINPUT116), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n812), .A2(G150), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT53), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n794), .A2(G128), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n278), .B1(new_n833), .B2(G125), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1151), .B(new_n1152), .C1(new_n202), .C2(new_n874), .ZN(new_n1153));
  INV_X1    g0953(.A(G137), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n826), .A2(new_n816), .B1(new_n819), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(G132), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT54), .B(G143), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n799), .A2(new_n1156), .B1(new_n796), .B2(new_n1157), .ZN(new_n1158));
  OR4_X1    g0958(.A1(new_n1150), .A2(new_n1153), .A3(new_n1155), .A4(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1147), .A2(new_n1148), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1142), .B1(new_n1160), .B2(new_n788), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1134), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1161), .B1(new_n1162), .B2(new_n776), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT117), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1141), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n905), .B1(new_n866), .B2(new_n856), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1132), .B1(new_n1166), .B2(new_n1136), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n858), .B1(new_n866), .B2(KEYINPUT114), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT114), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n763), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n905), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1167), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n763), .A2(new_n676), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n675), .A2(new_n958), .A3(new_n1174), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n1173), .A2(new_n1175), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n941), .A2(new_n942), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1177), .A2(new_n953), .B1(new_n947), .B2(new_n951), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1138), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1126), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1175), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n942), .B1(new_n763), .B2(new_n858), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n941), .B1(new_n1182), .B2(new_n1126), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n856), .B1(new_n763), .B2(new_n1169), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n866), .A2(KEYINPUT114), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n942), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1136), .A2(new_n854), .A3(new_n1127), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1183), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1137), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1180), .A2(new_n1181), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1176), .A2(new_n729), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(KEYINPUT115), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT115), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1176), .A2(new_n1190), .A3(new_n1193), .A4(new_n729), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1165), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(G378));
  AOI211_X1 g0996(.A(new_n1037), .B(new_n1072), .C1(G283), .C2(new_n833), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n780), .A2(G41), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1197), .B(new_n1198), .C1(new_n253), .C2(new_n874), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n828), .A2(G97), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n797), .A2(new_n1069), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(new_n206), .B2(new_n799), .C1(new_n532), .C2(new_n793), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1199), .A2(new_n1203), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1204), .A2(KEYINPUT58), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(KEYINPUT58), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1205), .B(new_n1206), .C1(new_n1198), .C2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n796), .A2(new_n1154), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n826), .A2(new_n409), .B1(new_n819), .B2(new_n1156), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1209), .B(new_n1210), .C1(G125), .C2(new_n794), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1157), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n812), .A2(new_n1212), .B1(new_n831), .B2(G128), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT118), .ZN(new_n1214));
  AND2_X1   g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1211), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1217), .A2(KEYINPUT59), .ZN(new_n1218));
  AOI211_X1 g1018(.A(G33), .B(G41), .C1(new_n833), .C2(G124), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n874), .B2(new_n816), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n1217), .B2(KEYINPUT59), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1208), .B1(new_n1218), .B2(new_n1221), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n771), .B1(G50), .B2(new_n869), .C1(new_n1222), .C2(new_n791), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n909), .A2(new_n435), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n427), .A2(KEYINPUT89), .A3(new_n432), .ZN(new_n1228));
  AOI21_X1  g1028(.A(KEYINPUT89), .B1(new_n427), .B2(new_n432), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1227), .B1(new_n1230), .B2(new_n437), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n437), .ZN(new_n1232));
  NOR4_X1   g1032(.A1(new_n1228), .A2(new_n1229), .A3(new_n1232), .A4(new_n1226), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1225), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1226), .B1(new_n670), .B2(new_n1232), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1230), .A2(new_n437), .A3(new_n1227), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(new_n1236), .A3(new_n1224), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1234), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1223), .B1(new_n1239), .B2(new_n775), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1238), .B1(new_n936), .B2(G330), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n922), .A2(new_n923), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n865), .A2(new_n906), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n900), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n935), .A2(KEYINPUT40), .A3(new_n865), .A4(new_n906), .ZN(new_n1245));
  AND4_X1   g1045(.A1(G330), .A2(new_n1244), .A3(new_n1238), .A4(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(KEYINPUT119), .B1(new_n1241), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n957), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1244), .A2(new_n1245), .A3(G330), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n1239), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n936), .A2(G330), .A3(new_n1238), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n957), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1252), .A2(KEYINPUT119), .A3(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1248), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1240), .B1(new_n1255), .B2(new_n770), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1190), .A2(new_n1181), .ZN(new_n1257));
  AOI21_X1  g1057(.A(KEYINPUT57), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1250), .A2(new_n1251), .A3(new_n957), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n957), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1260));
  OAI21_X1  g1060(.A(KEYINPUT57), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1175), .B1(new_n1140), .B2(new_n1188), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n729), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1256), .B1(new_n1258), .B2(new_n1263), .ZN(G375));
  NAND2_X1  g1064(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1181), .A2(new_n1188), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n999), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1268));
  XOR2_X1   g1068(.A(new_n1268), .B(KEYINPUT120), .Z(new_n1269));
  OAI21_X1  g1069(.A(new_n771), .B1(new_n869), .B2(G68), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n258), .B1(new_n833), .B2(G303), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1041), .A2(new_n1070), .A3(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n831), .A2(G283), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n797), .A2(G107), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  OAI221_X1 g1075(.A(new_n1275), .B1(new_n532), .B2(new_n819), .C1(new_n825), .C2(new_n793), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n1272), .B(new_n1276), .C1(G97), .C2(new_n812), .ZN(new_n1277));
  OR2_X1    g1077(.A1(new_n1277), .A2(KEYINPUT121), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(KEYINPUT121), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(G58), .A2(new_n805), .B1(new_n812), .B2(G159), .ZN(new_n1280));
  OAI22_X1  g1080(.A1(new_n826), .A2(new_n202), .B1(new_n796), .B2(new_n409), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(G132), .B2(new_n794), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n831), .A2(G137), .B1(new_n828), .B2(new_n1212), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n881), .B1(G128), .B2(new_n833), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1280), .A2(new_n1282), .A3(new_n1283), .A4(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1278), .A2(new_n1279), .A3(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1270), .B1(new_n1286), .B2(new_n788), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1287), .B1(new_n942), .B2(new_n776), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1288), .B1(new_n1173), .B2(new_n769), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1269), .A2(new_n1290), .ZN(G381));
  INV_X1    g1091(.A(G396), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1097), .B(new_n1292), .C1(new_n1101), .C2(new_n1100), .ZN(new_n1293));
  OR4_X1    g1093(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1293), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1191), .A2(new_n1164), .A3(new_n1141), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  NOR4_X1   g1096(.A1(new_n1294), .A2(G375), .A3(G381), .A4(new_n1296), .ZN(new_n1297));
  XOR2_X1   g1097(.A(new_n1297), .B(KEYINPUT122), .Z(G407));
  NOR2_X1   g1098(.A1(new_n844), .A2(new_n706), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1299), .B(KEYINPUT123), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1295), .A2(new_n1300), .ZN(new_n1301));
  OAI211_X1 g1101(.A(G407), .B(G213), .C1(G375), .C2(new_n1301), .ZN(G409));
  INV_X1    g1102(.A(G390), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(G387), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(G393), .A2(G396), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1293), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1023), .A2(G390), .A3(new_n1053), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1304), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  AND3_X1   g1109(.A1(new_n1023), .A2(G390), .A3(new_n1053), .ZN(new_n1310));
  AOI21_X1  g1110(.A(G390), .B1(new_n1023), .B2(new_n1053), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1306), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1309), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1254), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1253), .B1(new_n1252), .B2(KEYINPUT119), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n1257), .B(new_n1267), .C1(new_n1314), .C2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1250), .A2(new_n1251), .A3(new_n957), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1240), .B1(new_n1319), .B2(new_n770), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1316), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1295), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1322), .B1(G375), .B2(new_n1195), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1300), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT60), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1326), .B1(new_n1181), .B2(new_n1188), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1181), .A2(new_n1188), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n729), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT125), .ZN(new_n1330));
  NOR3_X1   g1130(.A1(new_n1181), .A2(new_n1188), .A3(new_n1326), .ZN(new_n1331));
  NOR3_X1   g1131(.A1(new_n1329), .A2(new_n1330), .A3(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(KEYINPUT60), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n730), .B1(new_n1333), .B2(new_n1265), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1331), .ZN(new_n1335));
  AOI21_X1  g1135(.A(KEYINPUT125), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1290), .B1(new_n1332), .B2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(G384), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1330), .B1(new_n1329), .B2(new_n1331), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1334), .A2(KEYINPUT125), .A3(new_n1335), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1342), .A2(G384), .A3(new_n1290), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1339), .A2(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT62), .ZN(new_n1345));
  NOR3_X1   g1145(.A1(new_n1325), .A2(new_n1344), .A3(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1323), .A2(KEYINPUT124), .ZN(new_n1347));
  AOI21_X1  g1147(.A(G384), .B1(new_n1342), .B2(new_n1290), .ZN(new_n1348));
  AOI211_X1 g1148(.A(new_n1338), .B(new_n1289), .C1(new_n1340), .C2(new_n1341), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT124), .ZN(new_n1351));
  OAI211_X1 g1151(.A(new_n1322), .B(new_n1351), .C1(G375), .C2(new_n1195), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1347), .A2(new_n1324), .A3(new_n1350), .A4(new_n1352), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1346), .B1(new_n1345), .B2(new_n1353), .ZN(new_n1354));
  NAND4_X1  g1154(.A1(new_n1339), .A2(G2897), .A3(new_n1300), .A4(new_n1343), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1300), .A2(G2897), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1356), .B1(new_n1348), .B2(new_n1349), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1355), .A2(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1358), .A2(new_n1325), .ZN(new_n1359));
  INV_X1    g1159(.A(KEYINPUT61), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1359), .A2(new_n1360), .ZN(new_n1361));
  OAI21_X1  g1161(.A(new_n1313), .B1(new_n1354), .B2(new_n1361), .ZN(new_n1362));
  AND3_X1   g1162(.A1(new_n1309), .A2(new_n1312), .A3(new_n1360), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1339), .A2(KEYINPUT63), .A3(new_n1343), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1363), .B1(new_n1325), .B2(new_n1364), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1347), .A2(new_n1324), .A3(new_n1352), .ZN(new_n1366));
  AOI21_X1  g1166(.A(new_n1365), .B1(new_n1366), .B2(new_n1358), .ZN(new_n1367));
  XOR2_X1   g1167(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1368));
  NAND2_X1  g1168(.A1(new_n1353), .A2(new_n1368), .ZN(new_n1369));
  AOI21_X1  g1169(.A(KEYINPUT127), .B1(new_n1367), .B2(new_n1369), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1366), .A2(new_n1358), .ZN(new_n1371));
  NAND3_X1  g1171(.A1(new_n1309), .A2(new_n1312), .A3(new_n1360), .ZN(new_n1372));
  INV_X1    g1172(.A(new_n1325), .ZN(new_n1373));
  INV_X1    g1173(.A(new_n1364), .ZN(new_n1374));
  AOI21_X1  g1174(.A(new_n1372), .B1(new_n1373), .B2(new_n1374), .ZN(new_n1375));
  AND4_X1   g1175(.A1(KEYINPUT127), .A2(new_n1369), .A3(new_n1371), .A4(new_n1375), .ZN(new_n1376));
  OAI21_X1  g1176(.A(new_n1362), .B1(new_n1370), .B2(new_n1376), .ZN(G405));
  AND2_X1   g1177(.A1(G375), .A2(new_n1295), .ZN(new_n1378));
  NOR2_X1   g1178(.A1(G375), .A2(new_n1195), .ZN(new_n1379));
  NOR2_X1   g1179(.A1(new_n1378), .A2(new_n1379), .ZN(new_n1380));
  XNOR2_X1  g1180(.A(new_n1380), .B(new_n1344), .ZN(new_n1381));
  XNOR2_X1  g1181(.A(new_n1381), .B(new_n1313), .ZN(G402));
endmodule


