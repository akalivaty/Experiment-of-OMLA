

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U546 ( .A(n725), .ZN(n709) );
  NOR2_X1 U547 ( .A1(n631), .A2(n515), .ZN(n647) );
  NOR2_X2 U548 ( .A1(G651), .A2(n631), .ZN(n644) );
  BUF_X2 U549 ( .A(n961), .Z(n508) );
  XNOR2_X1 U550 ( .A(n597), .B(n596), .ZN(n976) );
  XNOR2_X1 U551 ( .A(KEYINPUT75), .B(n577), .ZN(n961) );
  NOR2_X1 U552 ( .A1(n576), .A2(n575), .ZN(n577) );
  INV_X1 U553 ( .A(G2105), .ZN(n534) );
  XNOR2_X2 U554 ( .A(n535), .B(KEYINPUT64), .ZN(n544) );
  INV_X1 U555 ( .A(KEYINPUT13), .ZN(n572) );
  XOR2_X1 U556 ( .A(KEYINPUT89), .B(n530), .Z(n531) );
  NOR2_X2 U557 ( .A1(n548), .A2(n547), .ZN(G160) );
  XNOR2_X2 U558 ( .A(n521), .B(n520), .ZN(n586) );
  OR2_X1 U559 ( .A1(G299), .A2(n703), .ZN(n509) );
  OR2_X1 U560 ( .A1(n685), .A2(n684), .ZN(n510) );
  AND2_X1 U561 ( .A1(G8), .A2(n737), .ZN(n511) );
  AND2_X1 U562 ( .A1(n761), .A2(n764), .ZN(n512) );
  AND2_X1 U563 ( .A1(n767), .A2(n766), .ZN(n513) );
  AND2_X1 U564 ( .A1(n681), .A2(n683), .ZN(n682) );
  NOR2_X1 U565 ( .A1(n508), .A2(n510), .ZN(n687) );
  NOR2_X1 U566 ( .A1(n706), .A2(n705), .ZN(n707) );
  AND2_X1 U567 ( .A1(n736), .A2(n739), .ZN(n740) );
  NOR2_X1 U568 ( .A1(n512), .A2(n765), .ZN(n766) );
  INV_X1 U569 ( .A(KEYINPUT68), .ZN(n519) );
  XNOR2_X1 U570 ( .A(n519), .B(KEYINPUT1), .ZN(n520) );
  XNOR2_X1 U571 ( .A(n572), .B(KEYINPUT74), .ZN(n573) );
  INV_X1 U572 ( .A(KEYINPUT17), .ZN(n528) );
  XNOR2_X1 U573 ( .A(n574), .B(n573), .ZN(n575) );
  NAND2_X1 U574 ( .A1(n877), .A2(G137), .ZN(n540) );
  NOR2_X2 U575 ( .A1(G651), .A2(G543), .ZN(n651) );
  NAND2_X1 U576 ( .A1(n651), .A2(G89), .ZN(n514) );
  XNOR2_X1 U577 ( .A(n514), .B(KEYINPUT4), .ZN(n517) );
  XOR2_X1 U578 ( .A(KEYINPUT0), .B(G543), .Z(n631) );
  INV_X1 U579 ( .A(G651), .ZN(n515) );
  NAND2_X1 U580 ( .A1(G76), .A2(n647), .ZN(n516) );
  NAND2_X1 U581 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n518), .B(KEYINPUT5), .ZN(n526) );
  NAND2_X1 U583 ( .A1(n644), .A2(G51), .ZN(n523) );
  NOR2_X1 U584 ( .A1(n515), .A2(G543), .ZN(n521) );
  NAND2_X1 U585 ( .A1(G63), .A2(n586), .ZN(n522) );
  NAND2_X1 U586 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U587 ( .A(KEYINPUT6), .B(n524), .Z(n525) );
  NAND2_X1 U588 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U589 ( .A(n527), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U590 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U591 ( .A1(G2105), .A2(G2104), .ZN(n529) );
  XNOR2_X2 U592 ( .A(n529), .B(n528), .ZN(n877) );
  NAND2_X1 U593 ( .A1(n877), .A2(G138), .ZN(n532) );
  AND2_X2 U594 ( .A1(n534), .A2(G2104), .ZN(n876) );
  NAND2_X1 U595 ( .A1(G102), .A2(n876), .ZN(n530) );
  NAND2_X1 U596 ( .A1(n532), .A2(n531), .ZN(n539) );
  NAND2_X1 U597 ( .A1(G2104), .A2(G2105), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n533), .B(KEYINPUT65), .ZN(n871) );
  NAND2_X1 U599 ( .A1(G114), .A2(n871), .ZN(n537) );
  NOR2_X1 U600 ( .A1(n534), .A2(G2104), .ZN(n535) );
  NAND2_X1 U601 ( .A1(G126), .A2(n544), .ZN(n536) );
  NAND2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U603 ( .A1(n539), .A2(n538), .ZN(G164) );
  XNOR2_X1 U604 ( .A(n540), .B(KEYINPUT66), .ZN(n543) );
  NAND2_X1 U605 ( .A1(G101), .A2(n876), .ZN(n541) );
  XOR2_X1 U606 ( .A(KEYINPUT23), .B(n541), .Z(n542) );
  NAND2_X1 U607 ( .A1(n543), .A2(n542), .ZN(n548) );
  NAND2_X1 U608 ( .A1(G113), .A2(n871), .ZN(n546) );
  NAND2_X1 U609 ( .A1(G125), .A2(n544), .ZN(n545) );
  NAND2_X1 U610 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U611 ( .A1(n644), .A2(G53), .ZN(n550) );
  NAND2_X1 U612 ( .A1(G65), .A2(n586), .ZN(n549) );
  NAND2_X1 U613 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U614 ( .A1(G91), .A2(n651), .ZN(n552) );
  NAND2_X1 U615 ( .A1(G78), .A2(n647), .ZN(n551) );
  NAND2_X1 U616 ( .A1(n552), .A2(n551), .ZN(n553) );
  OR2_X1 U617 ( .A1(n554), .A2(n553), .ZN(G299) );
  AND2_X1 U618 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U619 ( .A(G132), .ZN(G219) );
  NAND2_X1 U620 ( .A1(G88), .A2(n651), .ZN(n556) );
  NAND2_X1 U621 ( .A1(G75), .A2(n647), .ZN(n555) );
  NAND2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U623 ( .A(KEYINPUT86), .B(n557), .Z(n561) );
  NAND2_X1 U624 ( .A1(n586), .A2(G62), .ZN(n559) );
  NAND2_X1 U625 ( .A1(n644), .A2(G50), .ZN(n558) );
  AND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(G303) );
  XOR2_X1 U628 ( .A(KEYINPUT72), .B(KEYINPUT11), .Z(n564) );
  NAND2_X1 U629 ( .A1(G7), .A2(G661), .ZN(n562) );
  XOR2_X1 U630 ( .A(n562), .B(KEYINPUT10), .Z(n907) );
  NAND2_X1 U631 ( .A1(G567), .A2(n907), .ZN(n563) );
  XNOR2_X1 U632 ( .A(n564), .B(n563), .ZN(G234) );
  NAND2_X1 U633 ( .A1(n586), .A2(G56), .ZN(n565) );
  XOR2_X1 U634 ( .A(KEYINPUT14), .B(n565), .Z(n566) );
  XNOR2_X1 U635 ( .A(n566), .B(KEYINPUT73), .ZN(n568) );
  NAND2_X1 U636 ( .A1(G43), .A2(n644), .ZN(n567) );
  NAND2_X1 U637 ( .A1(n568), .A2(n567), .ZN(n576) );
  NAND2_X1 U638 ( .A1(n651), .A2(G81), .ZN(n569) );
  XNOR2_X1 U639 ( .A(n569), .B(KEYINPUT12), .ZN(n571) );
  NAND2_X1 U640 ( .A1(G68), .A2(n647), .ZN(n570) );
  NAND2_X1 U641 ( .A1(n571), .A2(n570), .ZN(n574) );
  INV_X1 U642 ( .A(G860), .ZN(n602) );
  OR2_X1 U643 ( .A1(n508), .A2(n602), .ZN(G153) );
  NAND2_X1 U644 ( .A1(n586), .A2(G64), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n578), .B(KEYINPUT69), .ZN(n583) );
  NAND2_X1 U646 ( .A1(G90), .A2(n651), .ZN(n580) );
  NAND2_X1 U647 ( .A1(G77), .A2(n647), .ZN(n579) );
  NAND2_X1 U648 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U649 ( .A(KEYINPUT9), .B(n581), .Z(n582) );
  NOR2_X1 U650 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U651 ( .A1(n644), .A2(G52), .ZN(n584) );
  NAND2_X1 U652 ( .A1(n585), .A2(n584), .ZN(G301) );
  NAND2_X1 U653 ( .A1(G868), .A2(G301), .ZN(n599) );
  INV_X1 U654 ( .A(KEYINPUT15), .ZN(n597) );
  NAND2_X1 U655 ( .A1(G66), .A2(n586), .ZN(n587) );
  XNOR2_X1 U656 ( .A(n587), .B(KEYINPUT76), .ZN(n589) );
  NAND2_X1 U657 ( .A1(G92), .A2(n651), .ZN(n588) );
  NAND2_X1 U658 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U659 ( .A(n590), .B(KEYINPUT77), .ZN(n592) );
  NAND2_X1 U660 ( .A1(G79), .A2(n647), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U662 ( .A1(n644), .A2(G54), .ZN(n593) );
  XOR2_X1 U663 ( .A(KEYINPUT78), .B(n593), .Z(n594) );
  NOR2_X1 U664 ( .A1(n595), .A2(n594), .ZN(n596) );
  OR2_X1 U665 ( .A1(n976), .A2(G868), .ZN(n598) );
  NAND2_X1 U666 ( .A1(n599), .A2(n598), .ZN(G284) );
  NOR2_X1 U667 ( .A1(G868), .A2(G299), .ZN(n601) );
  INV_X1 U668 ( .A(G868), .ZN(n663) );
  NOR2_X1 U669 ( .A1(G286), .A2(n663), .ZN(n600) );
  NOR2_X1 U670 ( .A1(n601), .A2(n600), .ZN(G297) );
  NAND2_X1 U671 ( .A1(n602), .A2(G559), .ZN(n603) );
  NAND2_X1 U672 ( .A1(n603), .A2(n976), .ZN(n604) );
  XNOR2_X1 U673 ( .A(n604), .B(KEYINPUT16), .ZN(n605) );
  XOR2_X1 U674 ( .A(KEYINPUT79), .B(n605), .Z(G148) );
  NOR2_X1 U675 ( .A1(G868), .A2(n508), .ZN(n606) );
  XNOR2_X1 U676 ( .A(KEYINPUT80), .B(n606), .ZN(n609) );
  NAND2_X1 U677 ( .A1(G868), .A2(n976), .ZN(n607) );
  NOR2_X1 U678 ( .A1(G559), .A2(n607), .ZN(n608) );
  NOR2_X1 U679 ( .A1(n609), .A2(n608), .ZN(G282) );
  XOR2_X1 U680 ( .A(G2100), .B(KEYINPUT82), .Z(n619) );
  XOR2_X1 U681 ( .A(G2096), .B(KEYINPUT81), .Z(n617) );
  NAND2_X1 U682 ( .A1(n544), .A2(G123), .ZN(n610) );
  XNOR2_X1 U683 ( .A(n610), .B(KEYINPUT18), .ZN(n612) );
  NAND2_X1 U684 ( .A1(n876), .A2(G99), .ZN(n611) );
  NAND2_X1 U685 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U686 ( .A1(G135), .A2(n877), .ZN(n614) );
  NAND2_X1 U687 ( .A1(G111), .A2(n871), .ZN(n613) );
  NAND2_X1 U688 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U689 ( .A1(n616), .A2(n615), .ZN(n943) );
  XNOR2_X1 U690 ( .A(n617), .B(n943), .ZN(n618) );
  NAND2_X1 U691 ( .A1(n619), .A2(n618), .ZN(G156) );
  NAND2_X1 U692 ( .A1(n976), .A2(G559), .ZN(n661) );
  XNOR2_X1 U693 ( .A(n508), .B(n661), .ZN(n620) );
  NOR2_X1 U694 ( .A1(n620), .A2(G860), .ZN(n630) );
  NAND2_X1 U695 ( .A1(G67), .A2(n586), .ZN(n621) );
  XNOR2_X1 U696 ( .A(n621), .B(KEYINPUT84), .ZN(n623) );
  NAND2_X1 U697 ( .A1(G55), .A2(n644), .ZN(n622) );
  NAND2_X1 U698 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U699 ( .A(n624), .B(KEYINPUT85), .ZN(n626) );
  NAND2_X1 U700 ( .A1(G80), .A2(n647), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U702 ( .A1(G93), .A2(n651), .ZN(n627) );
  XNOR2_X1 U703 ( .A(KEYINPUT83), .B(n627), .ZN(n628) );
  OR2_X1 U704 ( .A1(n629), .A2(n628), .ZN(n664) );
  XOR2_X1 U705 ( .A(n630), .B(n664), .Z(G145) );
  NAND2_X1 U706 ( .A1(G87), .A2(n631), .ZN(n633) );
  NAND2_X1 U707 ( .A1(G74), .A2(G651), .ZN(n632) );
  NAND2_X1 U708 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U709 ( .A1(n586), .A2(n634), .ZN(n636) );
  NAND2_X1 U710 ( .A1(n644), .A2(G49), .ZN(n635) );
  NAND2_X1 U711 ( .A1(n636), .A2(n635), .ZN(G288) );
  NAND2_X1 U712 ( .A1(n644), .A2(G47), .ZN(n638) );
  NAND2_X1 U713 ( .A1(G60), .A2(n586), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U715 ( .A1(G85), .A2(n651), .ZN(n639) );
  XNOR2_X1 U716 ( .A(KEYINPUT67), .B(n639), .ZN(n640) );
  NOR2_X1 U717 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U718 ( .A1(n647), .A2(G72), .ZN(n642) );
  NAND2_X1 U719 ( .A1(n643), .A2(n642), .ZN(G290) );
  NAND2_X1 U720 ( .A1(n644), .A2(G48), .ZN(n646) );
  NAND2_X1 U721 ( .A1(G61), .A2(n586), .ZN(n645) );
  NAND2_X1 U722 ( .A1(n646), .A2(n645), .ZN(n650) );
  NAND2_X1 U723 ( .A1(n647), .A2(G73), .ZN(n648) );
  XOR2_X1 U724 ( .A(KEYINPUT2), .B(n648), .Z(n649) );
  NOR2_X1 U725 ( .A1(n650), .A2(n649), .ZN(n653) );
  NAND2_X1 U726 ( .A1(n651), .A2(G86), .ZN(n652) );
  NAND2_X1 U727 ( .A1(n653), .A2(n652), .ZN(G305) );
  XOR2_X1 U728 ( .A(KEYINPUT19), .B(KEYINPUT87), .Z(n654) );
  XNOR2_X1 U729 ( .A(G288), .B(n654), .ZN(n657) );
  XOR2_X1 U730 ( .A(G303), .B(G290), .Z(n655) );
  XNOR2_X1 U731 ( .A(n655), .B(G299), .ZN(n656) );
  XNOR2_X1 U732 ( .A(n657), .B(n656), .ZN(n659) );
  XOR2_X1 U733 ( .A(G305), .B(n664), .Z(n658) );
  XNOR2_X1 U734 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U735 ( .A(n660), .B(n508), .ZN(n888) );
  XOR2_X1 U736 ( .A(n888), .B(n661), .Z(n662) );
  NAND2_X1 U737 ( .A1(G868), .A2(n662), .ZN(n666) );
  NAND2_X1 U738 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U739 ( .A1(n666), .A2(n665), .ZN(G295) );
  NAND2_X1 U740 ( .A1(G2084), .A2(G2078), .ZN(n667) );
  XOR2_X1 U741 ( .A(KEYINPUT20), .B(n667), .Z(n668) );
  NAND2_X1 U742 ( .A1(G2090), .A2(n668), .ZN(n669) );
  XNOR2_X1 U743 ( .A(KEYINPUT21), .B(n669), .ZN(n670) );
  NAND2_X1 U744 ( .A1(n670), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U745 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U746 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  XOR2_X1 U747 ( .A(KEYINPUT70), .B(G57), .Z(G237) );
  NOR2_X1 U748 ( .A1(G219), .A2(G220), .ZN(n671) );
  XOR2_X1 U749 ( .A(KEYINPUT88), .B(n671), .Z(n672) );
  XNOR2_X1 U750 ( .A(n672), .B(KEYINPUT22), .ZN(n673) );
  NOR2_X1 U751 ( .A1(G218), .A2(n673), .ZN(n674) );
  NAND2_X1 U752 ( .A1(G96), .A2(n674), .ZN(n823) );
  NAND2_X1 U753 ( .A1(n823), .A2(G2106), .ZN(n678) );
  NAND2_X1 U754 ( .A1(G108), .A2(G120), .ZN(n675) );
  NOR2_X1 U755 ( .A1(G237), .A2(n675), .ZN(n676) );
  NAND2_X1 U756 ( .A1(G69), .A2(n676), .ZN(n822) );
  NAND2_X1 U757 ( .A1(G567), .A2(n822), .ZN(n677) );
  NAND2_X1 U758 ( .A1(n678), .A2(n677), .ZN(n824) );
  NAND2_X1 U759 ( .A1(G661), .A2(G483), .ZN(n679) );
  NOR2_X1 U760 ( .A1(n824), .A2(n679), .ZN(n821) );
  NAND2_X1 U761 ( .A1(n821), .A2(G36), .ZN(G176) );
  INV_X1 U762 ( .A(G301), .ZN(G171) );
  XOR2_X1 U763 ( .A(KEYINPUT32), .B(KEYINPUT105), .Z(n735) );
  AND2_X1 U764 ( .A1(G160), .A2(G1996), .ZN(n681) );
  NOR2_X1 U765 ( .A1(G164), .A2(G1384), .ZN(n769) );
  AND2_X1 U766 ( .A1(n769), .A2(G40), .ZN(n683) );
  XNOR2_X1 U767 ( .A(n682), .B(KEYINPUT26), .ZN(n685) );
  NAND2_X1 U768 ( .A1(G160), .A2(n683), .ZN(n688) );
  AND2_X1 U769 ( .A1(n688), .A2(G1341), .ZN(n684) );
  NOR2_X1 U770 ( .A1(n976), .A2(n687), .ZN(n686) );
  XNOR2_X1 U771 ( .A(n686), .B(KEYINPUT98), .ZN(n696) );
  NAND2_X1 U772 ( .A1(n687), .A2(n976), .ZN(n693) );
  BUF_X2 U773 ( .A(n688), .Z(n725) );
  NAND2_X1 U774 ( .A1(n709), .A2(G2067), .ZN(n690) );
  NAND2_X1 U775 ( .A1(G1348), .A2(n725), .ZN(n689) );
  NAND2_X1 U776 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U777 ( .A(n691), .B(KEYINPUT96), .ZN(n692) );
  NAND2_X1 U778 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U779 ( .A(n694), .B(KEYINPUT97), .ZN(n695) );
  OR2_X1 U780 ( .A1(n696), .A2(n695), .ZN(n701) );
  INV_X1 U781 ( .A(G2072), .ZN(n985) );
  NOR2_X1 U782 ( .A1(n725), .A2(n985), .ZN(n698) );
  XOR2_X1 U783 ( .A(KEYINPUT27), .B(KEYINPUT95), .Z(n697) );
  XNOR2_X1 U784 ( .A(n698), .B(n697), .ZN(n700) );
  NAND2_X1 U785 ( .A1(n725), .A2(G1956), .ZN(n699) );
  NAND2_X1 U786 ( .A1(n700), .A2(n699), .ZN(n703) );
  NAND2_X1 U787 ( .A1(n701), .A2(n509), .ZN(n702) );
  XNOR2_X1 U788 ( .A(n702), .B(KEYINPUT99), .ZN(n706) );
  NAND2_X1 U789 ( .A1(G299), .A2(n703), .ZN(n704) );
  XOR2_X1 U790 ( .A(KEYINPUT28), .B(n704), .Z(n705) );
  XNOR2_X1 U791 ( .A(n707), .B(KEYINPUT29), .ZN(n713) );
  XNOR2_X1 U792 ( .A(G2078), .B(KEYINPUT25), .ZN(n989) );
  NAND2_X1 U793 ( .A1(n709), .A2(n989), .ZN(n708) );
  XNOR2_X1 U794 ( .A(n708), .B(KEYINPUT94), .ZN(n711) );
  OR2_X1 U795 ( .A1(G1961), .A2(n709), .ZN(n710) );
  NAND2_X1 U796 ( .A1(n711), .A2(n710), .ZN(n717) );
  NAND2_X1 U797 ( .A1(G171), .A2(n717), .ZN(n712) );
  NAND2_X1 U798 ( .A1(n713), .A2(n712), .ZN(n723) );
  NAND2_X1 U799 ( .A1(G8), .A2(n725), .ZN(n764) );
  NOR2_X1 U800 ( .A1(G1966), .A2(n764), .ZN(n738) );
  NOR2_X1 U801 ( .A1(G2084), .A2(n725), .ZN(n737) );
  NOR2_X1 U802 ( .A1(n738), .A2(n737), .ZN(n714) );
  NAND2_X1 U803 ( .A1(G8), .A2(n714), .ZN(n715) );
  XNOR2_X1 U804 ( .A(KEYINPUT30), .B(n715), .ZN(n716) );
  NOR2_X1 U805 ( .A1(G168), .A2(n716), .ZN(n719) );
  NOR2_X1 U806 ( .A1(G171), .A2(n717), .ZN(n718) );
  NOR2_X1 U807 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U808 ( .A(n720), .B(KEYINPUT100), .Z(n721) );
  XNOR2_X1 U809 ( .A(KEYINPUT31), .B(n721), .ZN(n722) );
  NAND2_X1 U810 ( .A1(n723), .A2(n722), .ZN(n736) );
  NAND2_X1 U811 ( .A1(n736), .A2(G286), .ZN(n724) );
  XNOR2_X1 U812 ( .A(n724), .B(KEYINPUT102), .ZN(n732) );
  NOR2_X1 U813 ( .A1(G2090), .A2(n725), .ZN(n726) );
  XOR2_X1 U814 ( .A(KEYINPUT103), .B(n726), .Z(n728) );
  NOR2_X1 U815 ( .A1(G1971), .A2(n764), .ZN(n727) );
  NOR2_X1 U816 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U817 ( .A(n729), .B(KEYINPUT104), .ZN(n730) );
  NAND2_X1 U818 ( .A1(n730), .A2(G303), .ZN(n731) );
  NAND2_X1 U819 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U820 ( .A1(n733), .A2(G8), .ZN(n734) );
  XNOR2_X1 U821 ( .A(n735), .B(n734), .ZN(n757) );
  NOR2_X1 U822 ( .A1(n738), .A2(n511), .ZN(n739) );
  XNOR2_X1 U823 ( .A(n740), .B(KEYINPUT101), .ZN(n756) );
  NAND2_X1 U824 ( .A1(G288), .A2(G1976), .ZN(n741) );
  XNOR2_X1 U825 ( .A(n741), .B(KEYINPUT106), .ZN(n967) );
  INV_X1 U826 ( .A(n967), .ZN(n742) );
  OR2_X1 U827 ( .A1(n742), .A2(n764), .ZN(n746) );
  INV_X1 U828 ( .A(n746), .ZN(n743) );
  AND2_X1 U829 ( .A1(n756), .A2(n743), .ZN(n744) );
  AND2_X1 U830 ( .A1(n757), .A2(n744), .ZN(n750) );
  NOR2_X1 U831 ( .A1(G1976), .A2(G288), .ZN(n751) );
  NOR2_X1 U832 ( .A1(G1971), .A2(G303), .ZN(n745) );
  NOR2_X1 U833 ( .A1(n751), .A2(n745), .ZN(n966) );
  OR2_X1 U834 ( .A1(n746), .A2(n966), .ZN(n748) );
  INV_X1 U835 ( .A(KEYINPUT33), .ZN(n747) );
  NAND2_X1 U836 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U837 ( .A1(n750), .A2(n749), .ZN(n754) );
  NAND2_X1 U838 ( .A1(n751), .A2(KEYINPUT33), .ZN(n752) );
  NOR2_X1 U839 ( .A1(n752), .A2(n764), .ZN(n753) );
  NOR2_X1 U840 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U841 ( .A(G1981), .B(G305), .Z(n958) );
  NAND2_X1 U842 ( .A1(n755), .A2(n958), .ZN(n767) );
  NAND2_X1 U843 ( .A1(n757), .A2(n756), .ZN(n760) );
  NOR2_X1 U844 ( .A1(G2090), .A2(G303), .ZN(n758) );
  NAND2_X1 U845 ( .A1(G8), .A2(n758), .ZN(n759) );
  NAND2_X1 U846 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U847 ( .A1(G1981), .A2(G305), .ZN(n762) );
  XOR2_X1 U848 ( .A(n762), .B(KEYINPUT24), .Z(n763) );
  NOR2_X1 U849 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U850 ( .A(n513), .B(KEYINPUT107), .ZN(n803) );
  NAND2_X1 U851 ( .A1(G160), .A2(G40), .ZN(n768) );
  NOR2_X1 U852 ( .A1(n769), .A2(n768), .ZN(n813) );
  XNOR2_X1 U853 ( .A(G2067), .B(KEYINPUT37), .ZN(n770) );
  XNOR2_X1 U854 ( .A(n770), .B(KEYINPUT90), .ZN(n811) );
  NAND2_X1 U855 ( .A1(G104), .A2(n876), .ZN(n772) );
  NAND2_X1 U856 ( .A1(G140), .A2(n877), .ZN(n771) );
  NAND2_X1 U857 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U858 ( .A(n773), .B(KEYINPUT91), .ZN(n774) );
  XNOR2_X1 U859 ( .A(n774), .B(KEYINPUT34), .ZN(n780) );
  XNOR2_X1 U860 ( .A(KEYINPUT35), .B(KEYINPUT92), .ZN(n778) );
  NAND2_X1 U861 ( .A1(G116), .A2(n871), .ZN(n776) );
  NAND2_X1 U862 ( .A1(G128), .A2(n544), .ZN(n775) );
  NAND2_X1 U863 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U864 ( .A(n778), .B(n777), .ZN(n779) );
  NAND2_X1 U865 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U866 ( .A(KEYINPUT36), .B(n781), .Z(n866) );
  NOR2_X1 U867 ( .A1(n811), .A2(n866), .ZN(n951) );
  NAND2_X1 U868 ( .A1(n813), .A2(n951), .ZN(n809) );
  INV_X1 U869 ( .A(n809), .ZN(n799) );
  NAND2_X1 U870 ( .A1(G131), .A2(n877), .ZN(n783) );
  NAND2_X1 U871 ( .A1(G119), .A2(n544), .ZN(n782) );
  NAND2_X1 U872 ( .A1(n783), .A2(n782), .ZN(n787) );
  NAND2_X1 U873 ( .A1(G95), .A2(n876), .ZN(n785) );
  NAND2_X1 U874 ( .A1(G107), .A2(n871), .ZN(n784) );
  NAND2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n786) );
  OR2_X1 U876 ( .A1(n787), .A2(n786), .ZN(n883) );
  AND2_X1 U877 ( .A1(n883), .A2(G1991), .ZN(n796) );
  NAND2_X1 U878 ( .A1(G141), .A2(n877), .ZN(n789) );
  NAND2_X1 U879 ( .A1(G129), .A2(n544), .ZN(n788) );
  NAND2_X1 U880 ( .A1(n789), .A2(n788), .ZN(n792) );
  NAND2_X1 U881 ( .A1(n876), .A2(G105), .ZN(n790) );
  XOR2_X1 U882 ( .A(KEYINPUT38), .B(n790), .Z(n791) );
  NOR2_X1 U883 ( .A1(n792), .A2(n791), .ZN(n794) );
  NAND2_X1 U884 ( .A1(n871), .A2(G117), .ZN(n793) );
  NAND2_X1 U885 ( .A1(n794), .A2(n793), .ZN(n853) );
  AND2_X1 U886 ( .A1(G1996), .A2(n853), .ZN(n795) );
  NOR2_X1 U887 ( .A1(n796), .A2(n795), .ZN(n946) );
  INV_X1 U888 ( .A(n813), .ZN(n797) );
  NOR2_X1 U889 ( .A1(n946), .A2(n797), .ZN(n806) );
  XOR2_X1 U890 ( .A(KEYINPUT93), .B(n806), .Z(n798) );
  NOR2_X1 U891 ( .A1(n799), .A2(n798), .ZN(n801) );
  XNOR2_X1 U892 ( .A(G1986), .B(G290), .ZN(n963) );
  NAND2_X1 U893 ( .A1(n963), .A2(n813), .ZN(n800) );
  AND2_X1 U894 ( .A1(n801), .A2(n800), .ZN(n802) );
  NAND2_X1 U895 ( .A1(n803), .A2(n802), .ZN(n816) );
  NOR2_X1 U896 ( .A1(G1996), .A2(n853), .ZN(n939) );
  NOR2_X1 U897 ( .A1(G1991), .A2(n883), .ZN(n944) );
  NOR2_X1 U898 ( .A1(G1986), .A2(G290), .ZN(n804) );
  NOR2_X1 U899 ( .A1(n944), .A2(n804), .ZN(n805) );
  NOR2_X1 U900 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U901 ( .A1(n939), .A2(n807), .ZN(n808) );
  XNOR2_X1 U902 ( .A(n808), .B(KEYINPUT39), .ZN(n810) );
  NAND2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n812) );
  NAND2_X1 U904 ( .A1(n811), .A2(n866), .ZN(n949) );
  NAND2_X1 U905 ( .A1(n812), .A2(n949), .ZN(n814) );
  NAND2_X1 U906 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U907 ( .A1(n816), .A2(n815), .ZN(n818) );
  XNOR2_X1 U908 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n817) );
  XNOR2_X1 U909 ( .A(n818), .B(n817), .ZN(G329) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n907), .ZN(G217) );
  AND2_X1 U911 ( .A1(G15), .A2(G2), .ZN(n819) );
  NAND2_X1 U912 ( .A1(G661), .A2(n819), .ZN(G259) );
  NAND2_X1 U913 ( .A1(G3), .A2(G1), .ZN(n820) );
  NAND2_X1 U914 ( .A1(n821), .A2(n820), .ZN(G188) );
  XNOR2_X1 U915 ( .A(G96), .B(KEYINPUT109), .ZN(G221) );
  NOR2_X1 U916 ( .A1(n823), .A2(n822), .ZN(G325) );
  XOR2_X1 U917 ( .A(KEYINPUT110), .B(G325), .Z(G261) );
  INV_X1 U919 ( .A(G120), .ZN(G236) );
  INV_X1 U920 ( .A(G108), .ZN(G238) );
  INV_X1 U921 ( .A(G69), .ZN(G235) );
  INV_X1 U922 ( .A(n824), .ZN(G319) );
  XOR2_X1 U923 ( .A(KEYINPUT112), .B(G1976), .Z(n826) );
  INV_X1 U924 ( .A(G1971), .ZN(n968) );
  XOR2_X1 U925 ( .A(G1986), .B(n968), .Z(n825) );
  XNOR2_X1 U926 ( .A(n826), .B(n825), .ZN(n827) );
  XOR2_X1 U927 ( .A(n827), .B(KEYINPUT41), .Z(n830) );
  INV_X1 U928 ( .A(G1996), .ZN(n828) );
  XOR2_X1 U929 ( .A(n828), .B(G1991), .Z(n829) );
  XNOR2_X1 U930 ( .A(n830), .B(n829), .ZN(n834) );
  XOR2_X1 U931 ( .A(G1981), .B(G1956), .Z(n832) );
  XNOR2_X1 U932 ( .A(G1966), .B(G1961), .ZN(n831) );
  XNOR2_X1 U933 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U934 ( .A(n834), .B(n833), .Z(n836) );
  XNOR2_X1 U935 ( .A(G2474), .B(KEYINPUT113), .ZN(n835) );
  XNOR2_X1 U936 ( .A(n836), .B(n835), .ZN(G229) );
  XNOR2_X1 U937 ( .A(KEYINPUT111), .B(n985), .ZN(n838) );
  XNOR2_X1 U938 ( .A(G2084), .B(G2078), .ZN(n837) );
  XNOR2_X1 U939 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U940 ( .A(n839), .B(G2096), .Z(n841) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2090), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U943 ( .A(G2100), .B(KEYINPUT43), .Z(n843) );
  XNOR2_X1 U944 ( .A(G2678), .B(KEYINPUT42), .ZN(n842) );
  XNOR2_X1 U945 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U946 ( .A(n845), .B(n844), .Z(G227) );
  NAND2_X1 U947 ( .A1(n544), .A2(G124), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n846), .B(KEYINPUT44), .ZN(n848) );
  NAND2_X1 U949 ( .A1(n876), .A2(G100), .ZN(n847) );
  NAND2_X1 U950 ( .A1(n848), .A2(n847), .ZN(n852) );
  NAND2_X1 U951 ( .A1(G136), .A2(n877), .ZN(n850) );
  NAND2_X1 U952 ( .A1(G112), .A2(n871), .ZN(n849) );
  NAND2_X1 U953 ( .A1(n850), .A2(n849), .ZN(n851) );
  NOR2_X1 U954 ( .A1(n852), .A2(n851), .ZN(G162) );
  XOR2_X1 U955 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n855) );
  XOR2_X1 U956 ( .A(n853), .B(KEYINPUT117), .Z(n854) );
  XNOR2_X1 U957 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U958 ( .A(G160), .B(n856), .ZN(n870) );
  NAND2_X1 U959 ( .A1(G118), .A2(n871), .ZN(n858) );
  NAND2_X1 U960 ( .A1(G130), .A2(n544), .ZN(n857) );
  NAND2_X1 U961 ( .A1(n858), .A2(n857), .ZN(n864) );
  NAND2_X1 U962 ( .A1(n877), .A2(G142), .ZN(n859) );
  XNOR2_X1 U963 ( .A(n859), .B(KEYINPUT114), .ZN(n861) );
  NAND2_X1 U964 ( .A1(G106), .A2(n876), .ZN(n860) );
  NAND2_X1 U965 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U966 ( .A(KEYINPUT45), .B(n862), .Z(n863) );
  NOR2_X1 U967 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U968 ( .A(n943), .B(n865), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n866), .B(G162), .ZN(n867) );
  XNOR2_X1 U970 ( .A(n868), .B(n867), .ZN(n869) );
  XNOR2_X1 U971 ( .A(n870), .B(n869), .ZN(n886) );
  NAND2_X1 U972 ( .A1(G115), .A2(n871), .ZN(n873) );
  NAND2_X1 U973 ( .A1(G127), .A2(n544), .ZN(n872) );
  NAND2_X1 U974 ( .A1(n873), .A2(n872), .ZN(n875) );
  XOR2_X1 U975 ( .A(KEYINPUT47), .B(KEYINPUT116), .Z(n874) );
  XNOR2_X1 U976 ( .A(n875), .B(n874), .ZN(n882) );
  NAND2_X1 U977 ( .A1(G103), .A2(n876), .ZN(n879) );
  NAND2_X1 U978 ( .A1(G139), .A2(n877), .ZN(n878) );
  NAND2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U980 ( .A(KEYINPUT115), .B(n880), .Z(n881) );
  NOR2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n934) );
  XNOR2_X1 U982 ( .A(G164), .B(n934), .ZN(n884) );
  XNOR2_X1 U983 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U984 ( .A(n886), .B(n885), .Z(n887) );
  NOR2_X1 U985 ( .A1(G37), .A2(n887), .ZN(G395) );
  XOR2_X1 U986 ( .A(G301), .B(n976), .Z(n889) );
  XNOR2_X1 U987 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U988 ( .A(n890), .B(G286), .ZN(n891) );
  NOR2_X1 U989 ( .A1(G37), .A2(n891), .ZN(G397) );
  XOR2_X1 U990 ( .A(G2451), .B(G2430), .Z(n893) );
  XNOR2_X1 U991 ( .A(G2438), .B(G2443), .ZN(n892) );
  XNOR2_X1 U992 ( .A(n893), .B(n892), .ZN(n899) );
  XOR2_X1 U993 ( .A(G2435), .B(G2454), .Z(n895) );
  XNOR2_X1 U994 ( .A(G1341), .B(G1348), .ZN(n894) );
  XNOR2_X1 U995 ( .A(n895), .B(n894), .ZN(n897) );
  XOR2_X1 U996 ( .A(G2446), .B(G2427), .Z(n896) );
  XNOR2_X1 U997 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U998 ( .A(n899), .B(n898), .Z(n900) );
  NAND2_X1 U999 ( .A1(G14), .A2(n900), .ZN(n906) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n906), .ZN(n903) );
  NOR2_X1 U1001 ( .A1(G229), .A2(G227), .ZN(n901) );
  XNOR2_X1 U1002 ( .A(KEYINPUT49), .B(n901), .ZN(n902) );
  NOR2_X1 U1003 ( .A1(n903), .A2(n902), .ZN(n905) );
  NOR2_X1 U1004 ( .A1(G395), .A2(G397), .ZN(n904) );
  NAND2_X1 U1005 ( .A1(n905), .A2(n904), .ZN(G225) );
  INV_X1 U1006 ( .A(G225), .ZN(G308) );
  INV_X1 U1007 ( .A(n906), .ZN(G401) );
  INV_X1 U1008 ( .A(n907), .ZN(G223) );
  INV_X1 U1009 ( .A(G303), .ZN(G166) );
  XOR2_X1 U1010 ( .A(G16), .B(KEYINPUT124), .Z(n932) );
  XOR2_X1 U1011 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n930) );
  XNOR2_X1 U1012 ( .A(G5), .B(G1961), .ZN(n908) );
  XNOR2_X1 U1013 ( .A(n908), .B(KEYINPUT125), .ZN(n926) );
  XOR2_X1 U1014 ( .A(G1348), .B(KEYINPUT59), .Z(n909) );
  XNOR2_X1 U1015 ( .A(G4), .B(n909), .ZN(n911) );
  XNOR2_X1 U1016 ( .A(G20), .B(G1956), .ZN(n910) );
  NOR2_X1 U1017 ( .A1(n911), .A2(n910), .ZN(n915) );
  XNOR2_X1 U1018 ( .A(G1341), .B(G19), .ZN(n913) );
  XNOR2_X1 U1019 ( .A(G1981), .B(G6), .ZN(n912) );
  NOR2_X1 U1020 ( .A1(n913), .A2(n912), .ZN(n914) );
  NAND2_X1 U1021 ( .A1(n915), .A2(n914), .ZN(n916) );
  XNOR2_X1 U1022 ( .A(n916), .B(KEYINPUT60), .ZN(n924) );
  XOR2_X1 U1023 ( .A(G1986), .B(G24), .Z(n920) );
  XOR2_X1 U1024 ( .A(n968), .B(G22), .Z(n918) );
  XNOR2_X1 U1025 ( .A(G23), .B(G1976), .ZN(n917) );
  NOR2_X1 U1026 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1027 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1028 ( .A(n921), .B(KEYINPUT58), .ZN(n922) );
  XNOR2_X1 U1029 ( .A(KEYINPUT126), .B(n922), .ZN(n923) );
  NOR2_X1 U1030 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1031 ( .A1(n926), .A2(n925), .ZN(n928) );
  XNOR2_X1 U1032 ( .A(G21), .B(G1966), .ZN(n927) );
  NOR2_X1 U1033 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1034 ( .A(n930), .B(n929), .ZN(n931) );
  NAND2_X1 U1035 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1036 ( .A1(G11), .A2(n933), .ZN(n1011) );
  XOR2_X1 U1037 ( .A(G164), .B(G2078), .Z(n936) );
  XOR2_X1 U1038 ( .A(G2072), .B(n934), .Z(n935) );
  NOR2_X1 U1039 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1040 ( .A(KEYINPUT50), .B(n937), .Z(n942) );
  XOR2_X1 U1041 ( .A(G2090), .B(G162), .Z(n938) );
  NOR2_X1 U1042 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1043 ( .A(KEYINPUT51), .B(n940), .ZN(n941) );
  NOR2_X1 U1044 ( .A1(n942), .A2(n941), .ZN(n954) );
  NOR2_X1 U1045 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1046 ( .A1(n946), .A2(n945), .ZN(n948) );
  XOR2_X1 U1047 ( .A(G160), .B(G2084), .Z(n947) );
  NOR2_X1 U1048 ( .A1(n948), .A2(n947), .ZN(n950) );
  NAND2_X1 U1049 ( .A1(n950), .A2(n949), .ZN(n952) );
  NOR2_X1 U1050 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1052 ( .A(KEYINPUT118), .B(n955), .ZN(n956) );
  XNOR2_X1 U1053 ( .A(n956), .B(KEYINPUT52), .ZN(n957) );
  NAND2_X1 U1054 ( .A1(n957), .A2(G29), .ZN(n1009) );
  XOR2_X1 U1055 ( .A(G16), .B(KEYINPUT56), .Z(n984) );
  XNOR2_X1 U1056 ( .A(G168), .B(G1966), .ZN(n959) );
  NAND2_X1 U1057 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1058 ( .A(n960), .B(KEYINPUT57), .ZN(n975) );
  XNOR2_X1 U1059 ( .A(G1341), .B(n508), .ZN(n962) );
  NOR2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n965) );
  XOR2_X1 U1061 ( .A(G1956), .B(G299), .Z(n964) );
  NAND2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n973) );
  NAND2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n970) );
  NOR2_X1 U1064 ( .A1(G166), .A2(n968), .ZN(n969) );
  NOR2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1066 ( .A(KEYINPUT122), .B(n971), .Z(n972) );
  NOR2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n981) );
  XOR2_X1 U1069 ( .A(n976), .B(G1348), .Z(n978) );
  XNOR2_X1 U1070 ( .A(G301), .B(G1961), .ZN(n977) );
  NOR2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1072 ( .A(n979), .B(KEYINPUT121), .ZN(n980) );
  NOR2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1074 ( .A(KEYINPUT123), .B(n982), .Z(n983) );
  NOR2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n1007) );
  XNOR2_X1 U1076 ( .A(G2067), .B(G26), .ZN(n987) );
  XOR2_X1 U1077 ( .A(G33), .B(n985), .Z(n986) );
  NOR2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n995) );
  XOR2_X1 U1079 ( .A(G25), .B(G1991), .Z(n988) );
  NAND2_X1 U1080 ( .A1(n988), .A2(G28), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(n989), .B(G27), .ZN(n991) );
  XOR2_X1 U1082 ( .A(G1996), .B(G32), .Z(n990) );
  NAND2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(n996), .B(KEYINPUT53), .ZN(n999) );
  XOR2_X1 U1087 ( .A(G2084), .B(G34), .Z(n997) );
  XNOR2_X1 U1088 ( .A(KEYINPUT54), .B(n997), .ZN(n998) );
  NAND2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(G35), .B(G2090), .ZN(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(n1002), .B(KEYINPUT120), .ZN(n1003) );
  NOR2_X1 U1093 ( .A1(G29), .A2(n1003), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(KEYINPUT55), .B(n1004), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(KEYINPUT119), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1099 ( .A(KEYINPUT62), .B(n1012), .Z(G150) );
  INV_X1 U1100 ( .A(G150), .ZN(G311) );
endmodule

