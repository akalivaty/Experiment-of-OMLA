

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578;

  INV_X1 U319 ( .A(KEYINPUT102), .ZN(n410) );
  XNOR2_X1 U320 ( .A(n298), .B(n297), .ZN(n302) );
  XNOR2_X1 U321 ( .A(n443), .B(KEYINPUT38), .ZN(n497) );
  NOR2_X1 U322 ( .A1(n570), .A2(n457), .ZN(n458) );
  XNOR2_X1 U323 ( .A(KEYINPUT48), .B(KEYINPUT113), .ZN(n462) );
  XNOR2_X1 U324 ( .A(n463), .B(n462), .ZN(n522) );
  XNOR2_X1 U325 ( .A(n335), .B(G134GAT), .ZN(n336) );
  INV_X1 U326 ( .A(G176GAT), .ZN(n295) );
  XNOR2_X1 U327 ( .A(KEYINPUT54), .B(KEYINPUT125), .ZN(n465) );
  XNOR2_X1 U328 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U329 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U330 ( .A(n466), .B(n465), .ZN(n563) );
  XNOR2_X1 U331 ( .A(n410), .B(KEYINPUT37), .ZN(n411) );
  XNOR2_X1 U332 ( .A(n412), .B(n411), .ZN(n510) );
  INV_X1 U333 ( .A(G43GAT), .ZN(n444) );
  XNOR2_X1 U334 ( .A(n304), .B(n303), .ZN(n525) );
  XNOR2_X1 U335 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U336 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U337 ( .A(n475), .B(n474), .ZN(G1349GAT) );
  XNOR2_X1 U338 ( .A(n447), .B(n446), .ZN(G1330GAT) );
  XOR2_X1 U339 ( .A(G99GAT), .B(G190GAT), .Z(n288) );
  XNOR2_X1 U340 ( .A(G43GAT), .B(G113GAT), .ZN(n287) );
  XNOR2_X1 U341 ( .A(n288), .B(n287), .ZN(n292) );
  XOR2_X1 U342 ( .A(KEYINPUT66), .B(KEYINPUT20), .Z(n290) );
  XNOR2_X1 U343 ( .A(G169GAT), .B(G71GAT), .ZN(n289) );
  XNOR2_X1 U344 ( .A(n290), .B(n289), .ZN(n291) );
  XNOR2_X1 U345 ( .A(n292), .B(n291), .ZN(n304) );
  XOR2_X1 U346 ( .A(G15GAT), .B(G127GAT), .Z(n310) );
  XOR2_X1 U347 ( .A(G120GAT), .B(KEYINPUT83), .Z(n294) );
  XNOR2_X1 U348 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n293) );
  XNOR2_X1 U349 ( .A(n294), .B(n293), .ZN(n375) );
  XOR2_X1 U350 ( .A(n310), .B(n375), .Z(n298) );
  NAND2_X1 U351 ( .A1(G227GAT), .A2(G233GAT), .ZN(n296) );
  XOR2_X1 U352 ( .A(G183GAT), .B(KEYINPUT18), .Z(n300) );
  XNOR2_X1 U353 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n299) );
  XNOR2_X1 U354 ( .A(n300), .B(n299), .ZN(n394) );
  XNOR2_X1 U355 ( .A(n394), .B(KEYINPUT84), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U357 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n306) );
  XNOR2_X1 U358 ( .A(G8GAT), .B(G1GAT), .ZN(n305) );
  XNOR2_X1 U359 ( .A(n306), .B(n305), .ZN(n309) );
  XOR2_X1 U360 ( .A(G57GAT), .B(KEYINPUT72), .Z(n308) );
  XNOR2_X1 U361 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n431) );
  XOR2_X1 U363 ( .A(n309), .B(n431), .Z(n312) );
  XOR2_X1 U364 ( .A(G22GAT), .B(G155GAT), .Z(n358) );
  XNOR2_X1 U365 ( .A(n310), .B(n358), .ZN(n311) );
  XNOR2_X1 U366 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U367 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n314) );
  NAND2_X1 U368 ( .A1(G231GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U369 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U370 ( .A(n316), .B(n315), .Z(n321) );
  XOR2_X1 U371 ( .A(G64GAT), .B(G78GAT), .Z(n318) );
  XNOR2_X1 U372 ( .A(G183GAT), .B(G211GAT), .ZN(n317) );
  XNOR2_X1 U373 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U374 ( .A(n319), .B(KEYINPUT12), .ZN(n320) );
  XOR2_X1 U375 ( .A(n321), .B(n320), .Z(n476) );
  INV_X1 U376 ( .A(n476), .ZN(n573) );
  INV_X1 U377 ( .A(KEYINPUT71), .ZN(n325) );
  XOR2_X1 U378 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n323) );
  XNOR2_X1 U379 ( .A(G43GAT), .B(G29GAT), .ZN(n322) );
  XNOR2_X1 U380 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n325), .B(n324), .ZN(n427) );
  XOR2_X1 U382 ( .A(n427), .B(G106GAT), .Z(n332) );
  XOR2_X1 U383 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n327) );
  XNOR2_X1 U384 ( .A(KEYINPUT11), .B(KEYINPUT69), .ZN(n326) );
  XNOR2_X1 U385 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U386 ( .A(n328), .B(KEYINPUT9), .Z(n330) );
  XOR2_X1 U387 ( .A(G50GAT), .B(G162GAT), .Z(n359) );
  XNOR2_X1 U388 ( .A(G218GAT), .B(n359), .ZN(n329) );
  XOR2_X1 U389 ( .A(n330), .B(n329), .Z(n331) );
  XNOR2_X1 U390 ( .A(n332), .B(n331), .ZN(n340) );
  XOR2_X1 U391 ( .A(KEYINPUT10), .B(KEYINPUT79), .Z(n334) );
  XNOR2_X1 U392 ( .A(KEYINPUT65), .B(KEYINPUT78), .ZN(n333) );
  XNOR2_X1 U393 ( .A(n334), .B(n333), .ZN(n337) );
  AND2_X1 U394 ( .A1(G232GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n338), .B(G92GAT), .ZN(n339) );
  XNOR2_X1 U396 ( .A(n340), .B(n339), .ZN(n344) );
  XNOR2_X1 U397 ( .A(G36GAT), .B(G190GAT), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n341), .B(KEYINPUT80), .ZN(n386) );
  XNOR2_X1 U399 ( .A(G99GAT), .B(G85GAT), .ZN(n342) );
  XNOR2_X1 U400 ( .A(n342), .B(KEYINPUT76), .ZN(n439) );
  XNOR2_X1 U401 ( .A(n386), .B(n439), .ZN(n343) );
  XNOR2_X1 U402 ( .A(n344), .B(n343), .ZN(n558) );
  XNOR2_X1 U403 ( .A(n558), .B(KEYINPUT36), .ZN(n454) );
  XOR2_X1 U404 ( .A(G204GAT), .B(KEYINPUT22), .Z(n346) );
  XNOR2_X1 U405 ( .A(KEYINPUT87), .B(KEYINPUT24), .ZN(n345) );
  XNOR2_X1 U406 ( .A(n346), .B(n345), .ZN(n363) );
  XOR2_X1 U407 ( .A(KEYINPUT85), .B(KEYINPUT23), .Z(n348) );
  NAND2_X1 U408 ( .A1(G228GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U409 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U410 ( .A(n349), .B(KEYINPUT86), .Z(n354) );
  XOR2_X1 U411 ( .A(G211GAT), .B(KEYINPUT21), .Z(n351) );
  XNOR2_X1 U412 ( .A(G197GAT), .B(G218GAT), .ZN(n350) );
  XNOR2_X1 U413 ( .A(n351), .B(n350), .ZN(n390) );
  XNOR2_X1 U414 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n352) );
  XNOR2_X1 U415 ( .A(n352), .B(KEYINPUT2), .ZN(n372) );
  XNOR2_X1 U416 ( .A(n390), .B(n372), .ZN(n353) );
  XNOR2_X1 U417 ( .A(n354), .B(n353), .ZN(n357) );
  XOR2_X1 U418 ( .A(G78GAT), .B(G148GAT), .Z(n356) );
  XNOR2_X1 U419 ( .A(G106GAT), .B(KEYINPUT75), .ZN(n355) );
  XNOR2_X1 U420 ( .A(n356), .B(n355), .ZN(n440) );
  XOR2_X1 U421 ( .A(n357), .B(n440), .Z(n361) );
  XNOR2_X1 U422 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U423 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U424 ( .A(n363), .B(n362), .Z(n467) );
  XOR2_X1 U425 ( .A(n467), .B(KEYINPUT28), .Z(n519) );
  INV_X1 U426 ( .A(n519), .ZN(n528) );
  XOR2_X1 U427 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n365) );
  XNOR2_X1 U428 ( .A(KEYINPUT5), .B(KEYINPUT89), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n365), .B(n364), .ZN(n383) );
  XOR2_X1 U430 ( .A(G85GAT), .B(G148GAT), .Z(n367) );
  XNOR2_X1 U431 ( .A(G127GAT), .B(G155GAT), .ZN(n366) );
  XNOR2_X1 U432 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U433 ( .A(KEYINPUT90), .B(KEYINPUT88), .Z(n369) );
  XNOR2_X1 U434 ( .A(G57GAT), .B(KEYINPUT91), .ZN(n368) );
  XNOR2_X1 U435 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U436 ( .A(n371), .B(n370), .Z(n381) );
  XOR2_X1 U437 ( .A(n372), .B(KEYINPUT4), .Z(n374) );
  NAND2_X1 U438 ( .A1(G225GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U439 ( .A(n374), .B(n373), .ZN(n379) );
  XOR2_X1 U440 ( .A(G162GAT), .B(n375), .Z(n377) );
  XOR2_X1 U441 ( .A(G113GAT), .B(G1GAT), .Z(n413) );
  XNOR2_X1 U442 ( .A(G29GAT), .B(n413), .ZN(n376) );
  XNOR2_X1 U443 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U444 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U445 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U446 ( .A(n383), .B(n382), .ZN(n562) );
  XNOR2_X1 U447 ( .A(KEYINPUT27), .B(KEYINPUT93), .ZN(n395) );
  XOR2_X1 U448 ( .A(G169GAT), .B(G8GAT), .Z(n416) );
  XOR2_X1 U449 ( .A(KEYINPUT92), .B(n416), .Z(n385) );
  NAND2_X1 U450 ( .A1(G226GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U451 ( .A(n385), .B(n384), .ZN(n387) );
  XOR2_X1 U452 ( .A(n387), .B(n386), .Z(n392) );
  XOR2_X1 U453 ( .A(G64GAT), .B(G92GAT), .Z(n389) );
  XNOR2_X1 U454 ( .A(G176GAT), .B(G204GAT), .ZN(n388) );
  XNOR2_X1 U455 ( .A(n389), .B(n388), .ZN(n432) );
  XNOR2_X1 U456 ( .A(n390), .B(n432), .ZN(n391) );
  XNOR2_X1 U457 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U458 ( .A(n394), .B(n393), .Z(n514) );
  XOR2_X1 U459 ( .A(n395), .B(n514), .Z(n402) );
  NOR2_X1 U460 ( .A1(n562), .A2(n402), .ZN(n523) );
  NAND2_X1 U461 ( .A1(n525), .A2(n523), .ZN(n396) );
  NOR2_X1 U462 ( .A1(n528), .A2(n396), .ZN(n397) );
  XOR2_X1 U463 ( .A(KEYINPUT94), .B(n397), .Z(n408) );
  NOR2_X1 U464 ( .A1(n525), .A2(n514), .ZN(n398) );
  NOR2_X1 U465 ( .A1(n467), .A2(n398), .ZN(n399) );
  XOR2_X1 U466 ( .A(KEYINPUT25), .B(n399), .Z(n404) );
  XOR2_X1 U467 ( .A(KEYINPUT26), .B(KEYINPUT95), .Z(n401) );
  NAND2_X1 U468 ( .A1(n467), .A2(n525), .ZN(n400) );
  XNOR2_X1 U469 ( .A(n401), .B(n400), .ZN(n565) );
  NOR2_X1 U470 ( .A1(n565), .A2(n402), .ZN(n403) );
  NOR2_X1 U471 ( .A1(n404), .A2(n403), .ZN(n405) );
  XOR2_X1 U472 ( .A(KEYINPUT96), .B(n405), .Z(n406) );
  NAND2_X1 U473 ( .A1(n406), .A2(n562), .ZN(n407) );
  NAND2_X1 U474 ( .A1(n408), .A2(n407), .ZN(n478) );
  NAND2_X1 U475 ( .A1(n454), .A2(n478), .ZN(n409) );
  NOR2_X1 U476 ( .A1(n573), .A2(n409), .ZN(n412) );
  XOR2_X1 U477 ( .A(n413), .B(KEYINPUT29), .Z(n415) );
  NAND2_X1 U478 ( .A1(G229GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U479 ( .A(n415), .B(n414), .ZN(n417) );
  XOR2_X1 U480 ( .A(n417), .B(n416), .Z(n425) );
  XOR2_X1 U481 ( .A(G22GAT), .B(G197GAT), .Z(n419) );
  XNOR2_X1 U482 ( .A(G36GAT), .B(G50GAT), .ZN(n418) );
  XNOR2_X1 U483 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U484 ( .A(KEYINPUT70), .B(KEYINPUT30), .Z(n421) );
  XNOR2_X1 U485 ( .A(G141GAT), .B(G15GAT), .ZN(n420) );
  XNOR2_X1 U486 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U487 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U488 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U489 ( .A(n427), .B(n426), .Z(n499) );
  XOR2_X1 U490 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n429) );
  NAND2_X1 U491 ( .A1(G230GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U492 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U493 ( .A(n430), .B(KEYINPUT32), .Z(n434) );
  XNOR2_X1 U494 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U495 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U496 ( .A(KEYINPUT74), .B(KEYINPUT77), .Z(n436) );
  XNOR2_X1 U497 ( .A(G120GAT), .B(KEYINPUT73), .ZN(n435) );
  XNOR2_X1 U498 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U499 ( .A(n438), .B(n437), .Z(n442) );
  XNOR2_X1 U500 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U501 ( .A(n442), .B(n441), .ZN(n570) );
  NOR2_X1 U502 ( .A1(n499), .A2(n570), .ZN(n480) );
  NAND2_X1 U503 ( .A1(n510), .A2(n480), .ZN(n443) );
  NOR2_X1 U504 ( .A1(n525), .A2(n497), .ZN(n447) );
  XNOR2_X1 U505 ( .A(KEYINPUT40), .B(KEYINPUT104), .ZN(n445) );
  INV_X1 U506 ( .A(n514), .ZN(n464) );
  XOR2_X1 U507 ( .A(KEYINPUT64), .B(KEYINPUT41), .Z(n448) );
  XNOR2_X1 U508 ( .A(n570), .B(n448), .ZN(n546) );
  INV_X1 U509 ( .A(n499), .ZN(n566) );
  NAND2_X1 U510 ( .A1(n546), .A2(n566), .ZN(n449) );
  XNOR2_X1 U511 ( .A(n449), .B(KEYINPUT110), .ZN(n450) );
  XNOR2_X1 U512 ( .A(KEYINPUT46), .B(n450), .ZN(n452) );
  NOR2_X1 U513 ( .A1(n558), .A2(n573), .ZN(n451) );
  NAND2_X1 U514 ( .A1(n452), .A2(n451), .ZN(n453) );
  XNOR2_X1 U515 ( .A(n453), .B(KEYINPUT47), .ZN(n461) );
  NAND2_X1 U516 ( .A1(n454), .A2(n573), .ZN(n456) );
  XOR2_X1 U517 ( .A(KEYINPUT45), .B(KEYINPUT111), .Z(n455) );
  XNOR2_X1 U518 ( .A(n456), .B(n455), .ZN(n457) );
  XOR2_X1 U519 ( .A(KEYINPUT112), .B(n458), .Z(n459) );
  NOR2_X1 U520 ( .A1(n566), .A2(n459), .ZN(n460) );
  NOR2_X1 U521 ( .A1(n461), .A2(n460), .ZN(n463) );
  NAND2_X1 U522 ( .A1(n464), .A2(n522), .ZN(n466) );
  INV_X1 U523 ( .A(n467), .ZN(n468) );
  AND2_X1 U524 ( .A1(n562), .A2(n468), .ZN(n469) );
  AND2_X1 U525 ( .A1(n563), .A2(n469), .ZN(n470) );
  XNOR2_X1 U526 ( .A(n470), .B(KEYINPUT55), .ZN(n471) );
  NOR2_X1 U527 ( .A1(n525), .A2(n471), .ZN(n559) );
  XOR2_X1 U528 ( .A(KEYINPUT105), .B(n546), .Z(n531) );
  NAND2_X1 U529 ( .A1(n559), .A2(n531), .ZN(n475) );
  XOR2_X1 U530 ( .A(G176GAT), .B(KEYINPUT56), .Z(n473) );
  XNOR2_X1 U531 ( .A(KEYINPUT126), .B(KEYINPUT57), .ZN(n472) );
  NOR2_X1 U532 ( .A1(n558), .A2(n476), .ZN(n477) );
  XNOR2_X1 U533 ( .A(KEYINPUT16), .B(n477), .ZN(n479) );
  AND2_X1 U534 ( .A1(n479), .A2(n478), .ZN(n500) );
  NAND2_X1 U535 ( .A1(n480), .A2(n500), .ZN(n491) );
  NOR2_X1 U536 ( .A1(n562), .A2(n491), .ZN(n485) );
  XOR2_X1 U537 ( .A(KEYINPUT34), .B(KEYINPUT99), .Z(n482) );
  XNOR2_X1 U538 ( .A(G1GAT), .B(KEYINPUT98), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U540 ( .A(KEYINPUT97), .B(n483), .ZN(n484) );
  XNOR2_X1 U541 ( .A(n485), .B(n484), .ZN(G1324GAT) );
  NOR2_X1 U542 ( .A1(n514), .A2(n491), .ZN(n486) );
  XOR2_X1 U543 ( .A(KEYINPUT100), .B(n486), .Z(n487) );
  XNOR2_X1 U544 ( .A(G8GAT), .B(n487), .ZN(G1325GAT) );
  NOR2_X1 U545 ( .A1(n525), .A2(n491), .ZN(n489) );
  XNOR2_X1 U546 ( .A(KEYINPUT101), .B(KEYINPUT35), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U548 ( .A(G15GAT), .B(n490), .Z(G1326GAT) );
  NOR2_X1 U549 ( .A1(n519), .A2(n491), .ZN(n492) );
  XOR2_X1 U550 ( .A(G22GAT), .B(n492), .Z(G1327GAT) );
  NOR2_X1 U551 ( .A1(n497), .A2(n562), .ZN(n494) );
  XNOR2_X1 U552 ( .A(KEYINPUT39), .B(KEYINPUT103), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U554 ( .A(G29GAT), .B(n495), .Z(G1328GAT) );
  NOR2_X1 U555 ( .A1(n514), .A2(n497), .ZN(n496) );
  XOR2_X1 U556 ( .A(G36GAT), .B(n496), .Z(G1329GAT) );
  NOR2_X1 U557 ( .A1(n519), .A2(n497), .ZN(n498) );
  XOR2_X1 U558 ( .A(G50GAT), .B(n498), .Z(G1331GAT) );
  AND2_X1 U559 ( .A1(n531), .A2(n499), .ZN(n511) );
  NAND2_X1 U560 ( .A1(n511), .A2(n500), .ZN(n507) );
  NOR2_X1 U561 ( .A1(n562), .A2(n507), .ZN(n502) );
  XNOR2_X1 U562 ( .A(KEYINPUT42), .B(KEYINPUT106), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U564 ( .A(G57GAT), .B(n503), .Z(G1332GAT) );
  NOR2_X1 U565 ( .A1(n514), .A2(n507), .ZN(n504) );
  XOR2_X1 U566 ( .A(G64GAT), .B(n504), .Z(G1333GAT) );
  NOR2_X1 U567 ( .A1(n525), .A2(n507), .ZN(n506) );
  XNOR2_X1 U568 ( .A(G71GAT), .B(KEYINPUT107), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n506), .B(n505), .ZN(G1334GAT) );
  NOR2_X1 U570 ( .A1(n519), .A2(n507), .ZN(n509) );
  XNOR2_X1 U571 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(G1335GAT) );
  NAND2_X1 U573 ( .A1(n511), .A2(n510), .ZN(n518) );
  NOR2_X1 U574 ( .A1(n562), .A2(n518), .ZN(n512) );
  XOR2_X1 U575 ( .A(KEYINPUT108), .B(n512), .Z(n513) );
  XNOR2_X1 U576 ( .A(G85GAT), .B(n513), .ZN(G1336GAT) );
  NOR2_X1 U577 ( .A1(n514), .A2(n518), .ZN(n516) );
  XNOR2_X1 U578 ( .A(G92GAT), .B(KEYINPUT109), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n516), .B(n515), .ZN(G1337GAT) );
  NOR2_X1 U580 ( .A1(n525), .A2(n518), .ZN(n517) );
  XOR2_X1 U581 ( .A(G99GAT), .B(n517), .Z(G1338GAT) );
  NOR2_X1 U582 ( .A1(n519), .A2(n518), .ZN(n520) );
  XOR2_X1 U583 ( .A(KEYINPUT44), .B(n520), .Z(n521) );
  XNOR2_X1 U584 ( .A(G106GAT), .B(n521), .ZN(G1339GAT) );
  NAND2_X1 U585 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U586 ( .A(n524), .B(KEYINPUT114), .ZN(n541) );
  NOR2_X1 U587 ( .A1(n525), .A2(n541), .ZN(n526) );
  XNOR2_X1 U588 ( .A(n526), .B(KEYINPUT115), .ZN(n527) );
  NOR2_X1 U589 ( .A1(n528), .A2(n527), .ZN(n538) );
  NAND2_X1 U590 ( .A1(n566), .A2(n538), .ZN(n529) );
  XNOR2_X1 U591 ( .A(n529), .B(KEYINPUT116), .ZN(n530) );
  XNOR2_X1 U592 ( .A(G113GAT), .B(n530), .ZN(G1340GAT) );
  XNOR2_X1 U593 ( .A(KEYINPUT117), .B(KEYINPUT49), .ZN(n533) );
  AND2_X1 U594 ( .A1(n538), .A2(n531), .ZN(n532) );
  XNOR2_X1 U595 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U596 ( .A(G120GAT), .B(n534), .Z(G1341GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n536) );
  NAND2_X1 U598 ( .A1(n538), .A2(n573), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U600 ( .A(G127GAT), .B(n537), .Z(G1342GAT) );
  XOR2_X1 U601 ( .A(G134GAT), .B(KEYINPUT51), .Z(n540) );
  NAND2_X1 U602 ( .A1(n538), .A2(n558), .ZN(n539) );
  XNOR2_X1 U603 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n544) );
  NOR2_X1 U605 ( .A1(n541), .A2(n565), .ZN(n542) );
  XOR2_X1 U606 ( .A(KEYINPUT119), .B(n542), .Z(n553) );
  NAND2_X1 U607 ( .A1(n553), .A2(n566), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U609 ( .A(G141GAT), .B(n545), .ZN(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n548) );
  NAND2_X1 U611 ( .A1(n553), .A2(n546), .ZN(n547) );
  XNOR2_X1 U612 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(n549), .ZN(G1345GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n551) );
  NAND2_X1 U615 ( .A1(n553), .A2(n573), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U617 ( .A(G155GAT), .B(n552), .ZN(G1346GAT) );
  NAND2_X1 U618 ( .A1(n553), .A2(n558), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n554), .B(KEYINPUT124), .ZN(n555) );
  XNOR2_X1 U620 ( .A(G162GAT), .B(n555), .ZN(G1347GAT) );
  NAND2_X1 U621 ( .A1(n559), .A2(n566), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U623 ( .A1(n559), .A2(n573), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(KEYINPUT58), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n568) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n575) );
  NAND2_X1 U631 ( .A1(n575), .A2(n566), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U634 ( .A(G204GAT), .B(KEYINPUT61), .Z(n572) );
  NAND2_X1 U635 ( .A1(n575), .A2(n570), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n572), .B(n571), .ZN(G1353GAT) );
  NAND2_X1 U637 ( .A1(n575), .A2(n573), .ZN(n574) );
  XNOR2_X1 U638 ( .A(n574), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n577) );
  NAND2_X1 U640 ( .A1(n575), .A2(n454), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U642 ( .A(G218GAT), .B(n578), .ZN(G1355GAT) );
endmodule

