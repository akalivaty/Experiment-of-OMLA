//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n995,
    new_n996, new_n997;
  INV_X1    g000(.A(G36gat), .ZN(new_n202));
  AND2_X1   g001(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n206), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n208), .A2(KEYINPUT15), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(KEYINPUT15), .ZN(new_n210));
  XNOR2_X1  g009(.A(G43gat), .B(G50gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(new_n210), .B2(new_n211), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n213), .B(KEYINPUT17), .ZN(new_n214));
  INV_X1    g013(.A(G8gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(G15gat), .B(G22gat), .ZN(new_n216));
  OR2_X1    g015(.A1(new_n216), .A2(G1gat), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n215), .B1(new_n217), .B2(KEYINPUT91), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n216), .B1(new_n219), .B2(G1gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n218), .B(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n214), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n213), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G229gat), .A2(G233gat), .ZN(new_n227));
  XOR2_X1   g026(.A(new_n227), .B(KEYINPUT92), .Z(new_n228));
  NAND3_X1  g027(.A1(new_n226), .A2(KEYINPUT18), .A3(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n224), .A2(new_n228), .A3(new_n225), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT18), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n222), .B(new_n213), .ZN(new_n233));
  XOR2_X1   g032(.A(new_n228), .B(KEYINPUT13), .Z(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT93), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n233), .A2(KEYINPUT93), .A3(new_n234), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n229), .A2(new_n232), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(G113gat), .B(G141gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(G169gat), .B(G197gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g042(.A(KEYINPUT90), .B(KEYINPUT11), .Z(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT12), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n240), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n229), .A2(new_n232), .A3(new_n239), .A4(new_n246), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  XOR2_X1   g050(.A(KEYINPUT72), .B(KEYINPUT33), .Z(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT26), .ZN(new_n254));
  INV_X1    g053(.A(G169gat), .ZN(new_n255));
  INV_X1    g054(.A(G176gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n257), .B(new_n258), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(G183gat), .A2(G190gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT27), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G183gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT68), .ZN(new_n268));
  INV_X1    g067(.A(G190gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G183gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT27), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT68), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n265), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n267), .A2(new_n272), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n275), .A2(KEYINPUT28), .A3(new_n269), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n264), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(KEYINPUT65), .B(KEYINPUT25), .Z(new_n278));
  NOR2_X1   g077(.A1(new_n263), .A2(KEYINPUT24), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n271), .A2(G190gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n269), .A2(G183gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n279), .B1(new_n282), .B2(KEYINPUT24), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT23), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(new_n255), .A3(new_n256), .ZN(new_n286));
  NAND2_X1  g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT66), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n284), .A2(new_n286), .B1(new_n289), .B2(new_n259), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n283), .B1(new_n290), .B2(KEYINPUT67), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n286), .A2(new_n284), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n289), .A2(new_n259), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n292), .A2(new_n293), .A3(KEYINPUT67), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n278), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  AND3_X1   g094(.A1(new_n283), .A2(KEYINPUT25), .A3(new_n290), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n277), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G113gat), .ZN(new_n299));
  INV_X1    g098(.A(G120gat), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT1), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G127gat), .B(G134gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT70), .B(G113gat), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n301), .B(new_n302), .C1(new_n303), .C2(new_n300), .ZN(new_n304));
  NAND2_X1  g103(.A1(G113gat), .A2(G120gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G134gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G127gat), .ZN(new_n308));
  INV_X1    g107(.A(G127gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(G134gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n304), .A2(new_n312), .A3(KEYINPUT71), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT71), .B1(new_n304), .B2(new_n312), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n315), .ZN(new_n316));
  OR2_X1    g115(.A1(new_n313), .A2(new_n314), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n292), .A2(new_n293), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT67), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n290), .A2(KEYINPUT67), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(new_n321), .A3(new_n283), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n296), .B1(new_n322), .B2(new_n278), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n317), .B1(new_n323), .B2(new_n277), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n316), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G227gat), .A2(G233gat), .ZN(new_n326));
  XOR2_X1   g125(.A(new_n326), .B(KEYINPUT64), .Z(new_n327));
  AOI21_X1  g126(.A(new_n253), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(G15gat), .B(G43gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(G71gat), .B(G99gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT34), .B1(new_n325), .B2(new_n327), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT34), .ZN(new_n334));
  INV_X1    g133(.A(new_n327), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n316), .A2(new_n324), .A3(new_n334), .A4(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n333), .B(new_n336), .C1(new_n328), .C2(new_n331), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n327), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT32), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n342), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n338), .A2(new_n344), .A3(new_n339), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(G78gat), .B(G106gat), .Z(new_n347));
  XNOR2_X1  g146(.A(new_n347), .B(G50gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(KEYINPUT82), .ZN(new_n349));
  XOR2_X1   g148(.A(new_n349), .B(KEYINPUT31), .Z(new_n350));
  INV_X1    g149(.A(G155gat), .ZN(new_n351));
  INV_X1    g150(.A(G162gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(G155gat), .A2(G162gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(KEYINPUT2), .ZN(new_n357));
  XNOR2_X1  g156(.A(G141gat), .B(G148gat), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n357), .B1(new_n358), .B2(KEYINPUT77), .ZN(new_n359));
  INV_X1    g158(.A(G141gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(G148gat), .ZN(new_n361));
  INV_X1    g160(.A(G148gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(G141gat), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n361), .A2(new_n363), .A3(KEYINPUT77), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n356), .B1(new_n359), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n367), .B1(new_n362), .B2(G141gat), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n360), .A2(KEYINPUT78), .A3(G148gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(new_n363), .A3(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n354), .B1(new_n353), .B2(KEYINPUT2), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n366), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT3), .ZN(new_n374));
  XOR2_X1   g173(.A(G211gat), .B(G218gat), .Z(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(G211gat), .A2(G218gat), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT22), .ZN(new_n378));
  OR2_X1    g177(.A1(G197gat), .A2(G204gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(G197gat), .A2(G204gat), .ZN(new_n380));
  AOI221_X4 g179(.A(KEYINPUT74), .B1(new_n377), .B2(new_n378), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT74), .ZN(new_n382));
  XNOR2_X1  g181(.A(G197gat), .B(G204gat), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n382), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n376), .B1(new_n381), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n383), .A2(new_n382), .A3(new_n385), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n375), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT29), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT83), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n374), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT29), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n383), .A2(new_n385), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT74), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n375), .B1(new_n395), .B2(new_n388), .ZN(new_n396));
  INV_X1    g195(.A(new_n389), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n391), .B(new_n393), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n373), .B1(new_n392), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n366), .A2(new_n374), .A3(new_n372), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n393), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT84), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n389), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT84), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n401), .A2(new_n406), .A3(new_n393), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n403), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(G228gat), .ZN(new_n409));
  INV_X1    g208(.A(G233gat), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n400), .A2(new_n408), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(G22gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n361), .A2(new_n363), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT77), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n416), .A2(new_n364), .A3(new_n357), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n417), .A2(new_n356), .B1(new_n370), .B2(new_n371), .ZN(new_n418));
  INV_X1    g217(.A(new_n390), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n418), .B1(new_n419), .B2(new_n374), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n404), .B1(new_n393), .B2(new_n401), .ZN(new_n421));
  OAI22_X1  g220(.A1(new_n420), .A2(new_n421), .B1(new_n409), .B2(new_n410), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n412), .A2(new_n413), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n413), .B1(new_n412), .B2(new_n422), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT85), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n350), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT86), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n428), .B1(new_n425), .B2(new_n426), .ZN(new_n429));
  NOR4_X1   g228(.A1(new_n423), .A2(new_n424), .A3(KEYINPUT85), .A4(KEYINPUT86), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n427), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n350), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n412), .A2(new_n422), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(G22gat), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n412), .A2(new_n413), .A3(new_n422), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n432), .B1(new_n436), .B2(KEYINPUT85), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n425), .A2(new_n426), .A3(new_n428), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n434), .A2(new_n426), .A3(new_n435), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT86), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n437), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n346), .B1(new_n431), .B2(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(G8gat), .B(G36gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(G64gat), .B(G92gat), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n443), .B(new_n444), .Z(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT75), .ZN(new_n447));
  NAND2_X1  g246(.A1(G226gat), .A2(G233gat), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n448), .B1(new_n298), .B2(KEYINPUT29), .ZN(new_n449));
  OAI211_X1 g248(.A(G226gat), .B(G233gat), .C1(new_n323), .C2(new_n277), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n393), .B1(new_n323), .B2(new_n277), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT75), .B1(new_n452), .B2(new_n448), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n451), .A2(new_n405), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n404), .B1(new_n449), .B2(new_n450), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n446), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n449), .A2(new_n447), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n295), .A2(new_n297), .ZN(new_n458));
  INV_X1    g257(.A(new_n277), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n448), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n460), .B1(new_n448), .B2(new_n452), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n404), .B(new_n457), .C1(new_n461), .C2(new_n447), .ZN(new_n462));
  INV_X1    g261(.A(new_n455), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n462), .A2(KEYINPUT30), .A3(new_n463), .A4(new_n445), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n456), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n462), .A2(new_n463), .A3(new_n445), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT76), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT30), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n467), .B1(new_n466), .B2(new_n468), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n465), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n442), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT5), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT1), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n475), .B1(G113gat), .B2(G120gat), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n311), .A2(new_n476), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n299), .A2(KEYINPUT70), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n299), .A2(KEYINPUT70), .ZN(new_n479));
  OAI21_X1  g278(.A(G120gat), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI22_X1  g279(.A1(new_n477), .A2(new_n480), .B1(new_n306), .B2(new_n311), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT79), .B1(new_n418), .B2(new_n481), .ZN(new_n482));
  AND4_X1   g281(.A1(KEYINPUT79), .A2(new_n366), .A3(new_n481), .A4(new_n372), .ZN(new_n483));
  OAI22_X1  g282(.A1(new_n482), .A2(new_n483), .B1(new_n418), .B2(new_n481), .ZN(new_n484));
  NAND2_X1  g283(.A1(G225gat), .A2(G233gat), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n474), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT4), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n488), .B1(new_n482), .B2(new_n483), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n481), .B1(new_n373), .B2(KEYINPUT3), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n486), .B1(new_n490), .B2(new_n401), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n315), .A2(KEYINPUT4), .A3(new_n418), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n489), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT4), .B1(new_n315), .B2(new_n418), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n482), .A2(new_n483), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n494), .B1(new_n495), .B2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT2), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n497), .B1(G155gat), .B2(G162gat), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n498), .B1(new_n414), .B2(new_n415), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n355), .B1(new_n499), .B2(new_n364), .ZN(new_n500));
  INV_X1    g299(.A(new_n372), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT3), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n304), .A2(new_n312), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(new_n503), .A3(new_n401), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n504), .A2(new_n474), .A3(new_n485), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n487), .A2(new_n493), .B1(new_n496), .B2(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(G1gat), .B(G29gat), .Z(new_n507));
  XNOR2_X1  g306(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G57gat), .B(G85gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT88), .B1(new_n513), .B2(KEYINPUT6), .ZN(new_n514));
  INV_X1    g313(.A(new_n494), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT79), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(new_n373), .B2(new_n503), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n418), .A2(KEYINPUT79), .A3(new_n481), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n517), .A2(KEYINPUT4), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n505), .A2(new_n515), .A3(new_n519), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n489), .A2(new_n491), .A3(new_n492), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n517), .A2(new_n518), .B1(new_n373), .B2(new_n503), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT5), .B1(new_n522), .B2(new_n485), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n520), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n524), .A2(KEYINPUT6), .A3(new_n511), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT6), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n526), .B1(new_n506), .B2(new_n512), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n512), .B(new_n520), .C1(new_n521), .C2(new_n523), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n525), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n514), .B1(new_n530), .B2(KEYINPUT88), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n531), .A2(KEYINPUT35), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n473), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT81), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n469), .A2(new_n470), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n530), .A2(new_n456), .A3(new_n464), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n456), .A2(new_n464), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n511), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n540), .A2(new_n526), .A3(new_n528), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n539), .B1(new_n525), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n466), .A2(new_n468), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT76), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n542), .A2(new_n546), .A3(KEYINPUT81), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n442), .A2(new_n538), .A3(new_n547), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n548), .A2(KEYINPUT89), .A3(KEYINPUT35), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT89), .B1(new_n548), .B2(KEYINPUT35), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n534), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n496), .A2(new_n504), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n486), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT39), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n554), .B1(new_n522), .B2(new_n485), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n552), .A2(new_n554), .A3(new_n486), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n512), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT40), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n556), .A2(KEYINPUT40), .A3(new_n512), .A4(new_n557), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n561), .A2(new_n540), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n471), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n431), .A2(new_n441), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n449), .A2(new_n450), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n453), .B1(new_n565), .B2(KEYINPUT75), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(new_n405), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT37), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n568), .B1(new_n565), .B2(new_n404), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT38), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT87), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n455), .B1(new_n566), .B2(new_n404), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n571), .B1(new_n572), .B2(new_n568), .ZN(new_n573));
  NOR4_X1   g372(.A1(new_n454), .A2(KEYINPUT87), .A3(KEYINPUT37), .A4(new_n455), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n446), .B(new_n570), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n575), .A2(new_n531), .A3(new_n466), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT38), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n462), .A2(new_n463), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT87), .B1(new_n578), .B2(KEYINPUT37), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n572), .A2(new_n571), .A3(new_n568), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n445), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(KEYINPUT37), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n577), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n563), .B(new_n564), .C1(new_n576), .C2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n346), .A2(KEYINPUT73), .A3(KEYINPUT36), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT36), .B1(new_n346), .B2(KEYINPUT73), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n564), .B1(new_n538), .B2(new_n547), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n251), .B1(new_n551), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G85gat), .A2(G92gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT7), .ZN(new_n595));
  NAND2_X1  g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  INV_X1    g395(.A(G85gat), .ZN(new_n597));
  INV_X1    g396(.A(G92gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(KEYINPUT8), .A2(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G99gat), .B(G106gat), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n600), .B(new_n601), .Z(new_n602));
  NAND2_X1  g401(.A1(new_n214), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n602), .ZN(new_n604));
  AND2_X1   g403(.A1(G232gat), .A2(G233gat), .ZN(new_n605));
  AOI22_X1  g404(.A1(new_n604), .A2(new_n213), .B1(KEYINPUT41), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G190gat), .B(G218gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(G134gat), .B(G162gat), .Z(new_n610));
  NOR2_X1   g409(.A1(new_n605), .A2(KEYINPUT41), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT97), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT97), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n615), .B1(new_n617), .B2(new_n609), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  AND2_X1   g418(.A1(G71gat), .A2(G78gat), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n620), .A2(KEYINPUT9), .ZN(new_n621));
  XNOR2_X1  g420(.A(G57gat), .B(G64gat), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(G71gat), .A2(G78gat), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n620), .A2(KEYINPUT94), .ZN(new_n626));
  OR3_X1    g425(.A1(new_n623), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n625), .B1(new_n623), .B2(new_n626), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n629), .B(KEYINPUT96), .Z(new_n630));
  AOI21_X1  g429(.A(new_n222), .B1(new_n630), .B2(KEYINPUT21), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n629), .A2(KEYINPUT21), .ZN(new_n632));
  XNOR2_X1  g431(.A(G127gat), .B(G155gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n631), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(G231gat), .A2(G233gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT95), .ZN(new_n637));
  XOR2_X1   g436(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G183gat), .B(G211gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n635), .B(new_n641), .Z(new_n642));
  NAND2_X1  g441(.A1(new_n619), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n630), .A2(KEYINPUT10), .A3(new_n604), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n602), .B(new_n629), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT10), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n645), .A2(KEYINPUT98), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT98), .B1(new_n645), .B2(new_n646), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n644), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(G230gat), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n650), .A2(new_n410), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n653), .B1(new_n652), .B2(new_n645), .ZN(new_n654));
  XNOR2_X1  g453(.A(G120gat), .B(G148gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n654), .A2(new_n658), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n643), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n593), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT99), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n593), .A2(KEYINPUT99), .A3(new_n662), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n530), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g469(.A(KEYINPUT16), .B(G8gat), .Z(new_n671));
  AND3_X1   g470(.A1(new_n667), .A2(new_n471), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n215), .B1(new_n667), .B2(new_n471), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT42), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(KEYINPUT42), .B2(new_n672), .ZN(G1325gat));
  INV_X1    g474(.A(G15gat), .ZN(new_n676));
  INV_X1    g475(.A(new_n346), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n667), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n588), .B1(new_n665), .B2(new_n666), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n678), .B1(new_n679), .B2(new_n676), .ZN(G1326gat));
  INV_X1    g479(.A(new_n564), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n667), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT43), .B(G22gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1327gat));
  INV_X1    g483(.A(KEYINPUT101), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n250), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n248), .A2(KEYINPUT101), .A3(new_n249), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n688), .A2(new_n642), .A3(new_n661), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n619), .A2(KEYINPUT44), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n584), .B(new_n588), .C1(new_n590), .C2(KEYINPUT102), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n590), .A2(KEYINPUT102), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n694), .B1(new_n551), .B2(KEYINPUT103), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT103), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n696), .B(new_n534), .C1(new_n549), .C2(new_n550), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n691), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n551), .A2(new_n592), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n699), .B1(new_n700), .B2(new_n618), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n668), .B(new_n689), .C1(new_n698), .C2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(KEYINPUT104), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n692), .A2(new_n693), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n538), .A2(new_n547), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n437), .A2(new_n440), .A3(new_n438), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n437), .B1(new_n440), .B2(new_n438), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n677), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT35), .B1(new_n705), .B2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT89), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n548), .A2(KEYINPUT89), .A3(KEYINPUT35), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n533), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n704), .B1(new_n713), .B2(new_n696), .ZN(new_n714));
  INV_X1    g513(.A(new_n697), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n690), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n592), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n618), .B1(new_n717), .B2(new_n713), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT44), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n720), .A2(new_n721), .A3(new_n668), .A4(new_n689), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n703), .A2(new_n722), .A3(G29gat), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n619), .A2(new_n642), .A3(new_n661), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n593), .A2(new_n724), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n725), .A2(G29gat), .A3(new_n530), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT100), .B(KEYINPUT45), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n723), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT105), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n723), .A2(new_n731), .A3(new_n728), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(G1328gat));
  NAND2_X1  g532(.A1(new_n720), .A2(new_n689), .ZN(new_n734));
  OAI21_X1  g533(.A(G36gat), .B1(new_n734), .B2(new_n472), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n471), .A2(new_n202), .ZN(new_n736));
  OAI21_X1  g535(.A(KEYINPUT46), .B1(new_n725), .B2(new_n736), .ZN(new_n737));
  OR3_X1    g536(.A1(new_n725), .A2(KEYINPUT46), .A3(new_n736), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n735), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n735), .A2(KEYINPUT106), .A3(new_n737), .A4(new_n738), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(G1329gat));
  OAI21_X1  g542(.A(G43gat), .B1(new_n734), .B2(new_n588), .ZN(new_n744));
  OR3_X1    g543(.A1(new_n725), .A2(G43gat), .A3(new_n346), .ZN(new_n745));
  XNOR2_X1  g544(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n746), .B1(new_n744), .B2(new_n745), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(G1330gat));
  OAI211_X1 g548(.A(new_n681), .B(new_n689), .C1(new_n698), .C2(new_n701), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G50gat), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n564), .A2(G50gat), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n593), .A2(new_n724), .A3(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n751), .A2(KEYINPUT48), .A3(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT108), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n753), .B(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(KEYINPUT48), .B1(new_n751), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(KEYINPUT109), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n759));
  AOI211_X1 g558(.A(new_n759), .B(KEYINPUT48), .C1(new_n751), .C2(new_n756), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n754), .B1(new_n758), .B2(new_n760), .ZN(G1331gat));
  NAND2_X1  g560(.A1(new_n551), .A2(KEYINPUT103), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n762), .A2(new_n697), .A3(new_n704), .ZN(new_n763));
  INV_X1    g562(.A(new_n688), .ZN(new_n764));
  INV_X1    g563(.A(new_n661), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n764), .A2(new_n643), .A3(new_n765), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n668), .ZN(new_n768));
  XOR2_X1   g567(.A(KEYINPUT110), .B(G57gat), .Z(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(G1332gat));
  INV_X1    g569(.A(KEYINPUT49), .ZN(new_n771));
  INV_X1    g570(.A(G64gat), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n471), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT111), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n767), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n771), .A2(new_n772), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n775), .B(new_n776), .ZN(G1333gat));
  INV_X1    g576(.A(G71gat), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n767), .A2(new_n778), .A3(new_n677), .ZN(new_n779));
  INV_X1    g578(.A(new_n588), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n767), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n781), .B2(new_n778), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n782), .B(new_n783), .ZN(G1334gat));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n681), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(G78gat), .ZN(G1335gat));
  INV_X1    g585(.A(new_n642), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n688), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT112), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n763), .A2(new_n618), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n763), .A2(KEYINPUT51), .A3(new_n618), .A4(new_n789), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n765), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n794), .A2(new_n597), .A3(new_n668), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n796));
  AOI22_X1  g595(.A1(new_n763), .A2(new_n690), .B1(new_n718), .B2(KEYINPUT44), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n789), .A2(new_n661), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n798), .ZN(new_n800));
  OAI211_X1 g599(.A(KEYINPUT113), .B(new_n800), .C1(new_n698), .C2(new_n701), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n799), .A2(new_n668), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n795), .B1(new_n802), .B2(new_n597), .ZN(G1336gat));
  NOR2_X1   g602(.A1(new_n472), .A2(G92gat), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n794), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n720), .A2(new_n800), .ZN(new_n807));
  OAI21_X1  g606(.A(G92gat), .B1(new_n807), .B2(new_n472), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n805), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n799), .A2(new_n471), .A3(new_n801), .ZN(new_n810));
  AOI22_X1  g609(.A1(new_n810), .A2(G92gat), .B1(new_n794), .B2(new_n804), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n809), .B1(new_n811), .B2(new_n806), .ZN(G1337gat));
  NAND3_X1  g611(.A1(new_n799), .A2(new_n780), .A3(new_n801), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n799), .A2(KEYINPUT114), .A3(new_n780), .A4(new_n801), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n815), .A2(G99gat), .A3(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(G99gat), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n794), .A2(new_n818), .A3(new_n677), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(G1338gat));
  NOR2_X1   g619(.A1(new_n564), .A2(G106gat), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n794), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(G106gat), .B1(new_n807), .B2(new_n564), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n799), .A2(new_n681), .A3(new_n801), .ZN(new_n826));
  AOI22_X1  g625(.A1(new_n826), .A2(G106gat), .B1(new_n794), .B2(new_n821), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n825), .B1(new_n827), .B2(new_n824), .ZN(G1339gat));
  NAND2_X1  g627(.A1(new_n662), .A2(new_n688), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n658), .B1(new_n653), .B2(KEYINPUT54), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n651), .B(new_n644), .C1(new_n647), .C2(new_n648), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n653), .A2(KEYINPUT54), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n831), .A2(KEYINPUT55), .A3(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835));
  INV_X1    g634(.A(new_n833), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n836), .B2(new_n830), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n618), .A2(new_n834), .A3(new_n659), .A4(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n226), .A2(new_n228), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n233), .A2(new_n234), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n245), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n249), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(KEYINPUT115), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n838), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n661), .A2(new_n249), .A3(new_n841), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n837), .A2(new_n834), .A3(new_n659), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n845), .B1(new_n688), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n844), .B1(new_n847), .B2(new_n619), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n829), .B1(new_n848), .B2(new_n642), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n668), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n850), .A2(new_n473), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n852), .A2(new_n303), .A3(new_n764), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n472), .A2(new_n668), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(new_n346), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n849), .A2(new_n856), .A3(new_n564), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n856), .B1(new_n849), .B2(new_n564), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n855), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT117), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n861), .B(new_n855), .C1(new_n857), .C2(new_n858), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n860), .A2(new_n250), .A3(new_n862), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n863), .A2(KEYINPUT118), .A3(G113gat), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT118), .B1(new_n863), .B2(G113gat), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n853), .B1(new_n864), .B2(new_n865), .ZN(G1340gat));
  AOI21_X1  g665(.A(G120gat), .B1(new_n852), .B2(new_n661), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n860), .A2(new_n862), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n765), .A2(new_n300), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(G1341gat));
  NAND3_X1  g669(.A1(new_n852), .A2(new_n309), .A3(new_n642), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n868), .A2(new_n642), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n871), .B1(new_n872), .B2(new_n309), .ZN(G1342gat));
  NOR3_X1   g672(.A1(new_n851), .A2(G134gat), .A3(new_n619), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT56), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n868), .A2(new_n618), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n876), .B2(new_n307), .ZN(G1343gat));
  NOR2_X1   g676(.A1(new_n780), .A2(new_n854), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n837), .A2(new_n834), .A3(new_n250), .A4(new_n659), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n618), .B1(new_n845), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n787), .B1(new_n880), .B2(new_n844), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n829), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n564), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT57), .B1(new_n849), .B2(new_n681), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n885), .B1(new_n886), .B2(KEYINPUT119), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n834), .A2(new_n659), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n888), .A2(new_n686), .A3(new_n687), .A4(new_n837), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n618), .B1(new_n889), .B2(new_n845), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n787), .B1(new_n890), .B2(new_n844), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n564), .B1(new_n891), .B2(new_n829), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n892), .A2(new_n893), .A3(KEYINPUT57), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n764), .B(new_n878), .C1(new_n887), .C2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(G141gat), .ZN(new_n896));
  INV_X1    g695(.A(new_n850), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n780), .A2(new_n564), .A3(new_n471), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n360), .A3(new_n250), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(KEYINPUT58), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n250), .B(new_n878), .C1(new_n887), .C2(new_n894), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT120), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n893), .B1(new_n892), .B2(KEYINPUT57), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n886), .A2(KEYINPUT119), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n907), .A2(new_n908), .A3(new_n885), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n909), .A2(KEYINPUT120), .A3(new_n250), .A4(new_n878), .ZN(new_n910));
  AND3_X1   g709(.A1(new_n906), .A2(G141gat), .A3(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT58), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n901), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n903), .B1(new_n911), .B2(new_n913), .ZN(G1344gat));
  NAND3_X1  g713(.A1(new_n900), .A2(new_n362), .A3(new_n661), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT59), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n878), .A2(new_n661), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n662), .A2(new_n251), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n881), .A2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n564), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n881), .A2(KEYINPUT121), .A3(new_n918), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(new_n883), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n849), .A2(new_n884), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n917), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n362), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT57), .B1(new_n921), .B2(new_n922), .ZN(new_n929));
  INV_X1    g728(.A(new_n925), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(KEYINPUT122), .B1(new_n931), .B2(new_n917), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n916), .B1(new_n928), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n916), .A2(G148gat), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n909), .A2(new_n878), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n935), .B2(new_n661), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n915), .B1(new_n933), .B2(new_n936), .ZN(G1345gat));
  AOI21_X1  g736(.A(new_n351), .B1(new_n935), .B2(new_n642), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n899), .A2(G155gat), .A3(new_n787), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n938), .A2(new_n939), .ZN(G1346gat));
  AOI21_X1  g739(.A(G162gat), .B1(new_n900), .B2(new_n618), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n619), .A2(new_n352), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n941), .B1(new_n935), .B2(new_n942), .ZN(G1347gat));
  NOR2_X1   g742(.A1(new_n472), .A2(new_n668), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n945), .A2(new_n708), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n849), .A2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(G169gat), .B1(new_n948), .B2(new_n764), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n677), .B(new_n944), .C1(new_n857), .C2(new_n858), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n251), .A2(new_n255), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(G1348gat));
  OAI21_X1  g752(.A(G176gat), .B1(new_n950), .B2(new_n765), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n948), .A2(new_n256), .A3(new_n661), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1349gat));
  OAI21_X1  g755(.A(G183gat), .B1(new_n950), .B2(new_n787), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n948), .A2(new_n275), .A3(new_n642), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g759(.A1(new_n948), .A2(new_n269), .A3(new_n618), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n951), .A2(new_n618), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n963));
  AND4_X1   g762(.A1(KEYINPUT123), .A2(new_n962), .A3(new_n963), .A4(G190gat), .ZN(new_n964));
  OAI21_X1  g763(.A(G190gat), .B1(new_n963), .B2(KEYINPUT123), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  AOI22_X1  g765(.A1(new_n962), .A2(new_n966), .B1(KEYINPUT123), .B2(new_n963), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n961), .B1(new_n964), .B2(new_n967), .ZN(G1351gat));
  NOR2_X1   g767(.A1(new_n780), .A2(new_n945), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n849), .A2(new_n681), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g769(.A(G197gat), .B1(new_n970), .B2(new_n764), .ZN(new_n971));
  NOR3_X1   g770(.A1(new_n931), .A2(new_n780), .A3(new_n945), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n250), .A2(G197gat), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(G1352gat));
  INV_X1    g773(.A(KEYINPUT62), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n975), .A2(KEYINPUT125), .ZN(new_n976));
  XNOR2_X1  g775(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n977));
  XNOR2_X1  g776(.A(KEYINPUT124), .B(G204gat), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n765), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n970), .A2(new_n979), .ZN(new_n980));
  MUX2_X1   g779(.A(new_n976), .B(new_n977), .S(new_n980), .Z(new_n981));
  OAI21_X1  g780(.A(new_n969), .B1(new_n929), .B2(new_n930), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n978), .B1(new_n982), .B2(new_n765), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT126), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n981), .A2(KEYINPUT126), .A3(new_n983), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n986), .A2(new_n987), .ZN(G1353gat));
  INV_X1    g787(.A(new_n970), .ZN(new_n989));
  OR3_X1    g788(.A1(new_n989), .A2(G211gat), .A3(new_n787), .ZN(new_n990));
  OAI211_X1 g789(.A(new_n642), .B(new_n969), .C1(new_n929), .C2(new_n930), .ZN(new_n991));
  AND3_X1   g790(.A1(new_n991), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n992));
  AOI21_X1  g791(.A(KEYINPUT63), .B1(new_n991), .B2(G211gat), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n990), .B1(new_n992), .B2(new_n993), .ZN(G1354gat));
  OAI21_X1  g793(.A(G218gat), .B1(new_n982), .B2(new_n619), .ZN(new_n995));
  OR3_X1    g794(.A1(new_n989), .A2(G218gat), .A3(new_n619), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n997), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


