//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1207,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  INV_X1    g0011(.A(G107), .ZN(new_n212));
  INV_X1    g0012(.A(G264), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G97), .A2(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI211_X1 g0020(.A(new_n214), .B(new_n220), .C1(G116), .C2(G270), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G77), .A2(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G226), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n221), .B(new_n222), .C1(new_n202), .C2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G58), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n208), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  INV_X1    g0031(.A(G20), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(G50), .B1(G58), .B2(G68), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n211), .B(new_n230), .C1(new_n233), .C2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT66), .B(G264), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n240), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n202), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G58), .ZN(new_n248));
  XOR2_X1   g0048(.A(G107), .B(G116), .Z(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(KEYINPUT76), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT14), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n256), .B(G274), .C1(G41), .C2(G45), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n257), .B(KEYINPUT67), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT3), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(G232), .A3(G1698), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G97), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n264), .B(new_n265), .C1(new_n267), .C2(new_n223), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G1), .A3(G13), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n258), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT13), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G238), .ZN(new_n277));
  AND3_X1   g0077(.A1(new_n272), .A2(new_n273), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n273), .B1(new_n272), .B2(new_n277), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G169), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n255), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(G179), .ZN(new_n283));
  OAI221_X1 g0083(.A(G169), .B1(new_n253), .B2(new_n254), .C1(new_n278), .C2(new_n279), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT71), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT70), .ZN(new_n288));
  AND3_X1   g0088(.A1(new_n287), .A2(new_n288), .A3(new_n231), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n288), .B1(new_n287), .B2(new_n231), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n286), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n287), .A2(new_n231), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT70), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n287), .A2(new_n288), .A3(new_n231), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(KEYINPUT71), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n216), .A2(G20), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n232), .A2(G33), .ZN(new_n299));
  NOR2_X1   g0099(.A1(G20), .A2(G33), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  OAI221_X1 g0101(.A(new_n298), .B1(new_n299), .B2(new_n205), .C1(new_n301), .C2(new_n202), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT73), .ZN(new_n304));
  INV_X1    g0104(.A(G13), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(G1), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G20), .ZN(new_n307));
  AND4_X1   g0107(.A1(new_n304), .A2(new_n293), .A3(new_n294), .A4(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n293), .A2(new_n294), .ZN(new_n310));
  INV_X1    g0110(.A(new_n307), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT73), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n309), .A2(new_n312), .B1(new_n256), .B2(G20), .ZN(new_n313));
  AOI22_X1  g0113(.A1(KEYINPUT11), .A2(new_n303), .B1(new_n313), .B2(G68), .ZN(new_n314));
  OR2_X1    g0114(.A1(new_n303), .A2(KEYINPUT11), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n306), .A2(G20), .A3(new_n216), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT75), .B(KEYINPUT12), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(KEYINPUT75), .A2(KEYINPUT12), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n314), .A2(new_n315), .A3(new_n319), .A4(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n285), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G200), .ZN(new_n324));
  INV_X1    g0124(.A(new_n279), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n272), .A2(new_n273), .A3(new_n277), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G190), .ZN(new_n328));
  NOR3_X1   g0128(.A1(new_n278), .A2(new_n279), .A3(new_n328), .ZN(new_n329));
  OR3_X1    g0129(.A1(new_n322), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n323), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n296), .A2(new_n307), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT72), .ZN(new_n333));
  XOR2_X1   g0133(.A(KEYINPUT8), .B(G58), .Z(new_n334));
  NAND2_X1  g0134(.A1(new_n256), .A2(G20), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n311), .B1(new_n291), .B2(new_n295), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT72), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n333), .A2(new_n334), .A3(new_n335), .A4(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n261), .A2(new_n232), .A3(new_n262), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT7), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT77), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n261), .A2(KEYINPUT7), .A3(new_n232), .A4(new_n262), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n340), .A2(KEYINPUT77), .A3(new_n341), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(G68), .A3(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n225), .A2(new_n216), .ZN(new_n348));
  OAI21_X1  g0148(.A(G20), .B1(new_n348), .B2(new_n201), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n300), .A2(G159), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n347), .A2(KEYINPUT16), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT16), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n216), .B1(new_n342), .B2(new_n344), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n354), .B1(new_n355), .B2(new_n351), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n353), .A2(new_n310), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n334), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n311), .ZN(new_n359));
  AND3_X1   g0159(.A1(new_n339), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n263), .B1(G226), .B2(new_n266), .ZN(new_n361));
  NOR2_X1   g0161(.A1(G223), .A2(G1698), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n361), .A2(new_n362), .B1(new_n260), .B2(new_n218), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n271), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT67), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n257), .B(new_n365), .ZN(new_n366));
  OR3_X1    g0166(.A1(new_n275), .A2(KEYINPUT78), .A3(new_n226), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT78), .B1(new_n275), .B2(new_n226), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n364), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(G200), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n364), .A2(new_n369), .A3(G190), .A4(new_n366), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n360), .A2(KEYINPUT17), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT17), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n339), .A2(new_n357), .A3(new_n372), .A4(new_n359), .ZN(new_n375));
  INV_X1    g0175(.A(new_n371), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n339), .A2(new_n357), .A3(new_n359), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n370), .A2(G169), .ZN(new_n379));
  INV_X1    g0179(.A(G179), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n379), .B1(new_n380), .B2(new_n370), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n378), .A2(new_n381), .A3(KEYINPUT18), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT18), .B1(new_n378), .B2(new_n381), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n373), .B(new_n377), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  AND2_X1   g0184(.A1(KEYINPUT3), .A2(G33), .ZN(new_n385));
  NOR2_X1   g0185(.A1(KEYINPUT3), .A2(G33), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n387), .A2(G1698), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n388), .A2(G232), .B1(G107), .B2(new_n387), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n263), .A2(G1698), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n389), .B1(new_n217), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n271), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n276), .A2(G244), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(new_n366), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n395), .A2(new_n324), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n289), .A2(new_n290), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n334), .A2(new_n300), .B1(G20), .B2(G77), .ZN(new_n398));
  XOR2_X1   g0198(.A(KEYINPUT15), .B(G87), .Z(new_n399));
  NAND3_X1  g0199(.A1(new_n399), .A2(new_n232), .A3(G33), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n397), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n401), .B1(new_n313), .B2(G77), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n311), .A2(new_n205), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n402), .B(new_n403), .C1(new_n394), .C2(new_n328), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n396), .A2(new_n404), .ZN(new_n405));
  OR3_X1    g0205(.A1(new_n331), .A2(new_n384), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n388), .A2(G222), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT69), .ZN(new_n408));
  XNOR2_X1  g0208(.A(new_n407), .B(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(G223), .ZN(new_n410));
  OAI22_X1  g0210(.A1(new_n390), .A2(new_n410), .B1(new_n205), .B2(new_n263), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n271), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n366), .B1(new_n223), .B2(new_n275), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n413), .B(KEYINPUT68), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n415), .A2(new_n328), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(G200), .B2(new_n415), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT74), .ZN(new_n418));
  AOI21_X1  g0218(.A(KEYINPUT10), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n311), .A2(new_n202), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n204), .A2(new_n232), .ZN(new_n421));
  INV_X1    g0221(.A(G150), .ZN(new_n422));
  OAI22_X1  g0222(.A1(new_n358), .A2(new_n299), .B1(new_n422), .B2(new_n301), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n297), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n333), .A2(new_n335), .A3(new_n338), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n420), .B(new_n424), .C1(new_n425), .C2(new_n202), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n426), .B(KEYINPUT9), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n417), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n419), .A2(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n427), .B(new_n417), .C1(new_n418), .C2(KEYINPUT10), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n415), .A2(G179), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(new_n281), .B2(new_n415), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n426), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n429), .A2(new_n430), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n395), .A2(new_n380), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n402), .A2(new_n403), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n394), .A2(new_n281), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NOR3_X1   g0239(.A1(new_n406), .A2(new_n434), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(G33), .A2(G116), .ZN(new_n442));
  OAI22_X1  g0242(.A1(new_n385), .A2(new_n386), .B1(G244), .B2(new_n266), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n217), .A2(new_n266), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n442), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT80), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT80), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n448), .B(new_n442), .C1(new_n443), .C2(new_n445), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n447), .A2(new_n271), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G45), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n219), .B1(new_n451), .B2(G1), .ZN(new_n452));
  INV_X1    g0252(.A(G274), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n256), .A2(new_n453), .A3(G45), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n270), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  XOR2_X1   g0255(.A(new_n455), .B(KEYINPUT79), .Z(new_n456));
  AND3_X1   g0256(.A1(new_n450), .A2(G179), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n281), .B1(new_n450), .B2(new_n456), .ZN(new_n458));
  OAI21_X1  g0258(.A(KEYINPUT81), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT81), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n450), .A2(new_n456), .A3(G179), .ZN(new_n461));
  XNOR2_X1  g0261(.A(new_n455), .B(KEYINPUT79), .ZN(new_n462));
  INV_X1    g0262(.A(new_n449), .ZN(new_n463));
  OAI221_X1 g0263(.A(new_n444), .B1(G244), .B2(new_n266), .C1(new_n385), .C2(new_n386), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n448), .B1(new_n464), .B2(new_n442), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n462), .B1(new_n466), .B2(new_n271), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n460), .B(new_n461), .C1(new_n467), .C2(new_n281), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT19), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n232), .B1(new_n265), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(G97), .A2(G107), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n218), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  OR2_X1    g0273(.A1(new_n473), .A2(KEYINPUT82), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n263), .A2(new_n232), .A3(G68), .ZN(new_n475));
  INV_X1    g0275(.A(G97), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n469), .B1(new_n299), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n473), .A2(KEYINPUT82), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n474), .A2(new_n475), .A3(new_n477), .A4(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n399), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n479), .A2(new_n310), .B1(new_n311), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n260), .A2(G1), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n336), .A2(new_n483), .A3(new_n399), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n459), .A2(new_n468), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(G244), .B1(new_n385), .B2(new_n386), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT4), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n487), .A2(new_n488), .B1(G33), .B2(G283), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n263), .A2(KEYINPUT4), .A3(G244), .A4(new_n266), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n263), .A2(G250), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n266), .B1(new_n492), .B2(KEYINPUT4), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n271), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  AND2_X1   g0294(.A1(KEYINPUT5), .A2(G41), .ZN(new_n495));
  NOR2_X1   g0295(.A1(KEYINPUT5), .A2(G41), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n256), .B(G45), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  OR2_X1    g0297(.A1(new_n497), .A2(new_n453), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n497), .A2(G257), .A3(new_n270), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n494), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G200), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n300), .A2(G77), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT6), .ZN(new_n504));
  NOR3_X1   g0304(.A1(new_n504), .A2(new_n476), .A3(G107), .ZN(new_n505));
  XNOR2_X1  g0305(.A(G97), .B(G107), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n505), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n503), .B1(new_n507), .B2(new_n232), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n212), .B1(new_n342), .B2(new_n344), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n310), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n311), .A2(new_n476), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n296), .A2(G97), .A3(new_n307), .A4(new_n483), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n494), .A2(G190), .A3(new_n498), .A4(new_n500), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n502), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n510), .A2(new_n512), .A3(new_n511), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n494), .A2(new_n380), .A3(new_n498), .A4(new_n500), .ZN(new_n517));
  INV_X1    g0317(.A(new_n498), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n488), .B1(new_n263), .B2(G250), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n489), .B(new_n490), .C1(new_n266), .C2(new_n519), .ZN(new_n520));
  AOI211_X1 g0320(.A(new_n499), .B(new_n518), .C1(new_n520), .C2(new_n271), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n516), .B(new_n517), .C1(new_n521), .C2(G169), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n515), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n296), .A2(G87), .A3(new_n307), .A4(new_n483), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT83), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT83), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n336), .A2(new_n526), .A3(G87), .A4(new_n483), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n450), .A2(new_n456), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G200), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n450), .A2(new_n456), .A3(G190), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n528), .A2(new_n481), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n486), .A2(new_n523), .A3(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n263), .B1(G250), .B2(G1698), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n266), .A2(G257), .ZN(new_n536));
  INV_X1    g0336(.A(G294), .ZN(new_n537));
  OAI22_X1  g0337(.A1(new_n535), .A2(new_n536), .B1(new_n260), .B2(new_n537), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n497), .A2(new_n270), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n538), .A2(new_n271), .B1(G264), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n498), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n281), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(G179), .B2(new_n541), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n232), .B(G87), .C1(new_n385), .C2(new_n386), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT84), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n263), .A2(KEYINPUT84), .A3(new_n232), .A4(G87), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT22), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT85), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT85), .A4(KEYINPUT22), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g0353(.A(KEYINPUT86), .B(KEYINPUT22), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n545), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT24), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n212), .A2(KEYINPUT23), .A3(G20), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT23), .B1(new_n212), .B2(G20), .ZN(new_n561));
  OAI22_X1  g0361(.A1(new_n560), .A2(new_n561), .B1(G20), .B2(new_n442), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n557), .A2(new_n558), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n555), .B1(new_n551), .B2(new_n552), .ZN(new_n565));
  OAI21_X1  g0365(.A(KEYINPUT24), .B1(new_n565), .B2(new_n562), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n397), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n332), .A2(new_n212), .A3(new_n482), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n306), .A2(G20), .A3(new_n212), .ZN(new_n569));
  XNOR2_X1  g0369(.A(new_n569), .B(KEYINPUT25), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n544), .B1(new_n567), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n558), .B1(new_n557), .B2(new_n563), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n565), .A2(KEYINPUT24), .A3(new_n562), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n310), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n541), .A2(G200), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n541), .A2(new_n328), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n576), .A2(new_n571), .A3(new_n577), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n266), .A2(G257), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n263), .B(new_n581), .C1(new_n213), .C2(new_n266), .ZN(new_n582));
  INV_X1    g0382(.A(G303), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n387), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n582), .A2(new_n271), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n497), .A2(G270), .A3(new_n270), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n585), .A2(G190), .A3(new_n498), .A4(new_n586), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n585), .A2(new_n498), .A3(new_n586), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n587), .B1(new_n588), .B2(new_n324), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n304), .B1(new_n397), .B2(new_n307), .ZN(new_n590));
  OAI211_X1 g0390(.A(G116), .B(new_n483), .C1(new_n590), .C2(new_n308), .ZN(new_n591));
  NAND2_X1  g0391(.A1(G33), .A2(G283), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n592), .B(new_n232), .C1(G33), .C2(new_n476), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n593), .B(new_n292), .C1(new_n232), .C2(G116), .ZN(new_n594));
  XOR2_X1   g0394(.A(new_n594), .B(KEYINPUT20), .Z(new_n595));
  INV_X1    g0395(.A(G116), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n306), .A2(G20), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n591), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  OR2_X1    g0398(.A1(new_n589), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(G179), .A3(new_n588), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT21), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n588), .A2(new_n281), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n598), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n601), .B1(new_n598), .B2(new_n602), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n599), .B(new_n600), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n534), .A2(new_n573), .A3(new_n580), .A4(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n441), .A2(new_n607), .ZN(G372));
  OR2_X1    g0408(.A1(new_n382), .A2(new_n383), .ZN(new_n609));
  INV_X1    g0409(.A(new_n323), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n330), .B1(new_n610), .B2(new_n439), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n373), .A2(new_n377), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n609), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n429), .A2(new_n430), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n613), .A2(new_n614), .B1(new_n426), .B2(new_n432), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n461), .B1(new_n467), .B2(new_n281), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n485), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n617), .A2(new_n532), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT26), .ZN(new_n619));
  INV_X1    g0419(.A(new_n522), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n459), .A2(new_n468), .A3(new_n485), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n622), .A2(new_n620), .A3(new_n532), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(KEYINPUT26), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n621), .A2(new_n624), .A3(new_n617), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n543), .B1(new_n576), .B2(new_n571), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n600), .B1(new_n603), .B2(new_n604), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n618), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n523), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n580), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(KEYINPUT87), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  NOR3_X1   g0431(.A1(new_n567), .A2(new_n572), .A3(new_n578), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n523), .B1(new_n632), .B2(new_n577), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n617), .A2(new_n532), .ZN(new_n634));
  INV_X1    g0434(.A(new_n600), .ZN(new_n635));
  INV_X1    g0435(.A(new_n604), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n598), .A2(new_n602), .A3(new_n601), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n634), .B1(new_n573), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT87), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n633), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n625), .B1(new_n631), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n615), .B1(new_n441), .B2(new_n642), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n643), .B(KEYINPUT88), .ZN(G369));
  INV_X1    g0444(.A(G330), .ZN(new_n645));
  INV_X1    g0445(.A(new_n306), .ZN(new_n646));
  OR3_X1    g0446(.A1(new_n646), .A2(KEYINPUT27), .A3(G20), .ZN(new_n647));
  OAI21_X1  g0447(.A(KEYINPUT27), .B1(new_n646), .B2(G20), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(G213), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(G343), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n598), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT89), .B1(new_n605), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n627), .A2(new_n652), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n627), .A2(KEYINPUT89), .A3(new_n652), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n645), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n657), .A2(KEYINPUT90), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(KEYINPUT90), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n580), .A2(new_n573), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n651), .B1(new_n567), .B2(new_n572), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n626), .A2(new_n651), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n651), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n626), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n638), .A2(new_n651), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n661), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n666), .A2(new_n668), .A3(new_n670), .ZN(G399));
  NOR2_X1   g0471(.A1(new_n472), .A2(G116), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT91), .ZN(new_n673));
  INV_X1    g0473(.A(new_n209), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(G41), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n673), .A2(new_n256), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n676), .B1(new_n235), .B2(new_n675), .ZN(new_n677));
  XOR2_X1   g0477(.A(new_n677), .B(KEYINPUT28), .Z(new_n678));
  NOR3_X1   g0478(.A1(new_n642), .A2(KEYINPUT29), .A3(new_n651), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT29), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT93), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n618), .A2(new_n681), .A3(KEYINPUT26), .A4(new_n620), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n620), .A2(new_n617), .A3(KEYINPUT26), .A4(new_n532), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(KEYINPUT93), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n623), .A2(new_n619), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT94), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n623), .A2(KEYINPUT94), .A3(new_n619), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n685), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n633), .A2(new_n639), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(new_n617), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n680), .B1(new_n692), .B2(new_n667), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n679), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n585), .A2(new_n498), .A3(new_n586), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n541), .A2(new_n529), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n521), .A2(G179), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(KEYINPUT92), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT30), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n521), .A2(new_n588), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n457), .A2(new_n540), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n501), .A2(new_n695), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n704), .A2(KEYINPUT30), .A3(new_n540), .A4(new_n457), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT92), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n501), .A2(new_n380), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n706), .B1(new_n696), .B2(new_n707), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n699), .A2(new_n703), .A3(new_n705), .A4(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n651), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT31), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n703), .A2(new_n705), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n696), .A2(new_n707), .ZN(new_n714));
  OAI211_X1 g0514(.A(KEYINPUT31), .B(new_n651), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n712), .B(new_n715), .C1(new_n607), .C2(new_n651), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G330), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n694), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n678), .B1(new_n719), .B2(G1), .ZN(G364));
  AOI21_X1  g0520(.A(new_n231), .B1(G20), .B2(new_n281), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n232), .A2(G179), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(new_n328), .A3(new_n324), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT97), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n724), .A2(KEYINPUT97), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n722), .A2(new_n328), .A3(G200), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n729), .A2(G329), .B1(G283), .B2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT98), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n328), .A2(G200), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n380), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G20), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n732), .A2(new_n733), .B1(G294), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(G322), .ZN(new_n738));
  NAND2_X1  g0538(.A1(G20), .A2(G179), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT95), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n734), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n737), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n740), .A2(new_n328), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n324), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G317), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n745), .B1(KEYINPUT33), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(KEYINPUT33), .B2(new_n746), .ZN(new_n748));
  INV_X1    g0548(.A(G311), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n743), .A2(G200), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI221_X1 g0551(.A(new_n748), .B1(new_n749), .B2(new_n751), .C1(new_n733), .C2(new_n732), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n328), .A2(new_n324), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n740), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n755), .A2(G326), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n753), .A2(new_n722), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n387), .B1(new_n757), .B2(new_n583), .ZN(new_n758));
  XOR2_X1   g0558(.A(new_n758), .B(KEYINPUT96), .Z(new_n759));
  NOR4_X1   g0559(.A1(new_n742), .A2(new_n752), .A3(new_n756), .A4(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n741), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n387), .B1(new_n761), .B2(G58), .ZN(new_n762));
  INV_X1    g0562(.A(new_n757), .ZN(new_n763));
  AOI22_X1  g0563(.A1(G97), .A2(new_n736), .B1(new_n763), .B2(G87), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n762), .B(new_n764), .C1(new_n745), .C2(new_n216), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n751), .A2(new_n205), .B1(new_n212), .B2(new_n730), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n754), .A2(new_n202), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n724), .A2(G159), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT32), .ZN(new_n769));
  NOR4_X1   g0569(.A1(new_n765), .A2(new_n766), .A3(new_n767), .A4(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n721), .B1(new_n760), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n263), .A2(G355), .A3(new_n209), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n248), .A2(new_n451), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n674), .A2(new_n263), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(G45), .B2(new_n234), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n772), .B1(G116), .B2(new_n209), .C1(new_n773), .C2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G13), .A2(G33), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n721), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n655), .A2(new_n656), .ZN(new_n782));
  INV_X1    g0582(.A(new_n779), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n771), .B(new_n781), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n658), .B(new_n659), .C1(G330), .C2(new_n782), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n305), .A2(G20), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n256), .B1(new_n786), .B2(G45), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n675), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  MUX2_X1   g0590(.A(new_n784), .B(new_n785), .S(new_n790), .Z(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT99), .ZN(G396));
  NAND2_X1  g0592(.A1(new_n631), .A2(new_n641), .ZN(new_n793));
  INV_X1    g0593(.A(new_n625), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n651), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n667), .B1(new_n402), .B2(new_n403), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n438), .B1(new_n405), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n439), .A2(new_n667), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n795), .B(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n717), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT100), .Z(new_n803));
  AOI21_X1  g0603(.A(new_n789), .B1(new_n801), .B2(new_n717), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n721), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n728), .A2(new_n749), .ZN(new_n807));
  INV_X1    g0607(.A(new_n736), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n476), .A2(new_n808), .B1(new_n754), .B2(new_n583), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n730), .A2(new_n218), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n807), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n744), .A2(G283), .B1(new_n761), .B2(G294), .ZN(new_n812));
  AND3_X1   g0612(.A1(new_n811), .A2(new_n387), .A3(new_n812), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n813), .B1(new_n212), .B2(new_n757), .C1(new_n596), .C2(new_n751), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n744), .A2(G150), .B1(new_n761), .B2(G143), .ZN(new_n815));
  INV_X1    g0615(.A(G137), .ZN(new_n816));
  INV_X1    g0616(.A(G159), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n815), .B1(new_n816), .B2(new_n754), .C1(new_n817), .C2(new_n751), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT34), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n808), .A2(new_n225), .B1(new_n757), .B2(new_n202), .ZN(new_n820));
  INV_X1    g0620(.A(G132), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n263), .B1(new_n728), .B2(new_n821), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n820), .B(new_n822), .C1(G68), .C2(new_n731), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n806), .B1(new_n814), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n721), .A2(new_n777), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n790), .B(new_n825), .C1(new_n205), .C2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n778), .B2(new_n800), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n805), .A2(new_n828), .ZN(G384));
  NAND3_X1  g0629(.A1(new_n709), .A2(KEYINPUT31), .A3(new_n651), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n712), .B(new_n830), .C1(new_n607), .C2(new_n651), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n322), .A2(new_n651), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n323), .A2(new_n330), .A3(new_n832), .ZN(new_n833));
  NOR3_X1   g0633(.A1(new_n322), .A2(new_n329), .A3(new_n327), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n322), .B(new_n651), .C1(new_n834), .C2(new_n285), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n799), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT103), .ZN(new_n838));
  INV_X1    g0638(.A(new_n649), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n347), .A2(new_n352), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n354), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n841), .A2(new_n297), .A3(new_n353), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n842), .A2(new_n359), .A3(new_n339), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n384), .A2(new_n839), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n360), .A2(new_n371), .A3(new_n372), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT37), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n379), .B(new_n649), .C1(new_n380), .C2(new_n370), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n378), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n375), .A2(new_n376), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(new_n847), .B2(new_n843), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n849), .B1(new_n851), .B2(new_n846), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT38), .B1(new_n844), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n844), .A2(new_n852), .A3(KEYINPUT38), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n837), .A2(new_n838), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n831), .B(new_n836), .C1(KEYINPUT103), .C2(KEYINPUT40), .ZN(new_n857));
  AND3_X1   g0657(.A1(new_n844), .A2(new_n852), .A3(KEYINPUT38), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n384), .A2(new_n378), .A3(new_n839), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n845), .A2(new_n848), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT37), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n849), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT38), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n831), .B(new_n836), .C1(new_n858), .C2(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n856), .A2(new_n857), .B1(KEYINPUT40), .B2(new_n864), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT104), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n440), .A2(new_n831), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n866), .B(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(G330), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n440), .B1(new_n679), .B2(new_n693), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n615), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n869), .B(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT102), .ZN(new_n873));
  INV_X1    g0673(.A(new_n798), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(new_n795), .B2(new_n800), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n833), .A2(new_n835), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n873), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n854), .A2(new_n855), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n628), .A2(KEYINPUT87), .A3(new_n630), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n640), .B1(new_n633), .B2(new_n639), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n794), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n882), .A2(new_n667), .A3(new_n800), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n798), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n884), .A2(KEYINPUT102), .A3(new_n876), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n878), .A2(new_n879), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n609), .A2(new_n839), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n854), .A2(KEYINPUT39), .A3(new_n855), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT39), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n858), .B2(new_n863), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n323), .A2(new_n651), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n887), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n886), .A2(new_n894), .ZN(new_n895));
  XOR2_X1   g0695(.A(new_n872), .B(new_n895), .Z(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n256), .B2(new_n786), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n507), .B(KEYINPUT101), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n596), .B1(new_n898), .B2(KEYINPUT35), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n899), .B(new_n233), .C1(KEYINPUT35), .C2(new_n898), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT36), .ZN(new_n901));
  OAI21_X1  g0701(.A(G77), .B1(new_n225), .B2(new_n216), .ZN(new_n902));
  OAI22_X1  g0702(.A1(new_n902), .A2(new_n234), .B1(G50), .B2(new_n216), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(G1), .A3(new_n305), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n897), .A2(new_n901), .A3(new_n904), .ZN(G367));
  OAI21_X1  g0705(.A(new_n629), .B1(new_n513), .B2(new_n667), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n670), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n907), .B(KEYINPUT42), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n522), .B1(new_n906), .B2(new_n573), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n667), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n667), .B1(new_n528), .B2(new_n481), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n912), .A2(new_n485), .A3(new_n616), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n634), .B2(new_n912), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n620), .A2(new_n651), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n906), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n660), .A2(new_n665), .A3(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n911), .A2(new_n919), .A3(new_n915), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n923), .B(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n675), .B(KEYINPUT41), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n666), .A2(KEYINPUT108), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT108), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n660), .A2(new_n929), .A3(new_n665), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n918), .B1(new_n670), .B2(new_n668), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT44), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n670), .A2(new_n668), .A3(new_n918), .ZN(new_n933));
  XNOR2_X1  g0733(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT106), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n933), .B(new_n935), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n928), .A2(new_n930), .A3(new_n932), .A4(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n932), .A2(new_n936), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n938), .A2(KEYINPUT108), .A3(new_n666), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n665), .A2(new_n669), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT107), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n670), .B(new_n941), .C1(new_n660), .C2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n670), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n944), .A2(KEYINPUT107), .A3(new_n658), .A4(new_n659), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n946), .A2(new_n718), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n940), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n927), .B1(new_n948), .B2(new_n719), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n925), .B1(new_n949), .B2(new_n788), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n750), .A2(G50), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n763), .A2(G58), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n755), .A2(G143), .ZN(new_n953));
  AOI22_X1  g0753(.A1(G77), .A2(new_n731), .B1(new_n736), .B2(G68), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n951), .A2(new_n952), .A3(new_n953), .A4(new_n954), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n745), .A2(new_n817), .B1(new_n816), .B2(new_n723), .ZN(new_n956));
  NOR3_X1   g0756(.A1(new_n955), .A2(new_n956), .A3(new_n387), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n422), .B2(new_n741), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT111), .Z(new_n959));
  XNOR2_X1  g0759(.A(KEYINPUT110), .B(G317), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n724), .A2(new_n960), .B1(new_n731), .B2(G97), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n961), .B1(new_n212), .B2(new_n808), .C1(new_n745), .C2(new_n537), .ZN(new_n962));
  AOI21_X1  g0762(.A(KEYINPUT46), .B1(new_n763), .B2(G116), .ZN(new_n963));
  INV_X1    g0763(.A(G283), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n751), .A2(new_n964), .ZN(new_n965));
  NOR4_X1   g0765(.A1(new_n962), .A2(new_n263), .A3(new_n963), .A4(new_n965), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n966), .B1(new_n583), .B2(new_n741), .C1(new_n749), .C2(new_n754), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n763), .A2(KEYINPUT46), .A3(G116), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(KEYINPUT109), .Z(new_n969));
  OAI21_X1  g0769(.A(new_n959), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT47), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n721), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n914), .A2(new_n783), .ZN(new_n973));
  INV_X1    g0773(.A(new_n774), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n780), .B1(new_n209), .B2(new_n480), .C1(new_n244), .C2(new_n974), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n972), .A2(new_n789), .A3(new_n973), .A4(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n950), .A2(new_n976), .ZN(G387));
  INV_X1    g0777(.A(new_n946), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n663), .A2(new_n664), .A3(new_n779), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n774), .B1(new_n240), .B2(new_n451), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n673), .A2(new_n209), .A3(new_n263), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n673), .A2(G45), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n334), .A2(new_n202), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT50), .Z(new_n985));
  OAI211_X1 g0785(.A(new_n983), .B(new_n985), .C1(new_n216), .C2(new_n205), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n982), .A2(new_n986), .B1(new_n212), .B2(new_n674), .ZN(new_n987));
  INV_X1    g0787(.A(new_n780), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n789), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n263), .B1(new_n422), .B2(new_n723), .C1(new_n751), .C2(new_n216), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n808), .A2(new_n480), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n992), .B1(new_n205), .B2(new_n757), .C1(new_n754), .C2(new_n817), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n745), .A2(new_n358), .B1(new_n476), .B2(new_n730), .ZN(new_n994));
  NOR3_X1   g0794(.A1(new_n990), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n202), .B2(new_n741), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n750), .A2(G303), .B1(new_n755), .B2(G322), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n761), .A2(new_n960), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n997), .B(new_n998), .C1(new_n749), .C2(new_n745), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT48), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n964), .B2(new_n808), .C1(new_n537), .C2(new_n757), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT49), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n731), .A2(G116), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n724), .A2(G326), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1003), .A2(new_n387), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  AND2_X1   g0806(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n996), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n989), .B1(new_n1008), .B2(new_n721), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n978), .A2(new_n788), .B1(new_n979), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n675), .B1(new_n978), .B2(new_n719), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1010), .B1(new_n1011), .B2(new_n947), .ZN(G393));
  NAND2_X1  g0812(.A1(new_n940), .A2(new_n788), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n749), .A2(new_n741), .B1(new_n754), .B2(new_n746), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT52), .Z(new_n1015));
  OAI22_X1  g0815(.A1(new_n745), .A2(new_n583), .B1(new_n212), .B2(new_n730), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n387), .B1(new_n757), .B2(new_n964), .C1(new_n808), .C2(new_n596), .ZN(new_n1017));
  NOR3_X1   g0817(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n537), .B2(new_n751), .C1(new_n738), .C2(new_n723), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n422), .A2(new_n754), .B1(new_n741), .B2(new_n817), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT51), .Z(new_n1021));
  OAI21_X1  g0821(.A(new_n263), .B1(new_n751), .B2(new_n358), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G143), .A2(new_n724), .B1(new_n736), .B2(G77), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n218), .B2(new_n730), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1025), .B1(new_n202), .B2(new_n745), .C1(new_n216), .C2(new_n757), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n806), .B1(new_n1019), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n780), .B1(new_n251), .B2(new_n974), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G97), .B2(new_n674), .ZN(new_n1029));
  NOR3_X1   g0829(.A1(new_n1027), .A2(new_n790), .A3(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n783), .B2(new_n918), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1013), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n940), .A2(new_n947), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n675), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1032), .B1(new_n1035), .B2(new_n948), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(G390));
  AOI21_X1  g0837(.A(new_n877), .B1(new_n883), .B2(new_n798), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n891), .B1(new_n1038), .B2(new_n893), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n717), .A2(new_n799), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n876), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n692), .A2(new_n667), .A3(new_n797), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n798), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n876), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n858), .A2(new_n863), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1046), .A2(new_n893), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1039), .A2(new_n1042), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n893), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n875), .B2(new_n877), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1051), .A2(new_n891), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n831), .A2(new_n836), .A3(G330), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1049), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n788), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n826), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n789), .B1(new_n1057), .B2(new_n334), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT114), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n205), .A2(new_n808), .B1(new_n741), .B2(new_n596), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT116), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n731), .A2(G68), .B1(new_n763), .B2(G87), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G97), .A2(new_n750), .B1(new_n744), .B2(G107), .ZN(new_n1063));
  AND4_X1   g0863(.A1(new_n387), .A2(new_n1061), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(new_n964), .B2(new_n754), .C1(new_n537), .C2(new_n728), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n808), .A2(new_n817), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n755), .A2(G128), .B1(G50), .B2(new_n731), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1067), .B1(new_n821), .B2(new_n741), .C1(new_n816), .C2(new_n745), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1066), .B(new_n1068), .C1(G125), .C2(new_n729), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(KEYINPUT54), .B(G143), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT115), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1069), .B(new_n263), .C1(new_n751), .C2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n763), .A2(G150), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT53), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1065), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT117), .Z(new_n1077));
  OAI21_X1  g0877(.A(new_n1059), .B1(new_n1077), .B2(new_n806), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT118), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n892), .B2(new_n778), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1078), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1081), .B1(KEYINPUT118), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1053), .B1(new_n1040), .B2(new_n876), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n884), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n831), .A2(G330), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(KEYINPUT112), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT112), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n831), .A2(new_n1089), .A3(G330), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1088), .A2(new_n800), .A3(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1091), .A2(KEYINPUT113), .A3(new_n877), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n1041), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1044), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n799), .B1(new_n1087), .B2(KEYINPUT112), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n876), .B1(new_n1095), .B2(new_n1090), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1094), .B1(new_n1096), .B2(KEYINPUT113), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1086), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n867), .A2(G330), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1099), .A2(new_n615), .A3(new_n870), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  AND3_X1   g0902(.A1(new_n1039), .A2(new_n1048), .A3(new_n1042), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1054), .B1(new_n1039), .B2(new_n1048), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n675), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT113), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n831), .A2(new_n1089), .A3(G330), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1089), .B1(new_n831), .B2(G330), .ZN(new_n1109));
  NOR3_X1   g0909(.A1(new_n1108), .A2(new_n1109), .A3(new_n799), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1107), .B1(new_n1110), .B2(new_n876), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1111), .A2(new_n1094), .A3(new_n1041), .A4(new_n1092), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1100), .B1(new_n1112), .B2(new_n1086), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1113), .A2(new_n1055), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1056), .B(new_n1084), .C1(new_n1106), .C2(new_n1114), .ZN(G378));
  INV_X1    g0915(.A(KEYINPUT121), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1100), .A2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1099), .A2(KEYINPUT121), .A3(new_n615), .A4(new_n870), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n1122), .B(KEYINPUT119), .Z(new_n1123));
  NAND2_X1  g0923(.A1(new_n434), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1123), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n429), .A2(new_n430), .A3(new_n433), .A4(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n426), .A2(new_n839), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1124), .A2(new_n426), .A3(new_n839), .A4(new_n1126), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n865), .B2(new_n645), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n837), .A2(new_n838), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n1134), .A2(new_n879), .A3(new_n857), .ZN(new_n1135));
  AND2_X1   g0935(.A1(new_n864), .A2(KEYINPUT40), .ZN(new_n1136));
  OAI211_X1 g0936(.A(G330), .B(new_n1133), .C1(new_n1135), .C2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1132), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n895), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n886), .A2(new_n1132), .A3(new_n1137), .A4(new_n894), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1121), .A2(KEYINPUT57), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT57), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1119), .B1(new_n1113), .B2(new_n1055), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1142), .A2(new_n1146), .A3(new_n675), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1139), .A2(new_n788), .A3(new_n1140), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n790), .B1(new_n202), .B2(new_n826), .ZN(new_n1149));
  INV_X1    g0949(.A(G124), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n260), .B1(new_n723), .B2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n808), .A2(new_n422), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n751), .A2(new_n816), .B1(new_n1072), .B2(new_n757), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1152), .B(new_n1153), .C1(G125), .C2(new_n755), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n761), .A2(G128), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1154), .B(new_n1155), .C1(new_n821), .C2(new_n745), .ZN(new_n1156));
  AOI211_X1 g0956(.A(G41), .B(new_n1151), .C1(new_n1156), .C2(KEYINPUT59), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1157), .B1(KEYINPUT59), .B2(new_n1156), .C1(new_n817), .C2(new_n730), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n202), .B1(new_n385), .B2(G41), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n751), .A2(new_n480), .B1(new_n205), .B2(new_n757), .ZN(new_n1160));
  AOI211_X1 g0960(.A(G41), .B(new_n1160), .C1(G116), .C2(new_n755), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n730), .A2(new_n225), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n745), .A2(new_n476), .B1(new_n216), .B2(new_n808), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1162), .B(new_n1163), .C1(G283), .C2(new_n729), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n761), .A2(G107), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1161), .A2(new_n1164), .A3(new_n387), .A4(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT58), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1158), .A2(new_n1159), .A3(new_n1167), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1149), .B1(new_n806), .B2(new_n1168), .C1(new_n1131), .C2(new_n778), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1148), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT120), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1148), .A2(KEYINPUT120), .A3(new_n1169), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1147), .A2(new_n1174), .ZN(G375));
  OAI211_X1 g0975(.A(new_n1086), .B(new_n1100), .C1(new_n1093), .C2(new_n1097), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1102), .A2(new_n926), .A3(new_n1176), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n755), .A2(G294), .B1(G77), .B2(new_n731), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n744), .A2(G116), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n763), .A2(G97), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1178), .A2(new_n1179), .A3(new_n992), .A4(new_n1180), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n387), .B1(new_n964), .B2(new_n741), .C1(new_n751), .C2(new_n212), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(G303), .C2(new_n729), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT122), .Z(new_n1184));
  AOI22_X1  g0984(.A1(new_n744), .A2(new_n1071), .B1(new_n761), .B2(G137), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n821), .B2(new_n754), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT123), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n263), .B1(new_n751), .B2(new_n422), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1162), .B(new_n1189), .C1(G159), .C2(new_n763), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n729), .A2(G128), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n736), .A2(G50), .ZN(new_n1192));
  OR2_X1    g0992(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1184), .B1(new_n1188), .B2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n790), .B1(new_n1195), .B2(new_n721), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n876), .B2(new_n778), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n216), .B2(new_n826), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n1098), .B2(new_n788), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1177), .A2(new_n1199), .ZN(G381));
  NOR2_X1   g1000(.A1(G375), .A2(G378), .ZN(new_n1201));
  INV_X1    g1001(.A(G384), .ZN(new_n1202));
  INV_X1    g1002(.A(G381), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n950), .A2(new_n1036), .A3(new_n976), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n1204), .A2(G396), .A3(G393), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .A4(new_n1205), .ZN(G407));
  INV_X1    g1006(.A(new_n1201), .ZN(new_n1207));
  OAI211_X1 g1007(.A(G407), .B(G213), .C1(G343), .C2(new_n1207), .ZN(G409));
  INV_X1    g1008(.A(KEYINPUT124), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT60), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1176), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1209), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1034), .B1(new_n1212), .B2(KEYINPUT60), .ZN(new_n1214));
  OAI211_X1 g1014(.A(KEYINPUT124), .B(new_n1176), .C1(new_n1113), .C2(new_n1210), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1216), .A2(G384), .A3(new_n1199), .ZN(new_n1217));
  AOI21_X1  g1017(.A(G384), .B1(new_n1216), .B2(new_n1199), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(G375), .A2(G378), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n650), .A2(G213), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n1144), .A2(new_n1145), .A3(new_n927), .ZN(new_n1222));
  OR3_X1    g1022(.A1(G378), .A2(new_n1222), .A3(new_n1170), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .A4(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(KEYINPUT63), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(G375), .A2(G378), .B1(G213), .B2(new_n650), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT63), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1226), .A2(new_n1227), .A3(new_n1219), .A4(new_n1223), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1225), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT125), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n650), .A2(G213), .A3(G2897), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1217), .A2(new_n1218), .A3(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1231), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1216), .A2(new_n1199), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n1202), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1216), .A2(G384), .A3(new_n1199), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1233), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1230), .B1(new_n1232), .B2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1220), .A2(new_n1221), .A3(new_n1223), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1231), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1235), .A2(new_n1236), .A3(new_n1233), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1240), .A2(new_n1241), .A3(KEYINPUT125), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1238), .A2(new_n1239), .A3(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT61), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(G393), .B(G396), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1204), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1036), .B1(new_n950), .B2(new_n976), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1245), .B1(new_n1248), .B2(KEYINPUT127), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(KEYINPUT126), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1247), .ZN(new_n1251));
  AND4_X1   g1051(.A1(KEYINPUT126), .A2(new_n1251), .A3(new_n1204), .A4(new_n1245), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT127), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(G387), .A2(new_n1253), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1249), .A2(new_n1250), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1229), .A2(new_n1243), .A3(new_n1244), .A4(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1224), .A2(KEYINPUT62), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1239), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT62), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1226), .A2(new_n1260), .A3(new_n1219), .A4(new_n1223), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1257), .A2(new_n1259), .A3(new_n1244), .A4(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1255), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1256), .A2(new_n1264), .ZN(G405));
  NAND2_X1  g1065(.A1(new_n1207), .A2(new_n1220), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1219), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1207), .B(new_n1220), .C1(new_n1218), .C2(new_n1217), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1255), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1255), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(G402));
endmodule


