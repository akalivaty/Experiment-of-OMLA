//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 0 0 0 1 1 1 1 0 1 0 0 0 1 1 0 0 0 0 0 1 1 0 0 0 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n561, new_n562, new_n564,
    new_n565, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n617, new_n619,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  AND2_X1   g033(.A1(G101), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(KEYINPUT64), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(new_n460), .A3(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n461), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n459), .B1(new_n466), .B2(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT65), .B1(new_n467), .B2(G2105), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT65), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  AOI211_X1 g046(.A(new_n471), .B(new_n461), .C1(new_n463), .C2(new_n465), .ZN(new_n472));
  OAI211_X1 g047(.A(new_n469), .B(new_n470), .C1(new_n472), .C2(new_n459), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n460), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G125), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n474), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  INV_X1    g058(.A(new_n466), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(new_n470), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n484), .A2(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  NOR2_X1   g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(new_n470), .B2(G112), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n486), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  NAND2_X1  g067(.A1(new_n463), .A2(new_n465), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n493), .A2(G138), .A3(new_n470), .A4(new_n476), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT66), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n496), .A2(new_n497), .A3(new_n470), .A4(G138), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n498), .B1(new_n496), .B2(new_n497), .ZN(new_n499));
  INV_X1    g074(.A(new_n478), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n493), .A2(G126), .A3(G2105), .A4(new_n476), .ZN(new_n503));
  OR2_X1    g078(.A1(G102), .A2(G2105), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n504), .B(G2104), .C1(G114), .C2(new_n470), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n502), .A2(KEYINPUT67), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT67), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n494), .A2(KEYINPUT4), .B1(new_n500), .B2(new_n499), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(new_n506), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(KEYINPUT68), .A3(G62), .ZN(new_n519));
  NAND2_X1  g094(.A1(G75), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT68), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n515), .A2(new_n517), .ZN(new_n522));
  INV_X1    g097(.A(G62), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n519), .A2(new_n520), .A3(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n525), .A2(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT6), .B(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n518), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G88), .ZN(new_n529));
  INV_X1    g104(.A(G50), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n527), .A2(G543), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n528), .A2(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g107(.A(KEYINPUT69), .B1(new_n526), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n532), .B1(G651), .B2(new_n525), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT69), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n533), .A2(new_n536), .ZN(G166));
  NAND3_X1  g112(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  INV_X1    g115(.A(G89), .ZN(new_n541));
  OAI211_X1 g116(.A(new_n538), .B(new_n540), .C1(new_n528), .C2(new_n541), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n531), .A2(KEYINPUT70), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n531), .A2(KEYINPUT70), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n542), .B1(new_n545), .B2(G51), .ZN(G168));
  XOR2_X1   g121(.A(KEYINPUT71), .B(G52), .Z(new_n547));
  AOI21_X1  g122(.A(new_n547), .B1(new_n543), .B2(new_n544), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G651), .ZN(new_n550));
  INV_X1    g125(.A(G90), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n549), .A2(new_n550), .B1(new_n551), .B2(new_n528), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n548), .A2(new_n552), .ZN(G171));
  AOI22_X1  g128(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT72), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G651), .ZN(new_n556));
  INV_X1    g131(.A(new_n528), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n545), .A2(G43), .B1(G81), .B2(new_n557), .ZN(new_n558));
  AND2_X1   g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(new_n562));
  XOR2_X1   g137(.A(new_n562), .B(KEYINPUT73), .Z(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n561), .A2(new_n565), .ZN(G188));
  AND2_X1   g141(.A1(new_n527), .A2(G543), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G53), .ZN(new_n568));
  XOR2_X1   g143(.A(new_n568), .B(KEYINPUT9), .Z(new_n569));
  AOI22_X1  g144(.A1(new_n518), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G91), .ZN(new_n571));
  OAI22_X1  g146(.A1(new_n570), .A2(new_n550), .B1(new_n571), .B2(new_n528), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n569), .A2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  INV_X1    g149(.A(G168), .ZN(G286));
  XNOR2_X1  g150(.A(new_n534), .B(KEYINPUT69), .ZN(G303));
  INV_X1    g151(.A(G87), .ZN(new_n577));
  OR3_X1    g152(.A1(new_n528), .A2(KEYINPUT74), .A3(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(G74), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n550), .B1(new_n522), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n580), .B1(G49), .B2(new_n567), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT74), .B1(new_n528), .B2(new_n577), .ZN(new_n582));
  AND3_X1   g157(.A1(new_n578), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G288));
  INV_X1    g159(.A(G86), .ZN(new_n585));
  INV_X1    g160(.A(G48), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n528), .A2(new_n585), .B1(new_n586), .B2(new_n531), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n518), .A2(G61), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n550), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n588), .A2(new_n592), .ZN(G305));
  AOI22_X1  g168(.A1(new_n545), .A2(G47), .B1(G85), .B2(new_n557), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n595), .A2(KEYINPUT75), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(KEYINPUT75), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n596), .A2(G651), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n594), .A2(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  AND3_X1   g175(.A1(new_n518), .A2(G92), .A3(new_n527), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT10), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n545), .A2(G54), .ZN(new_n603));
  OR2_X1    g178(.A1(KEYINPUT76), .A2(G66), .ZN(new_n604));
  NAND2_X1  g179(.A1(KEYINPUT76), .A2(G66), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n518), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G79), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(new_n514), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G651), .ZN(new_n609));
  AND3_X1   g184(.A1(new_n602), .A2(new_n603), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n600), .B1(G868), .B2(new_n610), .ZN(G284));
  OAI21_X1  g186(.A(new_n600), .B1(G868), .B2(new_n610), .ZN(G321));
  NAND2_X1  g187(.A1(G286), .A2(G868), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n569), .A2(new_n572), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(G297));
  OAI21_X1  g190(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n610), .B1(new_n617), .B2(G860), .ZN(G148));
  OAI21_X1  g193(.A(KEYINPUT77), .B1(new_n559), .B2(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n610), .A2(new_n617), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  MUX2_X1   g196(.A(KEYINPUT77), .B(new_n619), .S(new_n621), .Z(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n485), .A2(G123), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n487), .A2(G135), .ZN(new_n625));
  NOR2_X1   g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  OAI21_X1  g201(.A(G2104), .B1(new_n470), .B2(G111), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n624), .B(new_n625), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(G2096), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n470), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  INV_X1    g208(.A(G2100), .ZN(new_n634));
  AND2_X1   g209(.A1(new_n634), .A2(KEYINPUT78), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n634), .A2(KEYINPUT78), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n630), .B(new_n637), .C1(new_n635), .C2(new_n633), .ZN(G156));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2435), .ZN(new_n640));
  XOR2_X1   g215(.A(G2427), .B(G2438), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(KEYINPUT14), .ZN(new_n643));
  XOR2_X1   g218(.A(G2451), .B(G2454), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G1341), .B(G1348), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n648), .B(new_n649), .Z(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(G14), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(G401));
  XNOR2_X1  g227(.A(G2084), .B(G2090), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT79), .Z(new_n654));
  XOR2_X1   g229(.A(G2072), .B(G2078), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT17), .ZN(new_n656));
  XOR2_X1   g231(.A(G2067), .B(G2678), .Z(new_n657));
  OAI21_X1  g232(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n657), .B2(new_n655), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT80), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n654), .A2(new_n657), .A3(new_n655), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT18), .ZN(new_n662));
  INV_X1    g237(.A(new_n654), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n663), .A2(new_n656), .A3(new_n657), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n660), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(new_n629), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(new_n634), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G227));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT81), .ZN(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  AND2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G1971), .B(G1976), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT20), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n670), .A2(new_n671), .ZN(new_n677));
  AOI22_X1  g252(.A1(new_n675), .A2(new_n676), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  OR3_X1    g253(.A1(new_n672), .A2(new_n677), .A3(new_n674), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n678), .B(new_n679), .C1(new_n676), .C2(new_n675), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT21), .B(G1986), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G1991), .B(G1996), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT82), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n682), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT22), .B(G1981), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n685), .B(new_n686), .Z(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(G229));
  XOR2_X1   g263(.A(KEYINPUT95), .B(KEYINPUT96), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT23), .ZN(new_n690));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G20), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n690), .B(new_n692), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(new_n614), .B2(new_n691), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(G1956), .Z(new_n695));
  INV_X1    g270(.A(G2090), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT83), .B(G29), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G35), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G162), .B2(new_n698), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n695), .B1(new_n696), .B2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT97), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OR2_X1    g281(.A1(G29), .A2(G33), .ZN(new_n707));
  NAND2_X1  g282(.A1(G115), .A2(G2104), .ZN(new_n708));
  INV_X1    g283(.A(G127), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n478), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G2105), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT89), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n487), .A2(G139), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT25), .Z(new_n715));
  NAND3_X1  g290(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n707), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G2072), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT30), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n717), .B1(new_n722), .B2(G28), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT92), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n722), .A2(G28), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n723), .A2(new_n724), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n718), .B2(new_n719), .ZN(new_n729));
  NOR2_X1   g304(.A1(G5), .A2(G16), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G171), .B2(G16), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n731), .A2(G1961), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n628), .A2(new_n698), .ZN(new_n733));
  NOR4_X1   g308(.A1(new_n721), .A2(new_n729), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT84), .ZN(new_n735));
  INV_X1    g310(.A(G25), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n697), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n697), .A2(new_n736), .ZN(new_n738));
  AOI22_X1  g313(.A1(G119), .A2(new_n485), .B1(new_n487), .B2(G131), .ZN(new_n739));
  OR2_X1    g314(.A1(G95), .A2(G2105), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n740), .B(G2104), .C1(G107), .C2(new_n470), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT85), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n738), .B1(new_n743), .B2(new_n697), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n737), .B1(new_n744), .B2(new_n735), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT35), .B(G1991), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G290), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G16), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n749), .B(G1986), .C1(G16), .C2(G24), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n749), .B1(G16), .B2(G24), .ZN(new_n751));
  INV_X1    g326(.A(G1986), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n745), .A2(new_n746), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n747), .A2(new_n750), .A3(new_n753), .A4(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G1971), .ZN(new_n756));
  NOR2_X1   g331(.A1(G16), .A2(G22), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n756), .B(new_n758), .C1(G303), .C2(new_n691), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n691), .B1(new_n533), .B2(new_n536), .ZN(new_n760));
  OAI21_X1  g335(.A(G1971), .B1(new_n760), .B2(new_n757), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n583), .A2(G16), .ZN(new_n763));
  OR2_X1    g338(.A1(G16), .A2(G23), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT33), .B(G1976), .Z(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  MUX2_X1   g342(.A(G6), .B(G305), .S(G16), .Z(new_n768));
  XOR2_X1   g343(.A(KEYINPUT32), .B(G1981), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n762), .A2(new_n767), .A3(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT34), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n762), .A2(new_n767), .A3(KEYINPUT34), .A4(new_n770), .ZN(new_n774));
  AOI211_X1 g349(.A(KEYINPUT36), .B(new_n755), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT36), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n773), .A2(new_n774), .ZN(new_n777));
  INV_X1    g352(.A(new_n755), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n706), .B(new_n734), .C1(new_n775), .C2(new_n779), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n698), .A2(KEYINPUT93), .A3(G27), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G164), .B2(new_n698), .ZN(new_n782));
  AOI21_X1  g357(.A(KEYINPUT93), .B1(new_n698), .B2(G27), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n784), .A2(G2078), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT24), .B(G34), .Z(new_n786));
  OAI22_X1  g361(.A1(new_n482), .A2(new_n717), .B1(new_n697), .B2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(G2084), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n785), .B(new_n789), .C1(G2090), .C2(new_n702), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n704), .A2(new_n705), .ZN(new_n791));
  NOR2_X1   g366(.A1(G168), .A2(new_n691), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n691), .B2(G21), .ZN(new_n793));
  INV_X1    g368(.A(G1966), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  INV_X1    g371(.A(G1961), .ZN(new_n797));
  INV_X1    g372(.A(new_n731), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n795), .B(new_n796), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  NOR4_X1   g374(.A1(new_n780), .A2(new_n790), .A3(new_n791), .A4(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(G29), .A2(G32), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n487), .A2(G141), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n485), .A2(G129), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n470), .A2(G105), .A3(G2104), .ZN(new_n804));
  NAND3_X1  g379(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT26), .Z(new_n806));
  NAND4_X1  g381(.A1(new_n802), .A2(new_n803), .A3(new_n804), .A4(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT91), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n801), .B1(new_n809), .B2(G29), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT27), .B(G1996), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n787), .A2(new_n788), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT90), .Z(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n784), .A2(G2078), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT31), .B(G11), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n800), .A2(new_n812), .A3(new_n815), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n691), .A2(G19), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n559), .B2(new_n691), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(G1341), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n698), .A2(G26), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n485), .A2(G128), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n487), .A2(G140), .ZN(new_n828));
  NOR2_X1   g403(.A1(G104), .A2(G2105), .ZN(new_n829));
  OAI21_X1  g404(.A(G2104), .B1(new_n470), .B2(G116), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n827), .B(new_n828), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  AND3_X1   g406(.A1(new_n831), .A2(KEYINPUT86), .A3(G29), .ZN(new_n832));
  AOI21_X1  g407(.A(KEYINPUT86), .B1(new_n831), .B2(G29), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n826), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(G2067), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n691), .A2(G4), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n610), .B2(new_n691), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(G1348), .Z(new_n839));
  NAND3_X1  g414(.A1(new_n823), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT88), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n820), .A2(new_n841), .ZN(G311));
  INV_X1    g417(.A(KEYINPUT98), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n820), .B2(new_n841), .ZN(new_n844));
  INV_X1    g419(.A(new_n734), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n777), .A2(new_n778), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(KEYINPUT36), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n777), .A2(new_n776), .A3(new_n778), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n791), .ZN(new_n850));
  INV_X1    g425(.A(new_n799), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n849), .A2(new_n850), .A3(new_n851), .A4(new_n706), .ZN(new_n852));
  NOR4_X1   g427(.A1(new_n852), .A2(new_n814), .A3(new_n818), .A4(new_n790), .ZN(new_n853));
  INV_X1    g428(.A(new_n841), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n853), .A2(KEYINPUT98), .A3(new_n854), .A4(new_n812), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n844), .A2(new_n855), .ZN(G150));
  AND2_X1   g431(.A1(new_n545), .A2(G55), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n858));
  INV_X1    g433(.A(G93), .ZN(new_n859));
  OAI22_X1  g434(.A1(new_n858), .A2(new_n550), .B1(new_n859), .B2(new_n528), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(G860), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT37), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n861), .A2(KEYINPUT99), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n865), .A2(new_n559), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n861), .A2(KEYINPUT99), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n559), .A2(KEYINPUT99), .A3(new_n861), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT38), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n610), .A2(G559), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT39), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(KEYINPUT100), .Z(new_n876));
  OAI21_X1  g451(.A(new_n862), .B1(new_n873), .B2(new_n874), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n864), .B1(new_n876), .B2(new_n877), .ZN(G145));
  MUX2_X1   g453(.A(new_n809), .B(new_n807), .S(new_n716), .Z(new_n879));
  INV_X1    g454(.A(KEYINPUT102), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n506), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n503), .A2(KEYINPUT102), .A3(new_n505), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n510), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n831), .B(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n879), .B(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n743), .B(new_n632), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n487), .A2(G142), .ZN(new_n887));
  NOR2_X1   g462(.A1(G106), .A2(G2105), .ZN(new_n888));
  OAI21_X1  g463(.A(G2104), .B1(new_n470), .B2(G118), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n890), .B1(G130), .B2(new_n485), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n886), .B(new_n891), .Z(new_n892));
  XNOR2_X1  g467(.A(new_n885), .B(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n482), .B(KEYINPUT101), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(G162), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n628), .ZN(new_n896));
  OR3_X1    g471(.A1(new_n893), .A2(KEYINPUT103), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(G37), .B1(new_n893), .B2(new_n896), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT103), .B1(new_n893), .B2(new_n896), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g476(.A(new_n583), .B(G305), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(G303), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(new_n748), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n868), .A2(new_n620), .A3(new_n869), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n620), .B1(new_n868), .B2(new_n869), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT104), .ZN(new_n909));
  NAND2_X1  g484(.A1(G299), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n610), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n614), .A2(KEYINPUT104), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n614), .A2(new_n610), .A3(KEYINPUT104), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n908), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT42), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n913), .A2(KEYINPUT41), .A3(new_n914), .ZN(new_n918));
  AOI21_X1  g493(.A(KEYINPUT41), .B1(new_n913), .B2(new_n914), .ZN(new_n919));
  OAI22_X1  g494(.A1(new_n906), .A2(new_n907), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n916), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n917), .B1(new_n916), .B2(new_n920), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n905), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n923), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n925), .A2(new_n921), .A3(new_n904), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n924), .A2(new_n926), .A3(G868), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n861), .A2(G868), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n924), .A2(new_n926), .A3(KEYINPUT105), .A4(G868), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n930), .A2(KEYINPUT106), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT106), .B1(new_n930), .B2(new_n931), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(G295));
  AND2_X1   g509(.A1(new_n930), .A2(new_n931), .ZN(G331));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n936));
  INV_X1    g511(.A(G37), .ZN(new_n937));
  XNOR2_X1  g512(.A(G171), .B(G168), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n870), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n940));
  INV_X1    g515(.A(new_n938), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n868), .A2(new_n869), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n939), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n918), .A2(new_n919), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n870), .A2(KEYINPUT107), .A3(new_n938), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n939), .A2(new_n914), .A3(new_n913), .A4(new_n942), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n936), .B(new_n937), .C1(new_n948), .C2(new_n904), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n946), .A2(new_n904), .A3(new_n947), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT109), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n946), .A2(new_n952), .A3(new_n904), .A4(new_n947), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n904), .B1(new_n946), .B2(new_n947), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT108), .B1(new_n955), .B2(G37), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n949), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n943), .A2(new_n945), .ZN(new_n960));
  INV_X1    g535(.A(new_n944), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n939), .A2(new_n942), .ZN(new_n962));
  OAI22_X1  g537(.A1(new_n960), .A2(new_n915), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n905), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n954), .A2(new_n937), .A3(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n965), .A2(new_n958), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT44), .B1(new_n959), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n958), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n949), .A2(new_n954), .A3(KEYINPUT43), .A4(new_n956), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n967), .A2(new_n971), .ZN(G397));
  INV_X1    g547(.A(G40), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n973), .B1(new_n480), .B2(G2105), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n468), .A2(new_n473), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n468), .A2(new_n473), .A3(KEYINPUT111), .A4(new_n974), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G2078), .ZN(new_n980));
  INV_X1    g555(.A(G1384), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n508), .A2(new_n511), .A3(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n882), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT102), .B1(new_n503), .B2(new_n505), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n502), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n987), .A2(KEYINPUT45), .A3(new_n981), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n979), .A2(new_n980), .A3(new_n984), .A4(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT53), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT121), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n977), .A2(new_n978), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT45), .B1(new_n987), .B2(new_n981), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT115), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n982), .A2(new_n983), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(new_n883), .B2(G1384), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT115), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n999), .A2(new_n1000), .A3(new_n977), .A4(new_n978), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n990), .A2(G2078), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n996), .A2(new_n997), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n982), .A2(KEYINPUT50), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n881), .A2(new_n882), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1384), .B1(new_n1005), .B2(new_n502), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n979), .A2(new_n1004), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n797), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n989), .A2(KEYINPUT121), .A3(new_n990), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n993), .A2(new_n1003), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT122), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n1012), .A2(new_n1013), .A3(G171), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1013), .B1(new_n1012), .B2(G171), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1006), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n983), .ZN(new_n1018));
  INV_X1    g593(.A(new_n975), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1018), .A2(new_n1019), .A3(new_n988), .A4(new_n1002), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n993), .A2(new_n1010), .A3(new_n1011), .A4(new_n1020), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n1021), .A2(G171), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT54), .B1(new_n1016), .B2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n996), .A2(new_n997), .A3(new_n1001), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n979), .A2(new_n1004), .A3(new_n1008), .ZN(new_n1025));
  AOI22_X1  g600(.A1(new_n1024), .A2(new_n794), .B1(new_n1025), .B2(new_n788), .ZN(new_n1026));
  INV_X1    g601(.A(G8), .ZN(new_n1027));
  OR3_X1    g602(.A1(new_n1026), .A2(new_n1027), .A3(G168), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1024), .A2(new_n794), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1025), .A2(new_n788), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1029), .A2(G168), .A3(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1027), .A2(KEYINPUT120), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1031), .A2(KEYINPUT51), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT51), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1028), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n984), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n988), .A2(new_n977), .A3(new_n978), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n756), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n979), .A2(new_n696), .A3(new_n1004), .A4(new_n1008), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1041), .B1(G303), .B2(G8), .ZN(new_n1042));
  NOR3_X1   g617(.A1(G166), .A2(KEYINPUT55), .A3(new_n1027), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1040), .A2(G8), .A3(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1006), .A2(new_n977), .A3(new_n978), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n583), .A2(G1976), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1046), .A2(G8), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT52), .ZN(new_n1049));
  INV_X1    g624(.A(G1981), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n588), .A2(new_n592), .A3(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(G1981), .B1(new_n587), .B2(new_n591), .ZN(new_n1052));
  OR2_X1    g627(.A1(KEYINPUT113), .A2(KEYINPUT49), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1053), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(G8), .A3(new_n1046), .ZN(new_n1057));
  INV_X1    g632(.A(G1976), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT52), .B1(G288), .B2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1059), .A2(new_n1046), .A3(G8), .A4(new_n1047), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1049), .A2(new_n1057), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1045), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1007), .B1(new_n987), .B2(new_n981), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n994), .A2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n508), .A2(new_n511), .A3(new_n1007), .A4(new_n981), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT114), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1064), .B(new_n696), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n1038), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1044), .B1(new_n1071), .B2(G8), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT123), .B1(new_n1062), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1044), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n977), .B(new_n978), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n512), .A2(KEYINPUT114), .A3(new_n1007), .A4(new_n981), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1075), .B1(new_n1067), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n979), .A2(new_n984), .A3(new_n988), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n1077), .A2(new_n696), .B1(new_n756), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1074), .B1(new_n1079), .B2(new_n1027), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1049), .A2(new_n1057), .A3(new_n1060), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1027), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1081), .B1(new_n1044), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT123), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1080), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1073), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1011), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT121), .B1(new_n989), .B2(new_n990), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1089), .A2(G301), .A3(new_n1003), .A4(new_n1010), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1021), .A2(G171), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1090), .A2(new_n1091), .A3(KEYINPUT54), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1035), .A2(new_n1086), .A3(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT124), .B1(new_n1023), .B2(new_n1093), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1035), .A2(new_n1086), .A3(new_n1092), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT124), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1012), .A2(G171), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT122), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1012), .A2(new_n1013), .A3(G171), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1098), .A2(new_n1099), .A3(new_n1022), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1095), .A2(new_n1096), .A3(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT56), .B(G2072), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  OAI22_X1  g680(.A1(new_n1077), .A2(G1956), .B1(new_n1078), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(new_n572), .B2(KEYINPUT116), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1108), .B(KEYINPUT117), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1109), .B(G299), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1106), .A2(new_n1111), .ZN(new_n1112));
  OAI22_X1  g687(.A1(new_n1025), .A2(G1348), .B1(G2067), .B2(new_n1046), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n610), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1114), .B(KEYINPUT118), .ZN(new_n1115));
  OAI221_X1 g690(.A(new_n1110), .B1(new_n1078), .B2(new_n1105), .C1(G1956), .C2(new_n1077), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT61), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1113), .A2(KEYINPUT60), .A3(new_n911), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1116), .A2(KEYINPUT61), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1046), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT58), .B(G1341), .ZN(new_n1124));
  OAI22_X1  g699(.A1(new_n1078), .A2(G1996), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1125), .A2(new_n559), .ZN(new_n1126));
  OR2_X1    g701(.A1(new_n1126), .A2(KEYINPUT59), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(KEYINPUT59), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1121), .A2(new_n1122), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT60), .ZN(new_n1130));
  OR2_X1    g705(.A1(new_n1113), .A2(new_n610), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1130), .B1(new_n1131), .B2(new_n1114), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1112), .B(new_n1117), .C1(new_n1129), .C2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1094), .A2(new_n1103), .A3(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1045), .A2(new_n1081), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1057), .A2(new_n1058), .A3(new_n583), .ZN(new_n1136));
  AOI211_X1 g711(.A(new_n1027), .B(new_n1123), .C1(new_n1136), .C2(new_n1051), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1026), .A2(new_n1027), .A3(G286), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1138), .A2(new_n1080), .A3(new_n1083), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT63), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1082), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1140), .B1(new_n1142), .B2(new_n1074), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1143), .A2(new_n1138), .A3(new_n1083), .ZN(new_n1144));
  AOI211_X1 g719(.A(new_n1135), .B(new_n1137), .C1(new_n1141), .C2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1146), .B(new_n1028), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1147), .A2(new_n1148), .A3(new_n1086), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(KEYINPUT125), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT125), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1147), .A2(new_n1148), .A3(new_n1151), .A4(new_n1086), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1035), .A2(KEYINPUT62), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT126), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1035), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1150), .A2(new_n1152), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1134), .A2(new_n1145), .A3(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n743), .B(new_n746), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n1159), .B(KEYINPUT112), .Z(new_n1160));
  XNOR2_X1  g735(.A(new_n831), .B(new_n835), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n807), .A2(G1996), .ZN(new_n1162));
  INV_X1    g737(.A(new_n809), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1161), .B(new_n1162), .C1(new_n1163), .C2(G1996), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1160), .A2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(G290), .B(new_n752), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1018), .A2(new_n994), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1158), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1168), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT46), .ZN(new_n1172));
  OR3_X1    g747(.A1(new_n1171), .A2(new_n1172), .A3(G1996), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1161), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1168), .B1(new_n807), .B2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1172), .B1(new_n1171), .B2(G1996), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1173), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT47), .ZN(new_n1178));
  NOR3_X1   g753(.A1(new_n1164), .A2(new_n746), .A3(new_n743), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n831), .A2(G2067), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1168), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1168), .A2(new_n752), .A3(new_n748), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1182), .B(KEYINPUT48), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1183), .B1(new_n1165), .B2(new_n1171), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1178), .A2(new_n1181), .A3(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1185), .B(KEYINPUT127), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1170), .A2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g762(.A1(new_n968), .A2(G319), .A3(new_n651), .A4(new_n970), .ZN(new_n1189));
  NAND3_X1  g763(.A1(new_n900), .A2(new_n667), .A3(new_n687), .ZN(new_n1190));
  NOR2_X1   g764(.A1(new_n1189), .A2(new_n1190), .ZN(G308));
  OR2_X1    g765(.A1(new_n1189), .A2(new_n1190), .ZN(G225));
endmodule


