//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 1 1 1 0 1 0 1 1 0 0 0 0 0 1 1 0 0 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n815, new_n816, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT89), .ZN(new_n203));
  OR3_X1    g002(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT15), .ZN(new_n204));
  INV_X1    g003(.A(G29gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n205), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n206));
  AND2_X1   g005(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n206), .B1(new_n209), .B2(G36gat), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT15), .B1(new_n202), .B2(new_n203), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n204), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT90), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n214), .B1(new_n210), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G8gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(G15gat), .B(G22gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT91), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n218), .B(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G1gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT16), .ZN(new_n222));
  XOR2_X1   g021(.A(new_n222), .B(KEYINPUT92), .Z(new_n223));
  NAND2_X1  g022(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n217), .B1(new_n224), .B2(KEYINPUT93), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n224), .B1(G1gat), .B2(new_n220), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI221_X1 g026(.A(new_n224), .B1(KEYINPUT93), .B2(new_n217), .C1(G1gat), .C2(new_n220), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n216), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n230), .B(KEYINPUT94), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n216), .B(KEYINPUT17), .ZN(new_n232));
  INV_X1    g031(.A(new_n229), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n231), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT18), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n231), .B1(new_n229), .B2(new_n216), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n235), .B(KEYINPUT13), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n231), .A2(new_n234), .A3(KEYINPUT18), .A4(new_n235), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n238), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G113gat), .B(G141gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(G197gat), .ZN(new_n245));
  XOR2_X1   g044(.A(KEYINPUT11), .B(G169gat), .Z(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n247), .B(KEYINPUT12), .Z(new_n248));
  NAND2_X1  g047(.A1(new_n243), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n248), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n238), .A2(new_n241), .A3(new_n250), .A4(new_n242), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(G8gat), .B(G36gat), .Z(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(KEYINPUT78), .ZN(new_n255));
  XNOR2_X1  g054(.A(G64gat), .B(G92gat), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n255), .B(new_n256), .Z(new_n257));
  INV_X1    g056(.A(KEYINPUT24), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n258), .A2(G183gat), .A3(G190gat), .ZN(new_n259));
  AND2_X1   g058(.A1(G183gat), .A2(G190gat), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n259), .B1(new_n260), .B2(new_n258), .ZN(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT67), .B(G190gat), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n261), .B1(G183gat), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT23), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n264), .B1(G169gat), .B2(G176gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(KEYINPUT65), .ZN(new_n266));
  INV_X1    g065(.A(G169gat), .ZN(new_n267));
  INV_X1    g066(.A(G176gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n269), .A2(new_n264), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n267), .A2(new_n268), .ZN(new_n271));
  OAI21_X1  g070(.A(KEYINPUT66), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n273));
  NAND2_X1  g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n273), .B(new_n274), .C1(new_n269), .C2(new_n264), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n263), .A2(new_n266), .A3(new_n272), .A4(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT25), .ZN(new_n277));
  XOR2_X1   g076(.A(KEYINPUT64), .B(G169gat), .Z(new_n278));
  NOR2_X1   g077(.A1(new_n264), .A2(G176gat), .ZN(new_n279));
  AOI211_X1 g078(.A(KEYINPUT25), .B(new_n271), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n261), .B1(G183gat), .B2(G190gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n280), .A2(new_n266), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n271), .B1(KEYINPUT26), .B2(new_n269), .ZN(new_n283));
  OR2_X1    g082(.A1(new_n269), .A2(KEYINPUT26), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n260), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n262), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT27), .B(G183gat), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n286), .A2(KEYINPUT28), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT28), .B1(new_n286), .B2(new_n287), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n285), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n277), .A2(new_n282), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G226gat), .A2(G233gat), .ZN(new_n292));
  XOR2_X1   g091(.A(new_n292), .B(KEYINPUT76), .Z(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT29), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n293), .B1(new_n291), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G211gat), .B(G218gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT22), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT74), .B(G218gat), .ZN(new_n303));
  INV_X1    g102(.A(G211gat), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT75), .ZN(new_n306));
  XNOR2_X1  g105(.A(G197gat), .B(G204gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n306), .B1(new_n305), .B2(new_n307), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n301), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n305), .A2(new_n307), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT75), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n313), .A2(new_n308), .A3(new_n300), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n315), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT77), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n294), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n317), .B(new_n319), .C1(new_n298), .C2(new_n318), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n257), .B1(new_n321), .B2(KEYINPUT37), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT37), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n323), .B1(new_n299), .B2(new_n317), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n315), .B(new_n319), .C1(new_n298), .C2(new_n318), .ZN(new_n325));
  AND2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OR3_X1    g125(.A1(new_n322), .A2(KEYINPUT38), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n323), .B1(new_n320), .B2(new_n316), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT38), .B1(new_n322), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n257), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n316), .A2(new_n320), .A3(new_n330), .ZN(new_n331));
  AND3_X1   g130(.A1(new_n327), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G127gat), .B(G134gat), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT1), .ZN(new_n334));
  INV_X1    g133(.A(G120gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G113gat), .ZN(new_n336));
  INV_X1    g135(.A(G113gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(G120gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n333), .B1(new_n334), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n335), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n334), .B(new_n341), .C1(new_n339), .C2(KEYINPUT68), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n333), .B(KEYINPUT69), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n340), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT79), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n346), .B1(G155gat), .B2(G162gat), .ZN(new_n347));
  INV_X1    g146(.A(G141gat), .ZN(new_n348));
  INV_X1    g147(.A(G148gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G141gat), .A2(G148gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT2), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n353), .B1(G155gat), .B2(G162gat), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n347), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G155gat), .B(G162gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(G155gat), .ZN(new_n359));
  INV_X1    g158(.A(G162gat), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT2), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n361), .A2(new_n350), .A3(new_n351), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n362), .A2(new_n356), .A3(new_n347), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n345), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n340), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT69), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n333), .B(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n366), .B1(new_n368), .B2(new_n342), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n355), .A2(new_n357), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n356), .B1(new_n362), .B2(new_n347), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n365), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G225gat), .A2(G233gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n375), .B(KEYINPUT80), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT5), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n379), .B1(new_n370), .B2(new_n371), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n358), .A2(KEYINPUT3), .A3(new_n363), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(new_n369), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n376), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT82), .ZN(new_n385));
  XOR2_X1   g184(.A(KEYINPUT81), .B(KEYINPUT4), .Z(new_n386));
  OAI21_X1  g185(.A(new_n386), .B1(new_n369), .B2(new_n372), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n345), .A2(KEYINPUT4), .A3(new_n364), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n384), .A2(new_n385), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n387), .A2(new_n382), .A3(new_n388), .A4(new_n383), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT82), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n378), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  OR2_X1    g191(.A1(new_n365), .A2(new_n386), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT5), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT4), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n365), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n384), .A2(new_n393), .A3(new_n394), .A4(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n392), .A2(new_n398), .ZN(new_n399));
  XOR2_X1   g198(.A(G1gat), .B(G29gat), .Z(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G57gat), .B(G85gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT6), .B1(new_n399), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n378), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n390), .A2(KEYINPUT82), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n390), .A2(KEYINPUT82), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n397), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT87), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n404), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT88), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n410), .A2(KEYINPUT87), .A3(new_n397), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n412), .B1(new_n392), .B2(new_n398), .ZN(new_n417));
  INV_X1    g216(.A(new_n404), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n415), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT88), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n406), .B1(new_n416), .B2(new_n420), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n399), .A2(new_n404), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT6), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n332), .A2(new_n425), .ZN(new_n426));
  OR3_X1    g225(.A1(new_n321), .A2(KEYINPUT30), .A3(new_n257), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n393), .A2(new_n382), .A3(new_n396), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n376), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n429), .B(KEYINPUT39), .C1(new_n376), .C2(new_n374), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n430), .B(new_n404), .C1(KEYINPUT39), .C2(new_n429), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT40), .ZN(new_n432));
  OR2_X1    g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n321), .A2(new_n257), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n434), .A2(KEYINPUT30), .A3(new_n331), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n431), .A2(new_n432), .ZN(new_n436));
  AND4_X1   g235(.A1(new_n427), .A2(new_n433), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n416), .A2(new_n420), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n380), .A2(new_n296), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n315), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n440), .A2(G228gat), .A3(G233gat), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n311), .A2(new_n296), .A3(new_n314), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT3), .B1(new_n442), .B2(KEYINPUT86), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n443), .B1(KEYINPUT86), .B2(new_n442), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n441), .B1(new_n444), .B2(new_n372), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT84), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n440), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n315), .A2(KEYINPUT84), .A3(new_n439), .ZN(new_n449));
  AND2_X1   g248(.A1(new_n442), .A2(new_n379), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n448), .B(new_n449), .C1(new_n450), .C2(new_n364), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT85), .ZN(new_n452));
  NAND2_X1  g251(.A1(G228gat), .A2(G233gat), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n452), .B1(new_n451), .B2(new_n453), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n446), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(G22gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n448), .A2(new_n449), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n364), .B1(new_n442), .B2(new_n379), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n453), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT85), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n454), .ZN(new_n463));
  INV_X1    g262(.A(G22gat), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n463), .A2(new_n464), .A3(new_n446), .ZN(new_n465));
  XNOR2_X1  g264(.A(G78gat), .B(G106gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(KEYINPUT31), .B(G50gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n466), .B(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n458), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n468), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n464), .B1(new_n463), .B2(new_n446), .ZN(new_n471));
  AOI211_X1 g270(.A(G22gat), .B(new_n445), .C1(new_n462), .C2(new_n454), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n437), .A2(new_n438), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n426), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n435), .A2(new_n427), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n411), .A2(new_n418), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n405), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n423), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n480), .A2(new_n469), .A3(new_n473), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n282), .A2(new_n290), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT70), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n482), .A2(new_n483), .A3(new_n369), .A4(new_n277), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n345), .A2(KEYINPUT70), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n369), .A2(new_n483), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n291), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(G227gat), .A2(G233gat), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT72), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT34), .ZN(new_n491));
  OR2_X1    g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n491), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n484), .A2(new_n487), .A3(G227gat), .A4(G233gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT32), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT33), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(KEYINPUT71), .B(G71gat), .ZN(new_n499));
  INV_X1    g298(.A(G99gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  XOR2_X1   g300(.A(G15gat), .B(G43gat), .Z(new_n502));
  XOR2_X1   g301(.A(new_n501), .B(new_n502), .Z(new_n503));
  NAND3_X1  g302(.A1(new_n496), .A2(new_n498), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n503), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n495), .B(KEYINPUT32), .C1(new_n497), .C2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n494), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n492), .A2(new_n504), .A3(new_n493), .A4(new_n506), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n508), .A2(KEYINPUT73), .A3(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT36), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n475), .A2(new_n481), .A3(new_n511), .ZN(new_n512));
  AOI22_X1  g311(.A1(new_n435), .A2(new_n427), .B1(new_n478), .B2(new_n423), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n508), .A2(new_n509), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n471), .A2(new_n472), .A3(new_n470), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n468), .B1(new_n458), .B2(new_n465), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n513), .B(new_n514), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT35), .ZN(new_n518));
  INV_X1    g317(.A(new_n514), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n519), .B1(new_n473), .B2(new_n469), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n414), .B1(new_n413), .B2(new_n415), .ZN(new_n521));
  AND4_X1   g320(.A1(new_n414), .A2(new_n415), .A3(new_n417), .A4(new_n418), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n405), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(new_n423), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT35), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n520), .A2(new_n524), .A3(new_n525), .A4(new_n476), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n518), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n253), .B1(new_n512), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G99gat), .B(G106gat), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(G85gat), .A2(G92gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G99gat), .A2(G106gat), .ZN(new_n534));
  INV_X1    g333(.A(G85gat), .ZN(new_n535));
  INV_X1    g334(.A(G92gat), .ZN(new_n536));
  AOI22_X1  g335(.A1(KEYINPUT8), .A2(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n530), .B1(new_n533), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n532), .B1(G85gat), .B2(G92gat), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n531), .B1(KEYINPUT98), .B2(KEYINPUT7), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n529), .B(new_n537), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT99), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n539), .A2(KEYINPUT99), .A3(new_n542), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n232), .A2(new_n548), .ZN(new_n549));
  AND2_X1   g348(.A1(G232gat), .A2(G233gat), .ZN(new_n550));
  AOI22_X1  g349(.A1(new_n216), .A2(new_n547), .B1(KEYINPUT41), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  XOR2_X1   g351(.A(G190gat), .B(G218gat), .Z(new_n553));
  AND2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n552), .A2(new_n553), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n550), .A2(KEYINPUT41), .ZN(new_n557));
  XNOR2_X1  g356(.A(G134gat), .B(G162gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n559), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n561), .B1(new_n554), .B2(new_n555), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G71gat), .A2(G78gat), .ZN(new_n565));
  INV_X1    g364(.A(G71gat), .ZN(new_n566));
  INV_X1    g365(.A(G78gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G57gat), .B(G64gat), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT9), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n565), .B(new_n568), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT96), .ZN(new_n572));
  AND2_X1   g371(.A1(KEYINPUT95), .A2(G64gat), .ZN(new_n573));
  NOR2_X1   g372(.A1(KEYINPUT95), .A2(G64gat), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n572), .B(G57gat), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n565), .B1(new_n568), .B2(new_n570), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(G64gat), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT96), .B1(new_n578), .B2(G57gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(KEYINPUT95), .B(G64gat), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n579), .B1(new_n580), .B2(G57gat), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n571), .B1(new_n577), .B2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(KEYINPUT97), .B(KEYINPUT21), .Z(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(G127gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n568), .A2(new_n565), .ZN(new_n589));
  INV_X1    g388(.A(G57gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(G64gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n578), .A2(G57gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n589), .B1(KEYINPUT9), .B2(new_n593), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n575), .A2(new_n576), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n573), .A2(new_n574), .ZN(new_n596));
  OAI211_X1 g395(.A(KEYINPUT96), .B(new_n591), .C1(new_n596), .C2(new_n590), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n594), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n229), .B1(KEYINPUT21), .B2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n588), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(new_n359), .ZN(new_n602));
  XOR2_X1   g401(.A(G183gat), .B(G211gat), .Z(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n600), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT100), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n542), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n598), .A2(new_n543), .A3(new_n611), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n542), .B(new_n539), .C1(new_n582), .C2(new_n610), .ZN(new_n613));
  AND2_X1   g412(.A1(G230gat), .A2(G233gat), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT102), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT10), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n582), .A2(new_n617), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n547), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n612), .A2(new_n613), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(new_n617), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT101), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n620), .A2(KEYINPUT101), .A3(new_n617), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n619), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n614), .B(KEYINPUT103), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n616), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G120gat), .B(G148gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(G176gat), .B(G204gat), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n628), .B(new_n629), .Z(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n616), .B(new_n630), .C1(new_n625), .C2(new_n614), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n564), .A2(new_n609), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n528), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n636), .A2(new_n479), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(new_n221), .ZN(G1324gat));
  OR3_X1    g437(.A1(new_n636), .A2(KEYINPUT104), .A3(new_n476), .ZN(new_n639));
  OAI21_X1  g438(.A(KEYINPUT104), .B1(new_n636), .B2(new_n476), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n639), .A2(G8gat), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n636), .ZN(new_n642));
  INV_X1    g441(.A(new_n476), .ZN(new_n643));
  XOR2_X1   g442(.A(KEYINPUT16), .B(G8gat), .Z(new_n644));
  NAND4_X1  g443(.A1(new_n642), .A2(KEYINPUT42), .A3(new_n643), .A4(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n644), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n646), .B1(new_n639), .B2(new_n640), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n641), .B(new_n645), .C1(new_n647), .C2(KEYINPUT42), .ZN(G1325gat));
  AOI21_X1  g447(.A(G15gat), .B1(new_n642), .B2(new_n514), .ZN(new_n649));
  INV_X1    g448(.A(new_n511), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(G15gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT105), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n649), .B1(new_n642), .B2(new_n652), .ZN(G1326gat));
  NAND2_X1  g452(.A1(new_n473), .A2(new_n469), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n636), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT43), .B(G22gat), .Z(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(G1327gat));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n511), .A2(new_n481), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n659), .B1(new_n426), .B2(new_n474), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT108), .ZN(new_n661));
  OAI211_X1 g460(.A(new_n476), .B(new_n514), .C1(new_n515), .C2(new_n516), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n525), .B1(new_n421), .B2(new_n424), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n525), .B1(new_n520), .B2(new_n513), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n661), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n518), .A2(new_n526), .A3(KEYINPUT108), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n660), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n658), .B1(new_n668), .B2(new_n563), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n512), .A2(new_n527), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n670), .A2(KEYINPUT44), .A3(new_n564), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n634), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n609), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n253), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(G29gat), .B1(new_n676), .B2(new_n479), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n563), .A2(new_n674), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n678), .B(KEYINPUT106), .Z(new_n679));
  NAND2_X1  g478(.A1(new_n528), .A2(new_n679), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n680), .A2(G29gat), .A3(new_n479), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n677), .A2(new_n683), .ZN(G1328gat));
  OAI21_X1  g483(.A(G36gat), .B1(new_n676), .B2(new_n476), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n680), .A2(G36gat), .A3(new_n476), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT46), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT109), .ZN(G1329gat));
  OR3_X1    g488(.A1(new_n680), .A2(G43gat), .A3(new_n519), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n672), .A2(new_n650), .A3(new_n675), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT110), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(G43gat), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n691), .A2(new_n692), .ZN(new_n695));
  OAI211_X1 g494(.A(KEYINPUT47), .B(new_n690), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n691), .A2(G43gat), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n697), .A2(new_n690), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n696), .B1(KEYINPUT47), .B2(new_n698), .ZN(G1330gat));
  INV_X1    g498(.A(new_n654), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(G50gat), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n680), .A2(new_n654), .ZN(new_n702));
  OAI22_X1  g501(.A1(new_n676), .A2(new_n701), .B1(G50gat), .B2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT48), .ZN(G1331gat));
  AND3_X1   g503(.A1(new_n518), .A2(new_n526), .A3(KEYINPUT108), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT108), .B1(new_n518), .B2(new_n526), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n512), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n564), .A2(new_n609), .A3(new_n673), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n707), .A2(new_n253), .A3(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(new_n479), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(new_n590), .ZN(G1332gat));
  XNOR2_X1  g510(.A(new_n709), .B(KEYINPUT111), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n643), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n713), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n714));
  XOR2_X1   g513(.A(KEYINPUT49), .B(G64gat), .Z(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n713), .B2(new_n715), .ZN(G1333gat));
  NOR3_X1   g515(.A1(new_n709), .A2(G71gat), .A3(new_n519), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n712), .A2(new_n650), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n717), .B1(new_n718), .B2(G71gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g519(.A1(new_n712), .A2(new_n700), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g521(.A1(new_n252), .A2(new_n608), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n634), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT112), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n672), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(G85gat), .B1(new_n726), .B2(new_n479), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n707), .A2(new_n564), .A3(new_n723), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT51), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n707), .A2(KEYINPUT51), .A3(new_n564), .A4(new_n723), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OR2_X1    g531(.A1(new_n732), .A2(new_n673), .ZN(new_n733));
  INV_X1    g532(.A(new_n479), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n535), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n727), .B1(new_n733), .B2(new_n735), .ZN(G1336gat));
  NAND4_X1  g535(.A1(new_n669), .A2(new_n643), .A3(new_n671), .A4(new_n725), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G92gat), .ZN(new_n738));
  XOR2_X1   g537(.A(KEYINPUT116), .B(KEYINPUT52), .Z(new_n739));
  NAND2_X1  g538(.A1(new_n643), .A2(new_n536), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n738), .B(new_n739), .C1(new_n733), .C2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n738), .A2(KEYINPUT113), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n730), .A2(KEYINPUT114), .A3(new_n731), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT114), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n744), .A3(new_n729), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n740), .A2(new_n673), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n743), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT113), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n737), .A2(new_n748), .A3(G92gat), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n742), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n750), .A2(KEYINPUT115), .A3(KEYINPUT52), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT115), .B1(new_n750), .B2(KEYINPUT52), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n741), .B1(new_n751), .B2(new_n752), .ZN(G1337gat));
  OAI21_X1  g552(.A(G99gat), .B1(new_n726), .B2(new_n511), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n514), .A2(new_n500), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n754), .B1(new_n733), .B2(new_n755), .ZN(G1338gat));
  OAI21_X1  g555(.A(G106gat), .B1(new_n726), .B2(new_n654), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT53), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n654), .A2(G106gat), .A3(new_n673), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n757), .B(new_n758), .C1(new_n732), .C2(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n743), .A2(new_n745), .A3(new_n759), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n763), .B2(new_n758), .ZN(G1339gat));
  NAND2_X1  g563(.A1(new_n547), .A2(new_n618), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT101), .B1(new_n620), .B2(new_n617), .ZN(new_n766));
  AOI211_X1 g565(.A(new_n622), .B(KEYINPUT10), .C1(new_n612), .C2(new_n613), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n626), .B(new_n765), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  OAI211_X1 g567(.A(KEYINPUT54), .B(new_n768), .C1(new_n625), .C2(new_n614), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT54), .ZN(new_n771));
  INV_X1    g570(.A(new_n626), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n769), .A2(KEYINPUT55), .A3(new_n631), .A4(new_n773), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n774), .A2(new_n633), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n769), .A2(new_n631), .A3(new_n773), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT117), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n777), .B1(new_n776), .B2(new_n778), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n775), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT118), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI211_X1 g582(.A(KEYINPUT118), .B(new_n775), .C1(new_n779), .C2(new_n780), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(new_n252), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n240), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n231), .B(new_n786), .C1(new_n229), .C2(new_n216), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n235), .B1(new_n231), .B2(new_n234), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n247), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n251), .A2(new_n790), .A3(new_n634), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n785), .A2(KEYINPUT119), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT119), .B1(new_n785), .B2(new_n791), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n792), .A2(new_n793), .A3(new_n564), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n783), .A2(new_n784), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n251), .A2(new_n790), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n795), .A2(new_n563), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n609), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n635), .A2(new_n253), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n479), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n800), .A2(new_n476), .A3(new_n520), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(G113gat), .B1(new_n802), .B2(new_n252), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n700), .B1(new_n798), .B2(new_n799), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n643), .A2(new_n479), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n804), .A2(new_n514), .A3(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT120), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n806), .B(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n253), .A2(new_n337), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n803), .B1(new_n809), .B2(new_n810), .ZN(G1340gat));
  AOI21_X1  g610(.A(G120gat), .B1(new_n802), .B2(new_n634), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n673), .A2(new_n335), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n812), .B1(new_n809), .B2(new_n813), .ZN(G1341gat));
  OAI21_X1  g613(.A(G127gat), .B1(new_n808), .B2(new_n609), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n802), .A2(new_n587), .A3(new_n608), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(G1342gat));
  NOR3_X1   g616(.A1(new_n563), .A2(G134gat), .A3(new_n643), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n800), .A2(new_n520), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n819), .B1(KEYINPUT121), .B2(KEYINPUT56), .ZN(new_n820));
  NAND2_X1  g619(.A1(KEYINPUT121), .A2(KEYINPUT56), .ZN(new_n821));
  XOR2_X1   g620(.A(new_n820), .B(new_n821), .Z(new_n822));
  OAI21_X1  g621(.A(G134gat), .B1(new_n808), .B2(new_n563), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(G1343gat));
  AND2_X1   g623(.A1(new_n511), .A2(new_n805), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n785), .A2(new_n791), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n564), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n785), .A2(KEYINPUT119), .A3(new_n791), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n797), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n799), .B1(new_n830), .B2(new_n608), .ZN(new_n831));
  AOI21_X1  g630(.A(KEYINPUT57), .B1(new_n831), .B2(new_n700), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n700), .A2(KEYINPUT57), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n776), .A2(new_n778), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n252), .A2(new_n775), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n564), .B1(new_n835), .B2(new_n791), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n609), .B1(new_n797), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n833), .B1(new_n837), .B2(new_n799), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n825), .B1(new_n832), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(G141gat), .B1(new_n839), .B2(new_n253), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n700), .A2(new_n511), .ZN(new_n841));
  XOR2_X1   g640(.A(new_n841), .B(KEYINPUT122), .Z(new_n842));
  NAND3_X1  g641(.A1(new_n800), .A2(new_n476), .A3(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n844), .A2(new_n348), .A3(new_n252), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT58), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT58), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n840), .A2(new_n845), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(G1344gat));
  OR3_X1    g649(.A1(new_n839), .A2(KEYINPUT59), .A3(new_n673), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT59), .B1(new_n843), .B2(new_n673), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n349), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n833), .B1(new_n798), .B2(new_n799), .ZN(new_n854));
  OR3_X1    g653(.A1(new_n563), .A2(new_n781), .A3(new_n796), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n609), .B1(new_n856), .B2(new_n836), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n799), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT57), .B1(new_n858), .B2(new_n700), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n854), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n825), .A2(new_n634), .ZN(new_n861));
  OAI211_X1 g660(.A(KEYINPUT59), .B(G148gat), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n851), .A2(new_n853), .A3(new_n862), .ZN(G1345gat));
  OAI21_X1  g662(.A(G155gat), .B1(new_n839), .B2(new_n609), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n844), .A2(new_n359), .A3(new_n608), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(G1346gat));
  OAI21_X1  g665(.A(G162gat), .B1(new_n839), .B2(new_n563), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n563), .A2(G162gat), .A3(new_n643), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n800), .A2(new_n842), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(G1347gat));
  NOR2_X1   g669(.A1(new_n734), .A2(new_n476), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(new_n519), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n804), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(G169gat), .B1(new_n874), .B2(new_n253), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n734), .B1(new_n798), .B2(new_n799), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(new_n643), .A3(new_n520), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n252), .A2(new_n278), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(G1348gat));
  OAI21_X1  g678(.A(G176gat), .B1(new_n874), .B2(new_n673), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n634), .A2(new_n268), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n880), .B1(new_n877), .B2(new_n881), .ZN(G1349gat));
  OAI21_X1  g681(.A(G183gat), .B1(new_n874), .B2(new_n609), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n608), .A2(new_n287), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n883), .B1(new_n877), .B2(new_n884), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g685(.A1(new_n804), .A2(new_n564), .A3(new_n873), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT61), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n887), .A2(new_n888), .A3(G190gat), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n887), .B2(G190gat), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n564), .A2(new_n286), .ZN(new_n891));
  OAI22_X1  g690(.A1(new_n889), .A2(new_n890), .B1(new_n877), .B2(new_n891), .ZN(G1351gat));
  NOR2_X1   g691(.A1(new_n841), .A2(new_n476), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(G197gat), .B1(new_n895), .B2(new_n252), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n650), .A2(new_n872), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n897), .B1(new_n854), .B2(new_n859), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n252), .A2(G197gat), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n896), .B1(new_n899), .B2(new_n900), .ZN(G1352gat));
  OAI21_X1  g700(.A(G204gat), .B1(new_n898), .B2(new_n673), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n673), .A2(G204gat), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n876), .A2(new_n903), .A3(new_n893), .A4(new_n904), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n831), .A2(new_n479), .A3(new_n893), .A4(new_n904), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(KEYINPUT123), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n908));
  AND3_X1   g707(.A1(new_n905), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n908), .B1(new_n905), .B2(new_n907), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n902), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(KEYINPUT124), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT124), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n913), .B(new_n902), .C1(new_n909), .C2(new_n910), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(G1353gat));
  AOI21_X1  g714(.A(new_n304), .B1(new_n899), .B2(new_n608), .ZN(new_n916));
  NAND2_X1  g715(.A1(KEYINPUT125), .A2(KEYINPUT63), .ZN(new_n917));
  OR2_X1    g716(.A1(KEYINPUT125), .A2(KEYINPUT63), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n895), .A2(new_n304), .A3(new_n608), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n919), .B(new_n920), .C1(new_n916), .C2(new_n917), .ZN(G1354gat));
  INV_X1    g720(.A(KEYINPUT126), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n898), .A2(new_n922), .ZN(new_n923));
  OAI211_X1 g722(.A(KEYINPUT126), .B(new_n897), .C1(new_n854), .C2(new_n859), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n563), .A2(new_n303), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(G218gat), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n927), .B1(new_n894), .B2(new_n563), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT127), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n926), .A2(new_n928), .A3(KEYINPUT127), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1355gat));
endmodule


