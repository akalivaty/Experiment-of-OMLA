//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 0 0 0 0 0 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1291,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358;
  OR3_X1    g0000(.A1(KEYINPUT64), .A2(G58), .A3(G68), .ZN(new_n201));
  OAI21_X1  g0001(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n202));
  AOI211_X1 g0002(.A(G50), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G87), .ZN(new_n215));
  INV_X1    g0015(.A(G250), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n218));
  INV_X1    g0018(.A(G58), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n208), .B1(new_n217), .B2(new_n223), .ZN(new_n224));
  OR2_X1    g0024(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n201), .A2(new_n202), .ZN(new_n226));
  INV_X1    g0026(.A(G50), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n206), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n211), .A2(new_n225), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n220), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  INV_X1    g0041(.A(G107), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G97), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n221), .A2(G107), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  INV_X1    g0052(.A(G45), .ZN(new_n253));
  AOI21_X1  g0053(.A(G1), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G1), .A3(G13), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(new_n256), .A3(G274), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n256), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(new_n254), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n260), .A2(G226), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT3), .B(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n262), .A2(G222), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G77), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n262), .A2(G1698), .ZN(new_n266));
  INV_X1    g0066(.A(G223), .ZN(new_n267));
  OAI221_X1 g0067(.A(new_n264), .B1(new_n265), .B2(new_n262), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  AOI211_X1 g0068(.A(new_n258), .B(new_n261), .C1(new_n268), .C2(new_n259), .ZN(new_n269));
  INV_X1    g0069(.A(G200), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n271), .B1(G190), .B2(new_n269), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n227), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n229), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n273), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT67), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n279), .A2(new_n280), .B1(new_n205), .B2(G20), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n281), .B1(new_n280), .B2(new_n279), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n275), .B1(new_n282), .B2(new_n227), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT8), .B(G58), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT65), .ZN(new_n285));
  OR3_X1    g0085(.A1(new_n219), .A2(KEYINPUT65), .A3(KEYINPUT8), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G33), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(G20), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G150), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  OAI22_X1  g0093(.A1(new_n287), .A2(new_n290), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n206), .B1(new_n226), .B2(new_n227), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n277), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n283), .B1(KEYINPUT66), .B2(new_n296), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n296), .A2(KEYINPUT66), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(KEYINPUT9), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT9), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n301), .B1(new_n297), .B2(new_n298), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n272), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT10), .ZN(new_n304));
  INV_X1    g0104(.A(G179), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n269), .A2(new_n305), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n299), .B(new_n306), .C1(G169), .C2(new_n269), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n219), .A2(new_n213), .ZN(new_n309));
  OAI21_X1  g0109(.A(G20), .B1(new_n226), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n292), .A2(G159), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n288), .A2(KEYINPUT3), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  AND2_X1   g0115(.A1(KEYINPUT72), .A2(KEYINPUT3), .ZN(new_n316));
  NOR2_X1   g0116(.A1(KEYINPUT72), .A2(KEYINPUT3), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n315), .B1(new_n318), .B2(G33), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n206), .A2(KEYINPUT7), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT73), .ZN(new_n322));
  NOR3_X1   g0122(.A1(new_n316), .A2(new_n317), .A3(new_n288), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n322), .B1(new_n323), .B2(new_n315), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT72), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT3), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(KEYINPUT72), .A2(KEYINPUT3), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(G33), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n329), .A2(KEYINPUT73), .A3(new_n314), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n324), .A2(new_n206), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT7), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n321), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI211_X1 g0133(.A(KEYINPUT16), .B(new_n313), .C1(new_n333), .C2(new_n213), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT16), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n288), .B1(new_n316), .B2(new_n317), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n326), .A2(G33), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n320), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n314), .A2(new_n337), .ZN(new_n339));
  AOI21_X1  g0139(.A(KEYINPUT7), .B1(new_n339), .B2(new_n206), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n341), .A2(new_n213), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n335), .B1(new_n342), .B2(new_n312), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n334), .A2(new_n343), .A3(new_n277), .ZN(new_n344));
  INV_X1    g0144(.A(new_n287), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n282), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n287), .A2(new_n273), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT74), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT74), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n344), .A2(new_n351), .A3(new_n348), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n258), .B1(G232), .B2(new_n260), .ZN(new_n353));
  AND2_X1   g0153(.A1(G226), .A2(G1698), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n319), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT75), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n319), .A2(KEYINPUT75), .A3(new_n354), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n267), .A2(G1698), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n319), .A2(new_n360), .B1(G33), .B2(G87), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g0162(.A(G179), .B(new_n353), .C1(new_n362), .C2(new_n256), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n256), .B1(new_n359), .B2(new_n361), .ZN(new_n364));
  INV_X1    g0164(.A(new_n353), .ZN(new_n365));
  OAI21_X1  g0165(.A(G169), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n350), .A2(new_n352), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT18), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT18), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n350), .A2(new_n370), .A3(new_n352), .A4(new_n367), .ZN(new_n371));
  INV_X1    g0171(.A(G190), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n372), .A2(KEYINPUT76), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n372), .A2(KEYINPUT76), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n353), .B(new_n376), .C1(new_n362), .C2(new_n256), .ZN(new_n377));
  OAI21_X1  g0177(.A(G200), .B1(new_n364), .B2(new_n365), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n344), .A2(new_n377), .A3(new_n348), .A4(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT77), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n380), .A2(KEYINPUT17), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(KEYINPUT17), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n379), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n349), .ZN(new_n384));
  AND2_X1   g0184(.A1(new_n377), .A2(new_n378), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n384), .A2(new_n385), .A3(new_n380), .A4(KEYINPUT17), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n369), .A2(new_n371), .A3(new_n383), .A4(new_n386), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n292), .A2(G50), .B1(G20), .B2(new_n213), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n290), .B2(new_n265), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n277), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT11), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n389), .A2(KEYINPUT11), .A3(new_n277), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n394), .A2(KEYINPUT71), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(KEYINPUT71), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT12), .B1(new_n273), .B2(G68), .ZN(new_n397));
  OR3_X1    g0197(.A1(new_n273), .A2(KEYINPUT12), .A3(G68), .ZN(new_n398));
  INV_X1    g0198(.A(new_n279), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n213), .B1(new_n205), .B2(G20), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n397), .A2(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n395), .A2(new_n396), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n262), .A2(G232), .A3(G1698), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n262), .A2(G226), .A3(new_n263), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G97), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT70), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT70), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n403), .A2(new_n404), .A3(new_n408), .A4(new_n405), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n407), .A2(new_n259), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n258), .B1(G238), .B2(new_n260), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT13), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT13), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n410), .A2(new_n414), .A3(new_n411), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n413), .A2(G179), .A3(new_n415), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n410), .A2(new_n414), .A3(new_n411), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n414), .B1(new_n410), .B2(new_n411), .ZN(new_n418));
  OAI21_X1  g0218(.A(G169), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n416), .B1(new_n419), .B2(KEYINPUT14), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT14), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n413), .A2(new_n415), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n421), .B1(new_n422), .B2(G169), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n402), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n402), .ZN(new_n425));
  OAI21_X1  g0225(.A(G200), .B1(new_n417), .B2(new_n418), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n413), .A2(G190), .A3(new_n415), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  OAI22_X1  g0229(.A1(new_n266), .A2(new_n214), .B1(new_n242), .B2(new_n262), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n339), .A2(new_n220), .A3(G1698), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n259), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n258), .B1(G244), .B2(new_n260), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(G200), .ZN(new_n435));
  INV_X1    g0235(.A(new_n434), .ZN(new_n436));
  AOI22_X1  g0236(.A1(KEYINPUT68), .A2(new_n435), .B1(new_n436), .B2(G190), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT68), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n434), .A2(new_n438), .A3(new_n372), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n284), .B1(KEYINPUT69), .B2(new_n293), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(KEYINPUT69), .B2(new_n293), .ZN(new_n441));
  XNOR2_X1  g0241(.A(KEYINPUT15), .B(G87), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n443), .A2(new_n289), .B1(G20), .B2(G77), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n278), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(G77), .B1(new_n206), .B2(G1), .ZN(new_n446));
  OAI22_X1  g0246(.A1(new_n279), .A2(new_n446), .B1(G77), .B2(new_n273), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NOR3_X1   g0249(.A1(new_n437), .A2(new_n439), .A3(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n449), .B1(new_n436), .B2(G169), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n434), .A2(G179), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g0255(.A1(new_n308), .A2(new_n387), .A3(new_n429), .A4(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n273), .A2(G97), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n205), .A2(G33), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n273), .A2(new_n459), .A3(new_n229), .A4(new_n276), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n458), .B1(new_n461), .B2(G97), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n292), .A2(G77), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT6), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n464), .A2(new_n221), .A3(G107), .ZN(new_n465));
  XNOR2_X1  g0265(.A(G97), .B(G107), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n465), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n463), .B1(new_n467), .B2(new_n206), .ZN(new_n468));
  OAI21_X1  g0268(.A(G107), .B1(new_n338), .B2(new_n340), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n468), .B1(new_n469), .B2(KEYINPUT78), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT78), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n471), .B(G107), .C1(new_n338), .C2(new_n340), .ZN(new_n472));
  AOI211_X1 g0272(.A(KEYINPUT79), .B(new_n278), .C1(new_n470), .C2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT79), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n469), .A2(KEYINPUT78), .ZN(new_n475));
  INV_X1    g0275(.A(new_n468), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n475), .A2(new_n472), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n474), .B1(new_n477), .B2(new_n277), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n462), .B1(new_n473), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n253), .A2(G1), .ZN(new_n480));
  AND2_X1   g0280(.A1(KEYINPUT5), .A2(G41), .ZN(new_n481));
  NOR2_X1   g0281(.A1(KEYINPUT5), .A2(G41), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G274), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n483), .A2(new_n259), .A3(new_n484), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n483), .A2(new_n256), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n485), .B1(G257), .B2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G244), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(G1698), .ZN(new_n490));
  AOI21_X1  g0290(.A(KEYINPUT80), .B1(new_n319), .B2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n329), .A2(KEYINPUT80), .A3(new_n314), .A4(new_n490), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(KEYINPUT81), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n329), .A2(new_n314), .A3(new_n490), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT80), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT81), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n498), .A2(new_n499), .A3(new_n493), .A4(new_n492), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n262), .A2(KEYINPUT4), .A3(new_n490), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n262), .A2(G250), .A3(G1698), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G283), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n495), .A2(new_n500), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n488), .B1(new_n505), .B2(new_n259), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n506), .A2(new_n270), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n479), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT83), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n500), .A2(new_n504), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n492), .A2(new_n493), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n499), .B1(new_n511), .B2(new_n498), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n259), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n487), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT82), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT82), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n506), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n515), .A2(G190), .A3(new_n517), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n508), .A2(new_n509), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n509), .B1(new_n508), .B2(new_n518), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(G169), .B1(new_n515), .B2(new_n517), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n506), .A2(new_n305), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n479), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(G238), .A2(G1698), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n527), .B1(new_n489), .B2(G1698), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n528), .A2(new_n329), .A3(new_n314), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G116), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT86), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n529), .A2(KEYINPUT86), .A3(new_n530), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n533), .A2(new_n259), .A3(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT84), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n205), .A2(G45), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n256), .A2(new_n536), .A3(G250), .A4(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n256), .A2(G274), .A3(new_n480), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n480), .A2(new_n216), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n536), .B1(new_n541), .B2(new_n256), .ZN(new_n542));
  OAI21_X1  g0342(.A(KEYINPUT85), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n537), .A2(G250), .ZN(new_n544));
  OAI21_X1  g0344(.A(KEYINPUT84), .B1(new_n259), .B2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT85), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n545), .A2(new_n546), .A3(new_n539), .A4(new_n538), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n535), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(G169), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT19), .B1(new_n289), .B2(G97), .ZN(new_n551));
  XNOR2_X1  g0351(.A(KEYINPUT88), .B(G87), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n552), .A2(new_n221), .A3(new_n242), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT19), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(new_n405), .B2(new_n206), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n551), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n329), .A2(new_n206), .A3(G68), .A4(new_n314), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n278), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n443), .A2(new_n273), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n460), .A2(new_n442), .ZN(new_n561));
  XNOR2_X1  g0361(.A(new_n561), .B(KEYINPUT89), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n549), .A2(new_n550), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT87), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n549), .B2(G179), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n549), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n567), .A2(KEYINPUT87), .A3(new_n305), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n461), .A2(G87), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n560), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n270), .B1(new_n535), .B2(new_n548), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n567), .B2(G190), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n566), .A2(new_n568), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n526), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n329), .A2(new_n314), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n222), .A2(G1698), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(G250), .B2(G1698), .ZN(new_n578));
  INV_X1    g0378(.A(G294), .ZN(new_n579));
  OAI22_X1  g0379(.A1(new_n576), .A2(new_n578), .B1(new_n288), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n259), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT92), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT92), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n580), .A2(new_n583), .A3(new_n259), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n483), .A2(G264), .A3(new_n256), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT93), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT93), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n483), .A2(new_n587), .A3(G264), .A4(new_n256), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n485), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n582), .A2(new_n584), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G169), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n485), .B1(new_n580), .B2(new_n259), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT94), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n586), .A2(new_n593), .A3(new_n588), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n593), .B1(new_n586), .B2(new_n588), .ZN(new_n595));
  OAI211_X1 g0395(.A(G179), .B(new_n592), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT23), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(G20), .B2(new_n242), .ZN(new_n599));
  XNOR2_X1  g0399(.A(new_n599), .B(KEYINPUT91), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT22), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n206), .A2(G87), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n601), .B1(new_n339), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n598), .A2(new_n242), .A3(G20), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n600), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n329), .A2(KEYINPUT22), .A3(G87), .A4(new_n314), .ZN(new_n606));
  AOI21_X1  g0406(.A(G20), .B1(new_n606), .B2(new_n530), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT24), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n605), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n600), .A2(new_n603), .A3(new_n604), .ZN(new_n611));
  OAI21_X1  g0411(.A(KEYINPUT24), .B1(new_n611), .B2(new_n607), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n278), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n274), .A2(KEYINPUT25), .A3(new_n242), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT25), .B1(new_n274), .B2(new_n242), .ZN(new_n616));
  OAI22_X1  g0416(.A1(new_n615), .A2(new_n616), .B1(new_n242), .B2(new_n460), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n597), .B1(new_n613), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n610), .A2(new_n612), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n617), .B1(new_n619), .B2(new_n277), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n592), .B1(new_n594), .B2(new_n595), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n621), .A2(new_n270), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n590), .A2(G190), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n485), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n486), .A2(G270), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n339), .A2(G303), .ZN(new_n628));
  NAND2_X1  g0428(.A1(G264), .A2(G1698), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n628), .B1(new_n576), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT90), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n319), .A2(new_n631), .A3(G257), .A4(new_n263), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n263), .A2(G257), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT90), .B1(new_n576), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n630), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n626), .B(new_n627), .C1(new_n635), .C2(new_n256), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(G200), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n503), .B(new_n206), .C1(G33), .C2(new_n221), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n638), .B(new_n277), .C1(new_n206), .C2(G116), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT20), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n273), .A2(G116), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n461), .B2(G116), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n637), .B(new_n644), .C1(new_n375), .C2(new_n636), .ZN(new_n645));
  OR3_X1    g0445(.A1(new_n636), .A2(new_n644), .A3(new_n305), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT21), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n550), .B1(new_n641), .B2(new_n643), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n647), .B1(new_n636), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n636), .A2(new_n648), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(KEYINPUT21), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n645), .B(new_n646), .C1(new_n649), .C2(new_n651), .ZN(new_n652));
  NOR4_X1   g0452(.A1(new_n457), .A2(new_n575), .A3(new_n625), .A4(new_n652), .ZN(G372));
  INV_X1    g0453(.A(new_n304), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n349), .A2(new_n367), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT18), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n386), .A2(new_n383), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n428), .A2(new_n453), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n424), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n656), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n307), .B1(new_n654), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n567), .A2(new_n305), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n563), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n570), .A2(KEYINPUT95), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT95), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n560), .A2(new_n668), .A3(new_n569), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n670), .A2(new_n573), .B1(new_n664), .B2(new_n563), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n525), .A2(new_n666), .A3(new_n671), .ZN(new_n672));
  AOI211_X1 g0472(.A(KEYINPUT82), .B(new_n488), .C1(new_n505), .C2(new_n259), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n516), .B1(new_n513), .B2(new_n487), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n550), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n479), .A2(new_n523), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n574), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n665), .B(new_n672), .C1(new_n677), .C2(new_n666), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n675), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n618), .B(new_n646), .C1(new_n649), .C2(new_n651), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n679), .A2(new_n680), .A3(new_n624), .A4(new_n671), .ZN(new_n681));
  OAI21_X1  g0481(.A(KEYINPUT96), .B1(new_n521), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n646), .B1(new_n651), .B2(new_n649), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n620), .B1(new_n591), .B2(new_n596), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n671), .B(new_n624), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(new_n525), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT96), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n673), .A2(new_n674), .A3(new_n372), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n514), .A2(G200), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n477), .A2(new_n277), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT79), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n477), .A2(new_n474), .A3(new_n277), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n689), .A2(new_n693), .A3(new_n462), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT83), .B1(new_n688), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n508), .A2(new_n518), .A3(new_n509), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n686), .A2(new_n687), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n678), .B1(new_n682), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n663), .B1(new_n457), .B2(new_n699), .ZN(G369));
  INV_X1    g0500(.A(new_n652), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(G213), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(G343), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n644), .A2(new_n708), .ZN(new_n709));
  MUX2_X1   g0509(.A(new_n701), .B(new_n683), .S(new_n709), .Z(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G330), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n620), .A2(new_n708), .ZN(new_n713));
  OAI22_X1  g0513(.A1(new_n625), .A2(new_n713), .B1(new_n618), .B2(new_n708), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n683), .A2(new_n708), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(new_n625), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n618), .A2(new_n707), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n715), .A2(new_n719), .ZN(G399));
  INV_X1    g0520(.A(KEYINPUT29), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT99), .B1(new_n699), .B2(new_n707), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT99), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(new_n699), .B2(new_n707), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n521), .A2(new_n681), .ZN(new_n725));
  INV_X1    g0525(.A(new_n671), .ZN(new_n726));
  OAI21_X1  g0526(.A(KEYINPUT26), .B1(new_n679), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n525), .A2(new_n666), .A3(new_n574), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(new_n665), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n708), .B1(new_n725), .B2(new_n729), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n730), .A2(KEYINPUT29), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n721), .A2(new_n722), .B1(new_n724), .B2(new_n731), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n652), .A2(new_n625), .A3(new_n707), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n697), .A2(new_n733), .A3(new_n679), .A4(new_n574), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n627), .B1(new_n635), .B2(new_n256), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n596), .A2(new_n735), .A3(new_n549), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n515), .A2(new_n517), .A3(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT30), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n515), .A2(new_n736), .A3(new_n517), .A4(KEYINPUT30), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT98), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n549), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n535), .A2(KEYINPUT98), .A3(new_n548), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n636), .A2(new_n305), .A3(new_n621), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n744), .A2(new_n745), .A3(new_n506), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n739), .A2(new_n740), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n707), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT31), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n748), .A2(KEYINPUT31), .A3(new_n707), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n734), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G330), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n732), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n205), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT97), .ZN(new_n757));
  INV_X1    g0557(.A(new_n209), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n757), .B1(new_n758), .B2(G41), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n209), .A2(KEYINPUT97), .A3(new_n252), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n553), .A2(G116), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n761), .A2(G1), .A3(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n228), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n763), .B1(new_n764), .B2(new_n761), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT28), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n756), .A2(new_n766), .ZN(G364));
  INV_X1    g0567(.A(new_n761), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n206), .A2(G13), .ZN(new_n769));
  XOR2_X1   g0569(.A(new_n769), .B(KEYINPUT100), .Z(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G45), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G1), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n710), .A2(G330), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n712), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT101), .Z(new_n776));
  INV_X1    g0576(.A(new_n773), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n229), .B1(G20), .B2(new_n550), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n372), .A2(G179), .A3(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n206), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n579), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n206), .A2(new_n305), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G200), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(G190), .ZN(new_n785));
  XNOR2_X1  g0585(.A(KEYINPUT33), .B(G317), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n783), .A2(new_n270), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(G190), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G311), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n787), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n375), .A2(new_n784), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n782), .B(new_n792), .C1(G326), .C2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n375), .A2(new_n788), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT102), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n375), .A2(new_n788), .A3(KEYINPUT102), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G322), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n270), .A2(G179), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n802), .A2(G20), .A3(G190), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n262), .B1(new_n804), .B2(G303), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n206), .A2(G190), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n806), .A2(new_n305), .A3(new_n270), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n806), .A2(new_n802), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  AOI22_X1  g0610(.A1(G329), .A2(new_n808), .B1(new_n810), .B2(G283), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n794), .A2(new_n801), .A3(new_n805), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n800), .A2(G58), .ZN(new_n813));
  INV_X1    g0613(.A(new_n793), .ZN(new_n814));
  INV_X1    g0614(.A(new_n785), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n814), .A2(new_n227), .B1(new_n815), .B2(new_n213), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n790), .A2(new_n265), .B1(new_n221), .B2(new_n781), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(G159), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n807), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT32), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n262), .B1(new_n803), .B2(new_n552), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n809), .A2(new_n242), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n813), .A2(new_n818), .A3(new_n821), .A4(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n779), .B1(new_n812), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(G13), .A2(G33), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(G20), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(new_n778), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n324), .A2(new_n330), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n831), .A2(new_n758), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n250), .A2(G45), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n832), .B(new_n833), .C1(G45), .C2(new_n764), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n758), .A2(new_n339), .ZN(new_n835));
  INV_X1    g0635(.A(G116), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n835), .A2(G355), .B1(new_n836), .B2(new_n758), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n777), .B(new_n826), .C1(new_n830), .C2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n829), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n710), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n776), .A2(new_n841), .ZN(G396));
  NOR2_X1   g0642(.A1(new_n778), .A2(new_n827), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n777), .B1(new_n265), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n262), .B1(new_n810), .B2(G87), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n845), .B1(new_n242), .B2(new_n803), .C1(new_n791), .C2(new_n807), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n793), .A2(G303), .B1(new_n785), .B2(G283), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n847), .B1(new_n221), .B2(new_n781), .C1(new_n836), .C2(new_n790), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n846), .B(new_n848), .C1(G294), .C2(new_n800), .ZN(new_n849));
  INV_X1    g0649(.A(new_n831), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n809), .A2(new_n213), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(G50), .B2(new_n804), .ZN(new_n852));
  INV_X1    g0652(.A(G132), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n852), .B1(new_n219), .B2(new_n781), .C1(new_n853), .C2(new_n807), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n793), .A2(G137), .B1(new_n789), .B2(G159), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n291), .B2(new_n815), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(new_n800), .B2(G143), .ZN(new_n857));
  XOR2_X1   g0657(.A(KEYINPUT103), .B(KEYINPUT34), .Z(new_n858));
  AOI211_X1 g0658(.A(new_n850), .B(new_n854), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  OR2_X1    g0659(.A1(new_n857), .A2(new_n858), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n849), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n448), .A2(new_n708), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n450), .A2(new_n862), .B1(new_n452), .B2(new_n451), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n453), .A2(new_n708), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n844), .B1(new_n779), .B2(new_n861), .C1(new_n865), .C2(new_n828), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n455), .A2(new_n707), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n699), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n865), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n699), .B2(new_n707), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT104), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT104), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n873), .B(new_n870), .C1(new_n699), .C2(new_n707), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n869), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(G330), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n746), .B1(new_n737), .B2(new_n738), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n750), .B(new_n708), .C1(new_n877), .C2(new_n740), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT31), .B1(new_n748), .B2(new_n707), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n876), .B1(new_n880), .B2(new_n734), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n777), .B1(new_n875), .B2(new_n881), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n754), .B(new_n869), .C1(new_n872), .C2(new_n874), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n866), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT105), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(KEYINPUT105), .B(new_n866), .C1(new_n882), .C2(new_n883), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(G384));
  NAND2_X1  g0688(.A1(new_n722), .A2(new_n721), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n724), .A2(new_n731), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n662), .B1(new_n891), .B2(new_n456), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n892), .B(KEYINPUT106), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n334), .A2(new_n277), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n313), .B1(new_n333), .B2(new_n213), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n335), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n894), .A2(new_n896), .B1(new_n346), .B2(new_n347), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n897), .A2(new_n705), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n387), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n379), .B1(new_n897), .B2(new_n705), .ZN(new_n900));
  INV_X1    g0700(.A(new_n367), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT37), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n705), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n350), .A2(new_n352), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT37), .B1(new_n384), .B2(new_n385), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n368), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n899), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT38), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n899), .A2(KEYINPUT38), .A3(new_n908), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n911), .A2(KEYINPUT39), .A3(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT39), .ZN(new_n914));
  AOI221_X4 g0714(.A(new_n910), .B1(new_n903), .B2(new_n907), .C1(new_n387), .C2(new_n898), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n905), .A2(new_n379), .A3(new_n655), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT37), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n907), .ZN(new_n918));
  INV_X1    g0718(.A(new_n905), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n656), .B2(new_n657), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT38), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n914), .B1(new_n915), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n419), .A2(KEYINPUT14), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n422), .A2(new_n421), .A3(G169), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n923), .A2(new_n924), .A3(new_n416), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(new_n402), .A3(new_n708), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n913), .A2(new_n922), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n864), .B1(new_n699), .B2(new_n868), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n911), .A2(new_n912), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n402), .A2(new_n707), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n424), .A2(new_n428), .A3(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n428), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n402), .B(new_n707), .C1(new_n925), .C2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n929), .A2(new_n930), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n656), .A2(new_n705), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n928), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n893), .B(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n935), .A2(new_n865), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n880), .B2(new_n734), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT38), .B1(new_n899), .B2(new_n908), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n941), .B1(new_n915), .B2(new_n942), .ZN(new_n943));
  XOR2_X1   g0743(.A(KEYINPUT107), .B(KEYINPUT40), .Z(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n940), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n753), .A2(new_n946), .A3(KEYINPUT40), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n368), .A2(new_n906), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n948), .A2(new_n905), .B1(new_n916), .B2(KEYINPUT37), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n655), .B(new_n370), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n905), .B1(new_n658), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n910), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n912), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n943), .A2(new_n945), .B1(new_n947), .B2(new_n953), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n456), .A2(new_n753), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n954), .A2(new_n955), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n956), .A2(new_n957), .A3(new_n876), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n939), .A2(new_n958), .B1(new_n205), .B2(new_n770), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(new_n939), .B2(new_n958), .ZN(new_n960));
  INV_X1    g0760(.A(new_n467), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n961), .A2(KEYINPUT35), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(KEYINPUT35), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n962), .A2(G116), .A3(new_n230), .A4(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT36), .Z(new_n965));
  OAI211_X1 g0765(.A(new_n228), .B(G77), .C1(new_n219), .C2(new_n213), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n227), .A2(G68), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n205), .B(G13), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  OR3_X1    g0768(.A1(new_n960), .A2(new_n965), .A3(new_n968), .ZN(G367));
  NAND2_X1  g0769(.A1(new_n479), .A2(new_n707), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n526), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n525), .A2(new_n707), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n717), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n679), .B1(new_n971), .B2(new_n618), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n974), .A2(KEYINPUT42), .B1(new_n975), .B2(new_n708), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT109), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n974), .A2(KEYINPUT42), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n976), .A2(new_n977), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n671), .B1(new_n670), .B2(new_n708), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n982), .A2(KEYINPUT108), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(KEYINPUT108), .ZN(new_n984));
  OR3_X1    g0784(.A1(new_n665), .A2(new_n670), .A3(new_n708), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT43), .Z(new_n987));
  NAND2_X1  g0787(.A1(new_n981), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n978), .A2(new_n989), .A3(new_n979), .A4(new_n980), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n990), .A2(KEYINPUT110), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n990), .A2(KEYINPUT110), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n988), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n971), .A2(new_n972), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n994), .A2(new_n715), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n772), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n973), .A2(KEYINPUT45), .A3(new_n719), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT45), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n719), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1000), .B1(new_n994), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n994), .A2(KEYINPUT44), .A3(new_n1001), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT44), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n973), .B2(new_n719), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n999), .A2(new_n1002), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n715), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n717), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n716), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1009), .B1(new_n714), .B2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n711), .B(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n755), .B1(new_n1008), .B2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n761), .B(KEYINPUT41), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n998), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n995), .B(new_n988), .C1(new_n991), .C2(new_n992), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n997), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n832), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n830), .B1(new_n209), .B2(new_n442), .C1(new_n1019), .C2(new_n240), .ZN(new_n1020));
  AND2_X1   g0820(.A1(new_n1020), .A2(new_n773), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n800), .A2(G150), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n809), .A2(new_n265), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n262), .B1(new_n803), .B2(new_n219), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n1023), .B(new_n1024), .C1(G137), .C2(new_n808), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n781), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G68), .A2(new_n1026), .B1(new_n789), .B2(G50), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n793), .A2(G143), .B1(new_n785), .B2(G159), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1022), .A2(new_n1025), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(G283), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n803), .A2(new_n836), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n790), .A2(new_n1030), .B1(KEYINPUT46), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(KEYINPUT46), .B2(new_n1031), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n810), .A2(G97), .ZN(new_n1034));
  INV_X1    g0834(.A(G317), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1034), .B1(new_n1035), .B2(new_n807), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(G294), .B2(new_n785), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n793), .A2(G311), .B1(new_n1026), .B2(G107), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1033), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(G303), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n850), .B1(new_n799), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1029), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT47), .Z(new_n1043));
  OAI221_X1 g0843(.A(new_n1021), .B1(new_n779), .B2(new_n1043), .C1(new_n986), .C2(new_n840), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1018), .A2(new_n1044), .ZN(G387));
  AOI21_X1  g0845(.A(new_n850), .B1(new_n800), .B2(G50), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n781), .A2(new_n442), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n790), .A2(new_n213), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(G159), .C2(new_n793), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n804), .A2(G77), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1050), .B(new_n1034), .C1(new_n291), .C2(new_n807), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n345), .B2(new_n785), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1046), .A2(new_n1049), .A3(new_n1052), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G326), .A2(new_n808), .B1(new_n810), .B2(G116), .ZN(new_n1054));
  INV_X1    g0854(.A(G322), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n814), .A2(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n815), .A2(new_n791), .B1(new_n790), .B2(new_n1040), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(new_n800), .C2(G317), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1058), .A2(KEYINPUT48), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(KEYINPUT48), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1026), .A2(G283), .B1(new_n804), .B2(G294), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT111), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT49), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n850), .B(new_n1054), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1053), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n778), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n237), .A2(new_n253), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n762), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n1069), .A2(new_n832), .B1(new_n1070), .B2(new_n835), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n284), .A2(G50), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT50), .Z(new_n1073));
  OAI21_X1  g0873(.A(new_n253), .B1(new_n213), .B2(new_n265), .ZN(new_n1074));
  NOR3_X1   g0874(.A1(new_n1073), .A2(new_n1070), .A3(new_n1074), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n1071), .A2(new_n1075), .B1(G107), .B2(new_n209), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n777), .B1(new_n1076), .B2(new_n830), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1068), .B(new_n1077), .C1(new_n714), .C2(new_n840), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n732), .A2(new_n754), .A3(new_n1013), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n768), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1013), .B1(new_n732), .B2(new_n754), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1078), .B1(new_n998), .B2(new_n1012), .C1(new_n1080), .C2(new_n1081), .ZN(G393));
  INV_X1    g0882(.A(KEYINPUT113), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1002), .A2(new_n999), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1083), .B(new_n1007), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(KEYINPUT113), .B1(new_n1006), .B2(new_n715), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT114), .ZN(new_n1089));
  AOI21_X1  g0889(.A(KEYINPUT112), .B1(new_n1006), .B2(new_n715), .ZN(new_n1090));
  AND3_X1   g0890(.A1(new_n1006), .A2(KEYINPUT112), .A3(new_n715), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1088), .B(new_n1089), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1091), .A2(new_n1090), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1094));
  OAI21_X1  g0894(.A(KEYINPUT114), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1092), .A2(new_n1095), .A3(new_n772), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1079), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1008), .A2(new_n754), .A3(new_n732), .A4(new_n1013), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1097), .A2(new_n768), .A3(new_n1098), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n830), .B1(new_n221), .B2(new_n209), .C1(new_n1019), .C2(new_n247), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n773), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n799), .A2(new_n819), .B1(new_n291), .B2(new_n814), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT51), .Z(new_n1103));
  OAI22_X1  g0903(.A1(new_n815), .A2(new_n227), .B1(new_n790), .B2(new_n284), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT115), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G143), .A2(new_n808), .B1(new_n810), .B2(G87), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n1106), .B1(new_n213), .B2(new_n803), .C1(new_n265), .C2(new_n781), .ZN(new_n1107));
  OR3_X1    g0907(.A1(new_n1105), .A2(new_n850), .A3(new_n1107), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n799), .A2(new_n791), .B1(new_n1035), .B2(new_n814), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n1109), .B(KEYINPUT52), .Z(new_n1110));
  OAI22_X1  g0910(.A1(new_n803), .A2(new_n1030), .B1(new_n807), .B2(new_n1055), .ZN(new_n1111));
  NOR3_X1   g0911(.A1(new_n1111), .A2(new_n262), .A3(new_n823), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(G294), .A2(new_n789), .B1(new_n785), .B2(G303), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1112), .B(new_n1113), .C1(new_n836), .C2(new_n781), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n1103), .A2(new_n1108), .B1(new_n1110), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1101), .B1(new_n1115), .B2(new_n778), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n973), .B2(new_n840), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1096), .A2(new_n1099), .A3(new_n1117), .ZN(G390));
  NAND4_X1  g0918(.A1(new_n753), .A2(G330), .A3(new_n865), .A4(new_n935), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n864), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n682), .A2(new_n698), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n678), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1120), .B1(new_n1123), .B2(new_n867), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n935), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n926), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT117), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n913), .A2(new_n922), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n927), .B1(new_n929), .B2(new_n935), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(KEYINPUT117), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1128), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n927), .B1(new_n952), .B2(new_n912), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n708), .B(new_n863), .C1(new_n725), .C2(new_n729), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n864), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(KEYINPUT116), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT116), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1134), .A2(new_n1137), .A3(new_n864), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1133), .B1(new_n1139), .B2(new_n1125), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1119), .B1(new_n1132), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1129), .B1(new_n1130), .B2(KEYINPUT117), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1127), .B(new_n927), .C1(new_n929), .C2(new_n935), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1140), .B(new_n1119), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n457), .A2(new_n754), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1147), .B(new_n663), .C1(new_n732), .C2(new_n457), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT118), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1119), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1125), .B1(new_n754), .B2(new_n870), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1124), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n935), .B1(new_n881), .B2(new_n865), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1119), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1153), .B1(new_n1154), .B2(KEYINPUT118), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n1152), .A2(new_n1155), .B1(new_n1139), .B2(new_n1156), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n1141), .A2(new_n1145), .B1(new_n1148), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1140), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n1154), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1157), .A2(new_n1148), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1160), .A2(new_n1161), .A3(new_n1144), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1158), .A2(new_n768), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n777), .B1(new_n287), .B2(new_n843), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT119), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(KEYINPUT54), .B(G143), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(G137), .A2(new_n785), .B1(new_n789), .B2(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n800), .A2(G132), .B1(new_n1165), .B2(new_n1168), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n1168), .A2(new_n1165), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n804), .A2(G150), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT53), .ZN(new_n1173));
  INV_X1    g0973(.A(G128), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n814), .A2(new_n1174), .B1(new_n781), .B2(new_n819), .ZN(new_n1175));
  INV_X1    g0975(.A(G125), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n262), .B1(new_n809), .B2(new_n227), .C1(new_n1176), .C2(new_n807), .ZN(new_n1177));
  NOR3_X1   g0977(.A1(new_n1173), .A2(new_n1175), .A3(new_n1177), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n793), .A2(G283), .B1(new_n789), .B2(G97), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n265), .B2(new_n781), .C1(new_n242), .C2(new_n815), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n803), .A2(new_n215), .B1(new_n807), .B2(new_n579), .ZN(new_n1181));
  NOR4_X1   g0981(.A1(new_n1180), .A2(new_n262), .A3(new_n851), .A4(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n800), .A2(G116), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n1171), .A2(new_n1178), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1164), .B1(new_n1184), .B2(new_n779), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n1129), .B2(new_n827), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1141), .A2(new_n1145), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1186), .B1(new_n1187), .B2(new_n772), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1163), .A2(new_n1188), .ZN(G378));
  NAND2_X1  g0989(.A1(new_n943), .A2(new_n945), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n947), .A2(new_n953), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n299), .A2(new_n904), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n304), .A2(new_n307), .A3(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1194), .B1(new_n304), .B2(new_n307), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1193), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1197), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1199), .A2(new_n1195), .A3(new_n1192), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  AND4_X1   g1001(.A1(G330), .A2(new_n1190), .A3(new_n1191), .A4(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1201), .B1(new_n954), .B2(G330), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n938), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT121), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1190), .A2(G330), .A3(new_n1191), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1201), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  AND3_X1   g1008(.A1(new_n928), .A2(new_n936), .A3(new_n937), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n954), .A2(G330), .A3(new_n1201), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1204), .A2(new_n1205), .A3(new_n1211), .ZN(new_n1212));
  OAI211_X1 g1012(.A(KEYINPUT121), .B(new_n938), .C1(new_n1202), .C2(new_n1203), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1148), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1162), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1214), .A2(new_n1216), .A3(KEYINPUT57), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT120), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1204), .A2(new_n1218), .A3(new_n1211), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1208), .A2(new_n1209), .A3(KEYINPUT120), .A4(new_n1210), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n1215), .B2(new_n1162), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1217), .B(new_n768), .C1(new_n1222), .C2(KEYINPUT57), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1221), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n772), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n777), .B1(new_n227), .B2(new_n843), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n793), .A2(G125), .B1(new_n1026), .B2(G150), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G132), .B2(new_n785), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n789), .A2(G137), .B1(new_n804), .B2(new_n1167), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1229), .B(new_n1230), .C1(new_n799), .C2(new_n1174), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1231), .A2(KEYINPUT59), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(KEYINPUT59), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n288), .B(new_n252), .C1(new_n809), .C2(new_n819), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(G124), .B2(new_n808), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1232), .A2(new_n1233), .A3(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n850), .B1(new_n799), .B2(new_n242), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n808), .A2(G283), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n810), .A2(G58), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1050), .A2(new_n1238), .A3(new_n1239), .A4(new_n252), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n814), .A2(new_n836), .B1(new_n781), .B2(new_n213), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n221), .A2(new_n815), .B1(new_n790), .B2(new_n442), .ZN(new_n1242));
  NOR4_X1   g1042(.A1(new_n1237), .A2(new_n1240), .A3(new_n1241), .A4(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(KEYINPUT58), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n252), .B1(new_n850), .B2(new_n288), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n227), .ZN(new_n1246));
  OR2_X1    g1046(.A1(new_n1243), .A2(KEYINPUT58), .ZN(new_n1247));
  AND4_X1   g1047(.A1(new_n1236), .A2(new_n1244), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n1226), .B1(new_n779), .B2(new_n1248), .C1(new_n1201), .C2(new_n828), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1225), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1223), .A2(new_n1250), .ZN(G375));
  INV_X1    g1051(.A(KEYINPUT124), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1156), .A2(new_n1139), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n998), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(G128), .A2(new_n808), .B1(new_n804), .B2(G159), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n815), .B2(new_n1166), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(G50), .A2(new_n1026), .B1(new_n789), .B2(G150), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n853), .B2(new_n814), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n1257), .B(new_n1259), .C1(G137), .C2(new_n800), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n831), .A2(new_n1239), .ZN(new_n1261));
  XOR2_X1   g1061(.A(new_n1261), .B(KEYINPUT122), .Z(new_n1262));
  NAND2_X1  g1062(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n815), .A2(new_n836), .B1(new_n790), .B2(new_n242), .ZN(new_n1264));
  AOI211_X1 g1064(.A(new_n1047), .B(new_n1264), .C1(G294), .C2(new_n793), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n803), .A2(new_n221), .B1(new_n807), .B2(new_n1040), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n1266), .A2(new_n262), .A3(new_n1023), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1265), .B(new_n1267), .C1(new_n1030), .C2(new_n799), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n779), .B1(new_n1263), .B2(new_n1268), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n777), .B(new_n1269), .C1(new_n213), .C2(new_n843), .ZN(new_n1270));
  XOR2_X1   g1070(.A(new_n1270), .B(KEYINPUT123), .Z(new_n1271));
  NAND2_X1  g1071(.A1(new_n1125), .A2(new_n827), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1252), .B1(new_n1255), .B2(new_n1274), .ZN(new_n1275));
  OAI211_X1 g1075(.A(KEYINPUT124), .B(new_n1273), .C1(new_n1157), .C2(new_n998), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1161), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1015), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1157), .A2(new_n1148), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1278), .A2(new_n1279), .A3(new_n1280), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1277), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(G381));
  NOR4_X1   g1083(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1284), .A2(new_n1044), .A3(new_n1018), .A4(new_n1282), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT125), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(new_n1285), .B(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(G378), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1223), .A2(new_n1250), .A3(new_n1288), .ZN(new_n1289));
  OR2_X1    g1089(.A1(new_n1287), .A2(new_n1289), .ZN(G407));
  OR2_X1    g1090(.A1(new_n1289), .A2(G343), .ZN(new_n1291));
  OAI211_X1 g1091(.A(G213), .B(new_n1291), .C1(new_n1287), .C2(new_n1289), .ZN(G409));
  NAND3_X1  g1092(.A1(G390), .A2(new_n1018), .A3(new_n1044), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(KEYINPUT127), .ZN(new_n1294));
  XOR2_X1   g1094(.A(G393), .B(G396), .Z(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(G390), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G387), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1293), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1296), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT127), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1298), .A2(new_n1301), .A3(new_n1293), .A4(new_n1295), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1300), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT126), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n761), .B1(new_n1215), .B2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT60), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1280), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1157), .A2(KEYINPUT60), .A3(new_n1148), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1306), .A2(new_n1308), .A3(new_n1309), .ZN(new_n1310));
  AND3_X1   g1110(.A1(G384), .A2(new_n1310), .A3(new_n1277), .ZN(new_n1311));
  AOI21_X1  g1111(.A(G384), .B1(new_n1277), .B2(new_n1310), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1304), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1310), .A2(new_n1277), .ZN(new_n1314));
  INV_X1    g1114(.A(G384), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(G384), .A2(new_n1310), .A3(new_n1277), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1316), .A2(KEYINPUT126), .A3(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(G213), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1319), .A2(G343), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(G2897), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1313), .A2(new_n1318), .A3(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1323), .A2(G2897), .A3(new_n1320), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1288), .B1(new_n1223), .B2(new_n1250), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1212), .A2(new_n772), .A3(new_n1213), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1163), .A2(new_n1188), .A3(new_n1249), .A4(new_n1326), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1224), .A2(new_n1279), .A3(new_n1216), .ZN(new_n1328));
  OAI22_X1  g1128(.A1(new_n1327), .A2(new_n1328), .B1(new_n1319), .B2(G343), .ZN(new_n1329));
  OAI211_X1 g1129(.A(new_n1322), .B(new_n1324), .C1(new_n1325), .C2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT61), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1313), .A2(new_n1318), .ZN(new_n1332));
  NOR3_X1   g1132(.A1(new_n1325), .A2(new_n1332), .A3(new_n1329), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT62), .ZN(new_n1334));
  OAI211_X1 g1134(.A(new_n1330), .B(new_n1331), .C1(new_n1333), .C2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(G375), .A2(G378), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1332), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1329), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1336), .A2(new_n1337), .A3(new_n1338), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1339), .A2(KEYINPUT62), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1303), .B1(new_n1335), .B2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1336), .A2(new_n1338), .ZN(new_n1342));
  AND2_X1   g1142(.A1(new_n1322), .A2(new_n1324), .ZN(new_n1343));
  AOI21_X1  g1143(.A(KEYINPUT61), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1302), .ZN(new_n1345));
  AOI22_X1  g1145(.A1(new_n1294), .A2(new_n1295), .B1(new_n1298), .B2(new_n1293), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT63), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1339), .A2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1333), .A2(KEYINPUT63), .ZN(new_n1350));
  NAND4_X1  g1150(.A1(new_n1344), .A2(new_n1347), .A3(new_n1349), .A4(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1341), .A2(new_n1351), .ZN(G405));
  AOI21_X1  g1152(.A(new_n1323), .B1(new_n1336), .B2(new_n1289), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1336), .A2(new_n1289), .ZN(new_n1355));
  OAI211_X1 g1155(.A(new_n1303), .B(new_n1354), .C1(new_n1337), .C2(new_n1355), .ZN(new_n1356));
  NOR2_X1   g1156(.A1(new_n1355), .A2(new_n1337), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1347), .B1(new_n1357), .B2(new_n1353), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1356), .A2(new_n1358), .ZN(G402));
endmodule


