//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 0 1 0 0 1 0 1 0 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011;
  INV_X1    g000(.A(G137), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT65), .B1(new_n187), .B2(G134), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT65), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G137), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G131), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT11), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n194), .B1(new_n190), .B2(G137), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n187), .A2(KEYINPUT11), .A3(G134), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n192), .A2(new_n193), .A3(new_n195), .A4(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n190), .A2(G137), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n187), .A2(G134), .ZN(new_n199));
  OAI21_X1  g013(.A(G131), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT1), .B1(new_n204), .B2(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT67), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT68), .A2(G128), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT68), .A2(G128), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT67), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT1), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n206), .A2(new_n209), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n204), .A2(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n211), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(G143), .B(G146), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT1), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(G128), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n197), .A2(KEYINPUT66), .A3(new_n200), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n203), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT30), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n192), .A2(new_n195), .A3(new_n196), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G131), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n197), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT0), .B(G128), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT64), .B1(new_n218), .B2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n218), .A2(KEYINPUT0), .A3(G128), .ZN(new_n230));
  INV_X1    g044(.A(G128), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT0), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT0), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G128), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT64), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n216), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n229), .A2(new_n230), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n227), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n223), .A2(new_n224), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n238), .B1(new_n226), .B2(new_n197), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n216), .A2(new_n231), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n214), .A2(new_n216), .B1(new_n243), .B2(new_n219), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(new_n201), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT30), .B1(new_n242), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  AND2_X1   g061(.A1(KEYINPUT69), .A2(G119), .ZN(new_n248));
  NOR2_X1   g062(.A1(KEYINPUT69), .A2(G119), .ZN(new_n249));
  OAI21_X1  g063(.A(G116), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G116), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT71), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G116), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G119), .ZN(new_n258));
  OAI211_X1 g072(.A(KEYINPUT70), .B(G116), .C1(new_n248), .C2(new_n249), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n252), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT2), .B(G113), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n261), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n252), .A2(new_n258), .A3(new_n263), .A4(new_n259), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n262), .A2(KEYINPUT72), .A3(new_n264), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n247), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n268), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT72), .B1(new_n262), .B2(new_n264), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n221), .A2(new_n197), .A3(new_n200), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(new_n240), .A3(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(G237), .A2(G953), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G210), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n279), .B(G101), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n280), .B(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n247), .A2(KEYINPUT73), .A3(new_n269), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n272), .A2(new_n277), .A3(new_n282), .A4(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT31), .ZN(new_n285));
  AOI221_X4 g099(.A(new_n271), .B1(new_n267), .B2(new_n268), .C1(new_n241), .C2(new_n246), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT73), .B1(new_n247), .B2(new_n269), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT31), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n288), .A2(new_n289), .A3(new_n277), .A4(new_n282), .ZN(new_n290));
  XOR2_X1   g104(.A(new_n282), .B(KEYINPUT74), .Z(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n276), .A2(new_n240), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT75), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n276), .A2(new_n240), .A3(KEYINPUT75), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(new_n275), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT28), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n223), .A2(new_n240), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n269), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n298), .B1(new_n277), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n292), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n285), .A2(new_n290), .A3(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(G472), .A2(G902), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT32), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n305), .A2(KEYINPUT32), .A3(new_n306), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n272), .A2(new_n277), .A3(new_n283), .ZN(new_n311));
  INV_X1    g125(.A(new_n282), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT29), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n269), .A2(new_n293), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n315), .B1(new_n269), .B2(new_n301), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n299), .B(new_n291), .C1(new_n316), .C2(new_n298), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n313), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  AOI22_X1  g132(.A1(new_n267), .A2(new_n268), .B1(new_n240), .B2(new_n276), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT28), .B1(new_n315), .B2(new_n319), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n320), .A2(new_n299), .A3(KEYINPUT29), .A4(new_n282), .ZN(new_n321));
  INV_X1    g135(.A(G902), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G472), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n309), .A2(new_n310), .A3(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT25), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT22), .B(G137), .ZN(new_n328));
  INV_X1    g142(.A(G221), .ZN(new_n329));
  INV_X1    g143(.A(G234), .ZN(new_n330));
  NOR3_X1   g144(.A1(new_n329), .A2(new_n330), .A3(G953), .ZN(new_n331));
  XOR2_X1   g145(.A(new_n328), .B(new_n331), .Z(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT69), .B(G119), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n334), .B1(new_n335), .B2(G128), .ZN(new_n336));
  OAI21_X1  g150(.A(G128), .B1(new_n248), .B2(new_n249), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT23), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n248), .A2(new_n249), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(KEYINPUT77), .A3(new_n231), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n336), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G110), .ZN(new_n342));
  OAI211_X1 g156(.A(KEYINPUT23), .B(G119), .C1(new_n207), .C2(new_n208), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G119), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n337), .B1(new_n209), .B2(new_n347), .ZN(new_n348));
  XOR2_X1   g162(.A(KEYINPUT24), .B(G110), .Z(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n341), .A2(KEYINPUT78), .A3(new_n342), .A4(new_n343), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n346), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G125), .ZN(new_n354));
  NOR3_X1   g168(.A1(new_n354), .A2(KEYINPUT16), .A3(G140), .ZN(new_n355));
  XNOR2_X1  g169(.A(G125), .B(G140), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n355), .B1(new_n356), .B2(KEYINPUT16), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G146), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n210), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n353), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n356), .A2(KEYINPUT16), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n210), .B1(new_n363), .B2(new_n355), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n358), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n341), .A2(new_n343), .ZN(new_n366));
  OAI221_X1 g180(.A(new_n365), .B1(new_n348), .B2(new_n350), .C1(new_n366), .C2(new_n342), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n361), .A2(new_n362), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n362), .B1(new_n361), .B2(new_n367), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n333), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n361), .A2(new_n367), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(new_n333), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n327), .B1(new_n375), .B2(G902), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n372), .A2(KEYINPUT79), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n368), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n373), .B1(new_n378), .B2(new_n333), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(KEYINPUT25), .A3(new_n322), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G217), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n382), .B1(G234), .B2(new_n322), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n383), .B(KEYINPUT76), .ZN(new_n384));
  INV_X1    g198(.A(new_n383), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n322), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(KEYINPUT80), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  AOI22_X1  g202(.A1(new_n381), .A2(new_n384), .B1(new_n388), .B2(new_n379), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n326), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G122), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n391), .B1(new_n254), .B2(new_n256), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(KEYINPUT95), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT95), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G122), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n253), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  OR2_X1    g210(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(G107), .ZN(new_n398));
  OAI21_X1  g212(.A(G143), .B1(new_n207), .B2(new_n208), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n204), .A2(G128), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n209), .A2(new_n204), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n401), .B(G134), .C1(new_n402), .C2(KEYINPUT13), .ZN(new_n403));
  NAND2_X1  g217(.A1(KEYINPUT13), .A2(G134), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n399), .A2(new_n400), .A3(new_n404), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n398), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT97), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT96), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT14), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n410), .B1(new_n257), .B2(G122), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n409), .B1(new_n411), .B2(new_n396), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n392), .A2(new_n410), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n393), .A2(new_n395), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G116), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n415), .B(KEYINPUT96), .C1(new_n392), .C2(new_n410), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n412), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(G107), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n397), .A2(G107), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n401), .B(G134), .ZN(new_n421));
  AND4_X1   g235(.A1(new_n408), .A2(new_n418), .A3(new_n420), .A4(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n419), .B1(new_n417), .B2(G107), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n408), .B1(new_n423), .B2(new_n421), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n407), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  XOR2_X1   g239(.A(KEYINPUT9), .B(G234), .Z(new_n426));
  INV_X1    g240(.A(G953), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(G217), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n418), .A2(new_n420), .A3(new_n421), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT97), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n423), .A2(new_n408), .A3(new_n421), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(new_n407), .A3(new_n428), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n430), .A2(new_n435), .A3(new_n322), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT98), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G478), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n439), .A2(KEYINPUT15), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n430), .A2(new_n435), .A3(KEYINPUT98), .A4(new_n322), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  OR2_X1    g256(.A1(new_n436), .A2(new_n440), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT92), .B(G475), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT93), .ZN(new_n447));
  INV_X1    g261(.A(G237), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(new_n427), .A3(G214), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n204), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n278), .A2(G143), .A3(G214), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(KEYINPUT18), .A3(G131), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n356), .B(new_n210), .ZN(new_n454));
  NAND2_X1  g268(.A1(KEYINPUT18), .A2(G131), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n450), .A2(new_n451), .A3(new_n455), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n456), .A2(KEYINPUT90), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n456), .A2(KEYINPUT90), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n453), .B(new_n454), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n278), .A2(G143), .A3(G214), .ZN(new_n460));
  AOI21_X1  g274(.A(G143), .B1(new_n278), .B2(G214), .ZN(new_n461));
  OAI21_X1  g275(.A(G131), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT17), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n450), .A2(new_n193), .A3(new_n451), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n452), .A2(KEYINPUT17), .A3(G131), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n465), .A2(new_n364), .A3(new_n358), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n459), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(G113), .B(G122), .ZN(new_n469));
  INV_X1    g283(.A(G104), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n469), .B(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n447), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  AOI211_X1 g287(.A(KEYINPUT93), .B(new_n471), .C1(new_n459), .C2(new_n467), .ZN(new_n474));
  OAI22_X1  g288(.A1(new_n473), .A2(new_n474), .B1(new_n472), .B2(new_n468), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT94), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n475), .A2(new_n476), .A3(new_n322), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n476), .B1(new_n475), .B2(new_n322), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n446), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n468), .A2(new_n472), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n462), .A2(new_n464), .ZN(new_n481));
  XOR2_X1   g295(.A(new_n356), .B(KEYINPUT19), .Z(new_n482));
  OAI211_X1 g296(.A(new_n358), .B(new_n481), .C1(new_n482), .C2(G146), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n471), .B1(new_n459), .B2(new_n483), .ZN(new_n484));
  OR2_X1    g298(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(G475), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n486), .A3(new_n322), .ZN(new_n487));
  NAND2_X1  g301(.A1(KEYINPUT91), .A2(KEYINPUT20), .ZN(new_n488));
  OR2_X1    g302(.A1(KEYINPUT91), .A2(KEYINPUT20), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  OR2_X1    g304(.A1(new_n487), .A2(new_n488), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n479), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n444), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(G214), .B1(G237), .B2(G902), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n244), .A2(new_n354), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n238), .A2(G125), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G224), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n499), .A2(G953), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n498), .B(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT6), .ZN(new_n502));
  XOR2_X1   g316(.A(G110), .B(G122), .Z(new_n503));
  XOR2_X1   g317(.A(new_n503), .B(KEYINPUT86), .Z(new_n504));
  OAI21_X1  g318(.A(KEYINPUT3), .B1(new_n470), .B2(G107), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT3), .ZN(new_n506));
  INV_X1    g320(.A(G107), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n507), .A3(G104), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n470), .A2(G107), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n505), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(G101), .ZN(new_n511));
  INV_X1    g325(.A(G101), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n505), .A2(new_n508), .A3(new_n512), .A4(new_n509), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT81), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n513), .A2(new_n514), .ZN(new_n516));
  OAI211_X1 g330(.A(KEYINPUT4), .B(new_n511), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n511), .A2(KEYINPUT4), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n520), .B1(new_n267), .B2(new_n268), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT5), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n335), .A2(new_n522), .A3(G116), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n523), .B(G113), .C1(new_n260), .C2(new_n522), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT82), .B1(new_n507), .B2(G104), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n507), .A2(G104), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n507), .A2(KEYINPUT82), .A3(G104), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n512), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AND2_X1   g343(.A1(new_n505), .A2(new_n508), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n530), .A2(KEYINPUT81), .A3(new_n512), .A4(new_n509), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n513), .A2(new_n514), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n524), .A2(new_n264), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n504), .B1(new_n521), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT4), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n537), .B1(new_n531), .B2(new_n532), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n518), .B1(new_n538), .B2(new_n511), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n539), .B1(new_n273), .B2(new_n274), .ZN(new_n540));
  INV_X1    g354(.A(new_n503), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n534), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n502), .B1(new_n536), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n540), .A2(new_n534), .ZN(new_n544));
  AOI21_X1  g358(.A(KEYINPUT6), .B1(new_n544), .B2(new_n504), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n501), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n500), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT7), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n547), .B1(KEYINPUT87), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n549), .B1(KEYINPUT87), .B2(new_n548), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n550), .B1(new_n496), .B2(new_n497), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT88), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n498), .B1(new_n552), .B2(new_n500), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n548), .B1(new_n547), .B2(KEYINPUT88), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n551), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  XOR2_X1   g369(.A(new_n503), .B(KEYINPUT8), .Z(new_n556));
  AOI21_X1  g370(.A(new_n533), .B1(new_n524), .B2(new_n264), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n556), .B1(new_n535), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n555), .A2(new_n542), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n546), .A2(new_n322), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT89), .ZN(new_n561));
  OAI21_X1  g375(.A(G210), .B1(G237), .B2(G902), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n561), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n546), .A2(new_n322), .A3(new_n559), .A4(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n495), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n329), .B1(new_n426), .B2(new_n322), .ZN(new_n568));
  INV_X1    g382(.A(G469), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n569), .A2(new_n322), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n517), .A2(new_n239), .A3(new_n519), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n527), .A2(new_n528), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G101), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n231), .B1(new_n211), .B2(KEYINPUT1), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n220), .B1(new_n574), .B2(new_n218), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n573), .B(new_n575), .C1(new_n515), .C2(new_n516), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT10), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n227), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n577), .B1(new_n217), .B2(new_n220), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n533), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n571), .A2(new_n578), .A3(new_n579), .A4(new_n581), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n577), .A2(new_n576), .B1(new_n580), .B2(new_n533), .ZN(new_n583));
  AOI211_X1 g397(.A(KEYINPUT85), .B(new_n579), .C1(new_n583), .C2(new_n571), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT85), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n571), .A2(new_n578), .A3(new_n581), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n585), .B1(new_n586), .B2(new_n227), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n582), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(G110), .B(G140), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n427), .A2(G227), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT12), .B1(new_n227), .B2(KEYINPUT83), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n576), .B1(new_n533), .B2(new_n221), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n594), .B1(new_n596), .B2(new_n579), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n595), .B(new_n227), .C1(KEYINPUT83), .C2(KEYINPUT12), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n582), .A2(new_n591), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(G902), .B1(new_n593), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n570), .B1(new_n603), .B2(new_n569), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n591), .B1(new_n599), .B2(new_n582), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n586), .A2(new_n227), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT85), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n586), .A2(new_n585), .A3(new_n227), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n582), .A2(KEYINPUT84), .A3(new_n591), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT84), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n600), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n606), .A2(new_n614), .A3(G469), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n568), .B1(new_n604), .B2(new_n615), .ZN(new_n616));
  OR2_X1    g430(.A1(KEYINPUT99), .A2(G952), .ZN(new_n617));
  NAND2_X1  g431(.A1(KEYINPUT99), .A2(G952), .ZN(new_n618));
  AOI21_X1  g432(.A(G953), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n619), .B1(new_n330), .B2(new_n448), .ZN(new_n620));
  AOI211_X1 g434(.A(new_n322), .B(new_n427), .C1(G234), .C2(G237), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT21), .B(G898), .Z(new_n623));
  OAI21_X1  g437(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n493), .A2(new_n567), .A3(new_n616), .A4(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n390), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(new_n512), .ZN(G3));
  INV_X1    g441(.A(KEYINPUT101), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n305), .A2(new_n322), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(G472), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT100), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(G472), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n305), .B2(new_n322), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(KEYINPUT100), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n632), .A2(new_n307), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n389), .A2(new_n616), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n628), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT100), .B1(new_n629), .B2(G472), .ZN(new_n639));
  AOI211_X1 g453(.A(new_n631), .B(new_n633), .C1(new_n305), .C2(new_n322), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(KEYINPUT25), .B1(new_n379), .B2(new_n322), .ZN(new_n642));
  AND4_X1   g456(.A1(KEYINPUT25), .A2(new_n371), .A3(new_n322), .A4(new_n374), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n384), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n379), .A2(new_n388), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n591), .B1(new_n610), .B2(new_n582), .ZN(new_n647));
  INV_X1    g461(.A(new_n602), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n569), .B(new_n322), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n570), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n649), .A2(new_n650), .A3(new_n615), .ZN(new_n651));
  INV_X1    g465(.A(new_n568), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n641), .A2(new_n654), .A3(KEYINPUT101), .A4(new_n307), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n429), .A2(KEYINPUT103), .ZN(new_n656));
  AOI21_X1  g470(.A(KEYINPUT102), .B1(new_n656), .B2(KEYINPUT33), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(KEYINPUT102), .B2(KEYINPUT33), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n430), .A2(new_n435), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n657), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n661), .B1(new_n430), .B2(new_n435), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n322), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(G478), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n438), .A2(new_n441), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n439), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT104), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n664), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n428), .B1(new_n434), .B2(new_n407), .ZN(new_n669));
  AOI211_X1 g483(.A(new_n429), .B(new_n406), .C1(new_n432), .C2(new_n433), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n657), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n659), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n439), .B1(new_n672), .B2(new_n322), .ZN(new_n673));
  AOI21_X1  g487(.A(G478), .B1(new_n438), .B2(new_n441), .ZN(new_n674));
  OAI21_X1  g488(.A(KEYINPUT104), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n668), .A2(new_n675), .A3(new_n492), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n560), .A2(new_n562), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n546), .A2(new_n322), .A3(new_n559), .A4(new_n563), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n677), .A2(new_n494), .A3(new_n624), .A4(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n638), .A2(new_n655), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT34), .B(G104), .Z(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT105), .B(KEYINPUT106), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n681), .B(new_n684), .ZN(G6));
  AND3_X1   g499(.A1(new_n677), .A2(new_n494), .A3(new_n678), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n492), .B1(new_n443), .B2(new_n442), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n686), .A2(new_n687), .A3(new_n688), .A4(new_n624), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n479), .A2(new_n490), .A3(new_n491), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n444), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g505(.A(KEYINPUT107), .B1(new_n691), .B2(new_n679), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n638), .A2(new_n655), .A3(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT35), .B(G107), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G9));
  NOR2_X1   g510(.A1(new_n636), .A2(new_n625), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n333), .A2(KEYINPUT36), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n378), .B(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n644), .B1(new_n387), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G110), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT108), .B(KEYINPUT37), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G12));
  AND3_X1   g519(.A1(new_n305), .A2(KEYINPUT32), .A3(new_n306), .ZN(new_n706));
  AOI21_X1  g520(.A(KEYINPUT32), .B1(new_n305), .B2(new_n306), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n653), .B1(new_n708), .B2(new_n325), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n620), .B1(new_n622), .B2(G900), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n687), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n709), .A2(new_n686), .A3(new_n701), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G128), .ZN(G30));
  NAND2_X1  g527(.A1(new_n564), .A2(new_n566), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT38), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n444), .A2(new_n494), .A3(new_n492), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT40), .ZN(new_n719));
  XOR2_X1   g533(.A(new_n710), .B(KEYINPUT39), .Z(new_n720));
  NOR2_X1   g534(.A1(new_n653), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n718), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n292), .B1(new_n315), .B2(new_n319), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n284), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g538(.A(G472), .B1(new_n724), .B2(G902), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n701), .B1(new_n708), .B2(new_n725), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n722), .B(new_n726), .C1(new_n719), .C2(new_n721), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G143), .ZN(G45));
  NAND4_X1  g542(.A1(new_n668), .A2(new_n675), .A3(new_n492), .A4(new_n710), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n730), .A2(new_n709), .A3(new_n686), .A4(new_n701), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G146), .ZN(G48));
  AOI22_X1  g546(.A1(new_n588), .A2(new_n592), .B1(new_n601), .B2(new_n599), .ZN(new_n733));
  OAI21_X1  g547(.A(G469), .B1(new_n733), .B2(G902), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n649), .A3(new_n652), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n326), .A2(new_n389), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n680), .ZN(new_n738));
  XNOR2_X1  g552(.A(KEYINPUT41), .B(G113), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G15));
  NAND2_X1  g554(.A1(new_n737), .A2(new_n693), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G116), .ZN(G18));
  NAND3_X1  g556(.A1(new_n686), .A2(KEYINPUT109), .A3(new_n736), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n677), .A2(new_n494), .A3(new_n678), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n744), .B1(new_n745), .B2(new_n735), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n493), .A2(new_n624), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n747), .A2(new_n326), .A3(new_n748), .A4(new_n701), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G119), .ZN(G21));
  NAND2_X1  g564(.A1(new_n320), .A2(new_n299), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n291), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n320), .A2(new_n299), .A3(KEYINPUT110), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n285), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(KEYINPUT111), .ZN(new_n757));
  AOI22_X1  g571(.A1(new_n753), .A2(new_n754), .B1(KEYINPUT31), .B2(new_n284), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n757), .A2(new_n760), .A3(new_n290), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n634), .B1(new_n761), .B2(new_n306), .ZN(new_n762));
  INV_X1    g576(.A(new_n679), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n736), .A2(new_n444), .A3(new_n492), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n762), .A2(new_n389), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G122), .ZN(G24));
  NAND4_X1  g580(.A1(new_n730), .A2(new_n747), .A3(new_n701), .A4(new_n762), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G125), .ZN(G27));
  XNOR2_X1  g582(.A(KEYINPUT114), .B(KEYINPUT42), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n668), .A2(new_n675), .A3(new_n492), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n649), .A2(new_n650), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n613), .A2(new_n611), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n584), .A2(new_n587), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT112), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n610), .A2(new_n775), .A3(new_n611), .A4(new_n613), .ZN(new_n776));
  AOI211_X1 g590(.A(new_n569), .B(new_n605), .C1(new_n774), .C2(new_n776), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT113), .B1(new_n771), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n605), .B1(new_n774), .B2(new_n776), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(G469), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n604), .A3(new_n781), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n778), .A2(new_n782), .A3(new_n652), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n564), .A2(new_n566), .A3(new_n494), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n770), .A2(new_n783), .A3(new_n710), .A4(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n769), .B1(new_n786), .B2(new_n390), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT115), .B1(new_n309), .B2(new_n310), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n325), .B1(new_n706), .B2(new_n789), .ZN(new_n790));
  OAI211_X1 g604(.A(KEYINPUT42), .B(new_n389), .C1(new_n788), .C2(new_n790), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n786), .A2(KEYINPUT116), .A3(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n778), .A2(new_n782), .A3(new_n652), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n729), .A2(new_n794), .A3(new_n784), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT42), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n789), .B1(new_n706), .B2(new_n707), .ZN(new_n797));
  AOI22_X1  g611(.A1(new_n310), .A2(KEYINPUT115), .B1(new_n324), .B2(G472), .ZN(new_n798));
  AOI211_X1 g612(.A(new_n796), .B(new_n646), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n793), .B1(new_n795), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n787), .B1(new_n792), .B2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G131), .ZN(G33));
  NOR2_X1   g616(.A1(new_n390), .A2(new_n784), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n803), .A2(new_n711), .A3(new_n783), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G134), .ZN(G36));
  NAND3_X1  g619(.A1(new_n668), .A2(new_n675), .A3(new_n690), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT43), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n806), .B1(KEYINPUT118), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(KEYINPUT118), .B(KEYINPUT43), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n808), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n810), .A2(new_n701), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n636), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT44), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n811), .A2(KEYINPUT44), .A3(new_n636), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n614), .A2(new_n606), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n816), .A2(KEYINPUT45), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n779), .A2(new_n818), .A3(KEYINPUT45), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n818), .B1(new_n779), .B2(KEYINPUT45), .ZN(new_n820));
  OAI211_X1 g634(.A(G469), .B(new_n817), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n650), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT46), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n821), .A2(KEYINPUT46), .A3(new_n650), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n824), .A2(new_n649), .A3(new_n825), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n826), .A2(new_n568), .A3(new_n720), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n814), .A2(new_n785), .A3(new_n815), .A4(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(G137), .ZN(G39));
  INV_X1    g643(.A(new_n326), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n729), .A2(new_n389), .A3(new_n784), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n826), .A2(new_n568), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT47), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n832), .A2(KEYINPUT47), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n830), .B(new_n831), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(G140), .ZN(G42));
  AOI21_X1  g651(.A(new_n646), .B1(new_n797), .B2(new_n798), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n784), .A2(new_n620), .A3(new_n735), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n810), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT48), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(KEYINPUT120), .ZN(new_n842));
  XOR2_X1   g656(.A(new_n840), .B(new_n842), .Z(new_n843));
  OAI21_X1  g657(.A(new_n843), .B1(KEYINPUT120), .B2(new_n841), .ZN(new_n844));
  INV_X1    g658(.A(new_n620), .ZN(new_n845));
  INV_X1    g659(.A(new_n760), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n290), .B1(new_n758), .B2(new_n759), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n306), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n630), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n646), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n810), .A2(new_n845), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n747), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n844), .A2(new_n619), .A3(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n835), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n734), .A2(new_n649), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n568), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n854), .A2(new_n833), .A3(new_n856), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n857), .A2(new_n785), .A3(new_n851), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n811), .A2(new_n762), .A3(new_n839), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n715), .A2(new_n494), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n851), .A2(new_n736), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT50), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n851), .A2(KEYINPUT50), .A3(new_n736), .A4(new_n860), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n859), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n708), .A2(new_n389), .A3(new_n725), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n866), .A2(new_n839), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n668), .A2(new_n675), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n867), .A2(new_n690), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT51), .B1(new_n858), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n857), .A2(new_n785), .A3(new_n851), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT51), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n872), .A2(new_n873), .A3(new_n869), .A4(new_n865), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n853), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n867), .A2(new_n770), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n801), .A2(new_n804), .ZN(new_n878));
  AND4_X1   g692(.A1(new_n738), .A2(new_n749), .A3(new_n741), .A4(new_n765), .ZN(new_n879));
  INV_X1    g693(.A(new_n390), .ZN(new_n880));
  INV_X1    g694(.A(new_n625), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n697), .A2(new_n701), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n567), .A2(new_n624), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n883), .B1(new_n676), .B2(new_n691), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n638), .A2(new_n655), .A3(new_n884), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n849), .A2(new_n729), .A3(new_n794), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT119), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n493), .A2(new_n887), .A3(new_n710), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n690), .A2(new_n443), .A3(new_n442), .A4(new_n710), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT119), .ZN(new_n890));
  AND4_X1   g704(.A1(new_n326), .A2(new_n888), .A3(new_n616), .A4(new_n890), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n701), .B(new_n785), .C1(new_n886), .C2(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n879), .A2(new_n882), .A3(new_n885), .A4(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n878), .A2(new_n893), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n767), .A2(new_n712), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT52), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n677), .A2(new_n678), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n716), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n726), .A2(new_n710), .A3(new_n783), .A4(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n895), .A2(new_n896), .A3(new_n731), .A4(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n767), .A2(new_n731), .A3(new_n712), .A4(new_n899), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT52), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT53), .B1(new_n894), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n882), .A2(new_n885), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n738), .A2(new_n749), .A3(new_n741), .A4(new_n765), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n908), .A2(new_n801), .A3(new_n804), .A4(new_n892), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT53), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n909), .A2(new_n910), .A3(new_n903), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n877), .B1(new_n905), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n894), .A2(new_n904), .A3(KEYINPUT53), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n910), .B1(new_n909), .B2(new_n903), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n914), .A3(KEYINPUT54), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n875), .A2(new_n876), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n917), .B1(G952), .B2(G953), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n715), .A2(new_n495), .A3(new_n568), .ZN(new_n919));
  INV_X1    g733(.A(new_n806), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n855), .B(KEYINPUT49), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n919), .A2(new_n920), .A3(new_n866), .A4(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n918), .A2(new_n922), .ZN(G75));
  INV_X1    g737(.A(KEYINPUT56), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n913), .A2(new_n914), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(G902), .ZN(new_n926));
  INV_X1    g740(.A(G210), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n543), .A2(new_n545), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(new_n501), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT55), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n928), .A2(new_n931), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n427), .A2(G952), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT121), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n932), .A2(new_n933), .A3(new_n935), .ZN(G51));
  XNOR2_X1  g750(.A(new_n570), .B(KEYINPUT57), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n912), .A2(new_n915), .A3(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n733), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n938), .A2(KEYINPUT122), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT122), .B1(new_n938), .B2(new_n939), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n926), .A2(new_n821), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n934), .B1(new_n942), .B2(new_n943), .ZN(G54));
  INV_X1    g758(.A(KEYINPUT58), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT123), .B1(new_n945), .B2(new_n486), .ZN(new_n946));
  OR3_X1    g760(.A1(new_n945), .A2(new_n486), .A3(KEYINPUT123), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n925), .A2(G902), .A3(new_n946), .A4(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n485), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n948), .A2(new_n949), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n950), .A2(new_n951), .A3(new_n934), .ZN(G60));
  NAND2_X1  g766(.A1(G478), .A2(G902), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT59), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n912), .A2(new_n915), .A3(new_n954), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n672), .B(KEYINPUT124), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n955), .A2(new_n956), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n957), .A2(new_n958), .A3(new_n935), .ZN(G63));
  NOR2_X1   g773(.A1(new_n905), .A2(new_n911), .ZN(new_n960));
  NAND2_X1  g774(.A1(G217), .A2(G902), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT60), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n935), .B1(new_n963), .B2(new_n699), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n375), .B1(new_n960), .B2(new_n962), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT61), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n964), .A2(KEYINPUT61), .A3(new_n965), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(G66));
  INV_X1    g784(.A(new_n908), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n427), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT125), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n427), .B1(new_n623), .B2(G224), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(G898), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n929), .B1(new_n976), .B2(G953), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n975), .B(new_n977), .ZN(G69));
  XNOR2_X1  g792(.A(new_n247), .B(new_n482), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(G900), .A2(G953), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n838), .A2(new_n898), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n878), .B1(new_n827), .B2(new_n982), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n895), .A2(new_n731), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n836), .A2(new_n983), .A3(new_n828), .A4(new_n984), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n980), .B(new_n981), .C1(new_n985), .C2(G953), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n984), .A2(new_n727), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT62), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n984), .A2(KEYINPUT62), .A3(new_n727), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n803), .B(new_n721), .C1(new_n770), .C2(new_n687), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n991), .A2(new_n828), .A3(new_n836), .A4(new_n992), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n993), .A2(new_n427), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n986), .B1(new_n994), .B2(new_n980), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n427), .B1(G227), .B2(G900), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n995), .B(new_n996), .ZN(G72));
  NAND2_X1  g811(.A1(G472), .A2(G902), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT63), .Z(new_n999));
  OAI21_X1  g813(.A(new_n999), .B1(new_n985), .B2(new_n971), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n311), .B(KEYINPUT127), .Z(new_n1001));
  NAND3_X1  g815(.A1(new_n1000), .A2(new_n312), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n313), .A2(new_n284), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n925), .A2(new_n999), .A3(new_n1003), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n1002), .B(new_n1004), .C1(G952), .C2(new_n427), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n999), .B1(new_n993), .B2(new_n971), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT126), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1001), .ZN(new_n1009));
  OAI211_X1 g823(.A(KEYINPUT126), .B(new_n999), .C1(new_n993), .C2(new_n971), .ZN(new_n1010));
  AND3_X1   g824(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1005), .B1(new_n1011), .B2(new_n282), .ZN(G57));
endmodule


