

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766;

  AND2_X1 U377 ( .A1(n646), .A2(KEYINPUT68), .ZN(n439) );
  XNOR2_X1 U378 ( .A(n544), .B(KEYINPUT32), .ZN(n658) );
  INV_X1 U379 ( .A(n583), .ZN(n701) );
  BUF_X1 U380 ( .A(G107), .Z(n357) );
  NAND2_X1 U381 ( .A1(n358), .A2(n437), .ZN(n446) );
  NAND2_X1 U382 ( .A1(n439), .A2(n364), .ZN(n358) );
  NOR2_X2 U383 ( .A1(n592), .A2(n709), .ZN(n469) );
  XNOR2_X2 U384 ( .A(n467), .B(n466), .ZN(n592) );
  NOR2_X1 U385 ( .A1(G953), .A2(G237), .ZN(n526) );
  NOR2_X1 U386 ( .A1(n612), .A2(n613), .ZN(n742) );
  AND2_X1 U387 ( .A1(n388), .A2(n387), .ZN(n359) );
  XNOR2_X2 U388 ( .A(n560), .B(n559), .ZN(n424) );
  AND2_X4 U389 ( .A1(n444), .A2(n443), .ZN(n683) );
  XNOR2_X2 U390 ( .A(n429), .B(n369), .ZN(n547) );
  XNOR2_X2 U391 ( .A(n553), .B(n552), .ZN(n407) );
  NOR2_X1 U392 ( .A1(n545), .A2(n696), .ZN(n409) );
  INV_X2 U393 ( .A(G953), .ZN(n755) );
  XNOR2_X1 U394 ( .A(n379), .B(n413), .ZN(n633) );
  NOR2_X1 U395 ( .A1(n598), .A2(n726), .ZN(n599) );
  XNOR2_X1 U396 ( .A(n409), .B(n408), .ZN(n394) );
  XNOR2_X1 U397 ( .A(G104), .B(G107), .ZN(n449) );
  NAND2_X1 U398 ( .A1(n633), .A2(n626), .ZN(n647) );
  NAND2_X1 U399 ( .A1(n396), .A2(n542), .ZN(n657) );
  NAND2_X1 U400 ( .A1(n394), .A2(n604), .ZN(n429) );
  BUF_X1 U401 ( .A(n545), .Z(n525) );
  OR2_X1 U402 ( .A1(n710), .A2(n709), .ZN(n382) );
  XNOR2_X1 U403 ( .A(n660), .B(KEYINPUT125), .ZN(n661) );
  AND2_X1 U404 ( .A1(n393), .A2(n392), .ZN(n391) );
  XNOR2_X1 U405 ( .A(n665), .B(KEYINPUT123), .ZN(n666) );
  XNOR2_X1 U406 ( .A(n672), .B(n671), .ZN(n673) );
  INV_X1 U407 ( .A(n449), .ZN(n451) );
  BUF_X1 U408 ( .A(n546), .Z(n562) );
  INV_X1 U409 ( .A(n404), .ZN(n360) );
  AND2_X1 U410 ( .A1(n565), .A2(n657), .ZN(n405) );
  NAND2_X1 U411 ( .A1(n381), .A2(n600), .ZN(n380) );
  INV_X1 U412 ( .A(n763), .ZN(n381) );
  NAND2_X1 U413 ( .A1(G469), .A2(n390), .ZN(n389) );
  NAND2_X1 U414 ( .A1(n524), .A2(G902), .ZN(n392) );
  INV_X1 U415 ( .A(KEYINPUT75), .ZN(n408) );
  XNOR2_X1 U416 ( .A(KEYINPUT18), .B(KEYINPUT94), .ZN(n452) );
  NAND2_X1 U417 ( .A1(n438), .A2(KEYINPUT44), .ZN(n437) );
  AND2_X1 U418 ( .A1(n431), .A2(n367), .ZN(n415) );
  XNOR2_X1 U419 ( .A(n380), .B(n432), .ZN(n431) );
  INV_X1 U420 ( .A(G237), .ZN(n463) );
  NAND2_X1 U421 ( .A1(n391), .A2(n388), .ZN(n385) );
  XNOR2_X1 U422 ( .A(n376), .B(n375), .ZN(n374) );
  XNOR2_X1 U423 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n376) );
  XNOR2_X1 U424 ( .A(G119), .B(G128), .ZN(n375) );
  XNOR2_X1 U425 ( .A(n373), .B(KEYINPUT82), .ZN(n372) );
  XNOR2_X1 U426 ( .A(G137), .B(G110), .ZN(n373) );
  XNOR2_X1 U427 ( .A(n378), .B(n482), .ZN(n535) );
  XNOR2_X1 U428 ( .A(n481), .B(n480), .ZN(n378) );
  INV_X1 U429 ( .A(G125), .ZN(n457) );
  XNOR2_X1 U430 ( .A(KEYINPUT67), .B(G101), .ZN(n529) );
  XNOR2_X1 U431 ( .A(n395), .B(n361), .ZN(n410) );
  INV_X1 U432 ( .A(KEYINPUT83), .ZN(n430) );
  XNOR2_X1 U433 ( .A(n416), .B(KEYINPUT110), .ZN(n598) );
  INV_X1 U434 ( .A(n584), .ZN(n417) );
  XNOR2_X1 U435 ( .A(n420), .B(n419), .ZN(n418) );
  INV_X1 U436 ( .A(KEYINPUT64), .ZN(n438) );
  NAND2_X1 U437 ( .A1(n397), .A2(n608), .ZN(n565) );
  INV_X1 U438 ( .A(n733), .ZN(n422) );
  INV_X1 U439 ( .A(KEYINPUT46), .ZN(n432) );
  INV_X1 U440 ( .A(n746), .ZN(n433) );
  AND2_X1 U441 ( .A1(n570), .A2(n426), .ZN(n425) );
  NAND2_X1 U442 ( .A1(KEYINPUT44), .A2(KEYINPUT64), .ZN(n426) );
  XNOR2_X1 U443 ( .A(KEYINPUT97), .B(KEYINPUT5), .ZN(n527) );
  XNOR2_X1 U444 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n453) );
  INV_X1 U445 ( .A(KEYINPUT48), .ZN(n413) );
  NAND2_X1 U446 ( .A1(n415), .A2(n414), .ZN(n379) );
  XNOR2_X1 U447 ( .A(n618), .B(KEYINPUT81), .ZN(n414) );
  NAND2_X1 U448 ( .A1(G234), .A2(G237), .ZN(n470) );
  NOR2_X1 U449 ( .A1(n713), .A2(n382), .ZN(n714) );
  INV_X1 U450 ( .A(n709), .ZN(n436) );
  INV_X1 U451 ( .A(KEYINPUT28), .ZN(n419) );
  NAND2_X1 U452 ( .A1(n385), .A2(KEYINPUT1), .ZN(n384) );
  NAND2_X1 U453 ( .A1(n410), .A2(n580), .ZN(n696) );
  XNOR2_X1 U454 ( .A(n537), .B(n536), .ZN(n659) );
  XNOR2_X1 U455 ( .A(n377), .B(n371), .ZN(n537) );
  XNOR2_X1 U456 ( .A(n374), .B(n372), .ZN(n371) );
  XOR2_X1 U457 ( .A(n357), .B(G122), .Z(n485) );
  XNOR2_X1 U458 ( .A(KEYINPUT107), .B(KEYINPUT105), .ZN(n477) );
  XOR2_X1 U459 ( .A(KEYINPUT7), .B(KEYINPUT106), .Z(n478) );
  INV_X1 U460 ( .A(G134), .ZN(n486) );
  XNOR2_X1 U461 ( .A(G113), .B(G143), .ZN(n492) );
  XOR2_X1 U462 ( .A(G122), .B(G104), .Z(n493) );
  XOR2_X1 U463 ( .A(KEYINPUT102), .B(KEYINPUT100), .Z(n495) );
  XNOR2_X1 U464 ( .A(n596), .B(KEYINPUT39), .ZN(n624) );
  OR2_X1 U465 ( .A1(n639), .A2(G902), .ZN(n534) );
  XNOR2_X1 U466 ( .A(KEYINPUT16), .B(G122), .ZN(n448) );
  NAND2_X1 U467 ( .A1(n411), .A2(n447), .ZN(n444) );
  XNOR2_X1 U468 ( .A(G140), .B(KEYINPUT78), .ZN(n521) );
  NOR2_X1 U469 ( .A1(n755), .A2(G952), .ZN(n688) );
  XNOR2_X1 U470 ( .A(n599), .B(KEYINPUT42), .ZN(n763) );
  XNOR2_X1 U471 ( .A(n435), .B(n434), .ZN(n764) );
  XNOR2_X1 U472 ( .A(KEYINPUT40), .B(KEYINPUT111), .ZN(n434) );
  NAND2_X1 U473 ( .A1(n624), .A2(n742), .ZN(n435) );
  XNOR2_X1 U474 ( .A(n558), .B(n557), .ZN(n396) );
  INV_X1 U475 ( .A(KEYINPUT90), .ZN(n557) );
  INV_X1 U476 ( .A(G122), .ZN(n406) );
  XOR2_X1 U477 ( .A(n540), .B(n539), .Z(n361) );
  XOR2_X1 U478 ( .A(n532), .B(n531), .Z(n362) );
  NOR2_X1 U479 ( .A1(n585), .A2(n598), .ZN(n363) );
  INV_X1 U480 ( .A(n410), .ZN(n699) );
  AND2_X1 U481 ( .A1(n658), .A2(KEYINPUT44), .ZN(n364) );
  NAND2_X1 U482 ( .A1(n568), .A2(n567), .ZN(n365) );
  AND2_X1 U483 ( .A1(n405), .A2(n404), .ZN(n366) );
  AND2_X1 U484 ( .A1(n607), .A2(n433), .ZN(n367) );
  NOR2_X1 U485 ( .A1(n543), .A2(n525), .ZN(n368) );
  INV_X1 U486 ( .A(G902), .ZN(n390) );
  XOR2_X1 U487 ( .A(KEYINPUT91), .B(KEYINPUT33), .Z(n369) );
  INV_X1 U488 ( .A(KEYINPUT1), .ZN(n387) );
  XOR2_X1 U489 ( .A(n639), .B(n638), .Z(n370) );
  XNOR2_X1 U490 ( .A(n523), .B(n383), .ZN(n677) );
  NAND2_X1 U491 ( .A1(n535), .A2(G221), .ZN(n377) );
  INV_X1 U492 ( .A(n647), .ZN(n412) );
  NOR2_X1 U493 ( .A1(n382), .A2(n712), .ZN(n597) );
  XNOR2_X1 U494 ( .A(n383), .B(n362), .ZN(n639) );
  XNOR2_X2 U495 ( .A(n649), .B(G146), .ZN(n383) );
  NAND2_X1 U496 ( .A1(n386), .A2(n384), .ZN(n545) );
  NAND2_X1 U497 ( .A1(n359), .A2(n391), .ZN(n386) );
  NAND2_X1 U498 ( .A1(n391), .A2(n388), .ZN(n584) );
  XNOR2_X1 U499 ( .A(n442), .B(KEYINPUT65), .ZN(n541) );
  INV_X1 U500 ( .A(n424), .ZN(n423) );
  XNOR2_X1 U501 ( .A(n401), .B(n430), .ZN(n411) );
  NAND2_X1 U502 ( .A1(n659), .A2(n390), .ZN(n395) );
  NAND2_X1 U503 ( .A1(n677), .A2(n524), .ZN(n393) );
  OR2_X2 U504 ( .A1(n677), .A2(n389), .ZN(n388) );
  AND2_X1 U505 ( .A1(n394), .A2(n583), .ZN(n706) );
  NAND2_X1 U506 ( .A1(n423), .A2(n422), .ZN(n397) );
  XNOR2_X2 U507 ( .A(n398), .B(n515), .ZN(n556) );
  NAND2_X1 U508 ( .A1(n546), .A2(n514), .ZN(n398) );
  XNOR2_X2 U509 ( .A(n399), .B(n476), .ZN(n546) );
  OR2_X2 U510 ( .A1(n585), .A2(n475), .ZN(n399) );
  NAND2_X1 U511 ( .A1(n556), .A2(n368), .ZN(n544) );
  NAND2_X1 U512 ( .A1(n402), .A2(n412), .ZN(n401) );
  XNOR2_X1 U513 ( .A(n403), .B(KEYINPUT84), .ZN(n402) );
  NOR2_X2 U514 ( .A1(n634), .A2(n627), .ZN(n403) );
  INV_X1 U515 ( .A(n407), .ZN(n404) );
  XNOR2_X1 U516 ( .A(n360), .B(n406), .ZN(G24) );
  XNOR2_X1 U517 ( .A(n407), .B(KEYINPUT68), .ZN(n428) );
  NAND2_X1 U518 ( .A1(n363), .A2(n608), .ZN(n609) );
  NAND2_X1 U519 ( .A1(n363), .A2(n587), .ZN(n607) );
  NAND2_X1 U520 ( .A1(n363), .A2(n744), .ZN(n738) );
  NAND2_X1 U521 ( .A1(n363), .A2(n742), .ZN(n741) );
  NAND2_X1 U522 ( .A1(n418), .A2(n417), .ZN(n416) );
  NAND2_X1 U523 ( .A1(n582), .A2(n583), .ZN(n420) );
  XNOR2_X1 U524 ( .A(n421), .B(n751), .ZN(n462) );
  XNOR2_X2 U525 ( .A(n750), .B(n529), .ZN(n421) );
  XNOR2_X1 U526 ( .A(n421), .B(n522), .ZN(n523) );
  NAND2_X1 U527 ( .A1(n424), .A2(n742), .ZN(n743) );
  NAND2_X1 U528 ( .A1(n424), .A2(n744), .ZN(n745) );
  NOR2_X2 U529 ( .A1(n663), .A2(n688), .ZN(n664) );
  NOR2_X2 U530 ( .A1(n668), .A2(n688), .ZN(n669) );
  NOR2_X2 U531 ( .A1(n689), .A2(n688), .ZN(n691) );
  NOR2_X2 U532 ( .A1(n675), .A2(n688), .ZN(n676) );
  NAND2_X1 U533 ( .A1(n427), .A2(n425), .ZN(n571) );
  NAND2_X1 U534 ( .A1(n428), .A2(KEYINPUT64), .ZN(n427) );
  INV_X1 U535 ( .A(n547), .ZN(n717) );
  XNOR2_X2 U536 ( .A(n701), .B(KEYINPUT6), .ZN(n604) );
  AND2_X1 U537 ( .A1(n583), .A2(n436), .ZN(n589) );
  XNOR2_X2 U538 ( .A(n534), .B(n533), .ZN(n583) );
  XNOR2_X2 U539 ( .A(n441), .B(n440), .ZN(n531) );
  XNOR2_X2 U540 ( .A(KEYINPUT3), .B(G119), .ZN(n440) );
  XNOR2_X2 U541 ( .A(G113), .B(G116), .ZN(n441) );
  NAND2_X1 U542 ( .A1(n556), .A2(n445), .ZN(n442) );
  INV_X1 U543 ( .A(n694), .ZN(n443) );
  XNOR2_X1 U544 ( .A(n574), .B(n573), .ZN(n634) );
  AND2_X1 U545 ( .A1(n525), .A2(n701), .ZN(n445) );
  OR2_X1 U546 ( .A1(n629), .A2(n628), .ZN(n447) );
  XNOR2_X1 U547 ( .A(n640), .B(n370), .ZN(n642) );
  XNOR2_X1 U548 ( .A(n531), .B(n448), .ZN(n751) );
  XNOR2_X2 U549 ( .A(KEYINPUT76), .B(G110), .ZN(n450) );
  XNOR2_X2 U550 ( .A(n451), .B(n450), .ZN(n750) );
  XNOR2_X1 U551 ( .A(n453), .B(n452), .ZN(n456) );
  NAND2_X1 U552 ( .A1(n755), .A2(G224), .ZN(n454) );
  XNOR2_X1 U553 ( .A(n454), .B(KEYINPUT93), .ZN(n455) );
  XNOR2_X1 U554 ( .A(n456), .B(n455), .ZN(n460) );
  XNOR2_X2 U555 ( .A(G143), .B(G128), .ZN(n487) );
  XNOR2_X1 U556 ( .A(n457), .B(G146), .ZN(n503) );
  INV_X1 U557 ( .A(n503), .ZN(n458) );
  XNOR2_X1 U558 ( .A(n487), .B(n458), .ZN(n459) );
  XNOR2_X1 U559 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U560 ( .A(n462), .B(n461), .ZN(n685) );
  XNOR2_X2 U561 ( .A(KEYINPUT15), .B(G902), .ZN(n627) );
  NAND2_X1 U562 ( .A1(n685), .A2(n627), .ZN(n467) );
  NAND2_X1 U563 ( .A1(n390), .A2(n463), .ZN(n468) );
  NAND2_X1 U564 ( .A1(n468), .A2(G210), .ZN(n465) );
  INV_X1 U565 ( .A(KEYINPUT95), .ZN(n464) );
  XNOR2_X1 U566 ( .A(n465), .B(n464), .ZN(n466) );
  AND2_X1 U567 ( .A1(n468), .A2(G214), .ZN(n709) );
  XNOR2_X1 U568 ( .A(n469), .B(KEYINPUT19), .ZN(n585) );
  XNOR2_X1 U569 ( .A(n470), .B(KEYINPUT14), .ZN(n472) );
  NAND2_X1 U570 ( .A1(G952), .A2(n472), .ZN(n471) );
  XOR2_X1 U571 ( .A(KEYINPUT96), .B(n471), .Z(n723) );
  AND2_X1 U572 ( .A1(n723), .A2(n755), .ZN(n578) );
  NAND2_X1 U573 ( .A1(G902), .A2(n472), .ZN(n575) );
  INV_X1 U574 ( .A(G898), .ZN(n473) );
  NAND2_X1 U575 ( .A1(n473), .A2(G953), .ZN(n753) );
  NOR2_X1 U576 ( .A1(n575), .A2(n753), .ZN(n474) );
  NOR2_X1 U577 ( .A1(n578), .A2(n474), .ZN(n475) );
  INV_X1 U578 ( .A(KEYINPUT0), .ZN(n476) );
  XNOR2_X1 U579 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U580 ( .A(n479), .B(G116), .ZN(n484) );
  NAND2_X1 U581 ( .A1(n755), .A2(G234), .ZN(n481) );
  INV_X1 U582 ( .A(KEYINPUT70), .ZN(n480) );
  XOR2_X1 U583 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n482) );
  NAND2_X1 U584 ( .A1(n535), .A2(G217), .ZN(n483) );
  XNOR2_X1 U585 ( .A(n484), .B(n483), .ZN(n490) );
  XNOR2_X1 U586 ( .A(KEYINPUT9), .B(n485), .ZN(n488) );
  XNOR2_X2 U587 ( .A(n487), .B(n486), .ZN(n519) );
  XNOR2_X1 U588 ( .A(n519), .B(n488), .ZN(n489) );
  XNOR2_X1 U589 ( .A(n490), .B(n489), .ZN(n665) );
  NAND2_X1 U590 ( .A1(n665), .A2(n390), .ZN(n491) );
  XNOR2_X1 U591 ( .A(n491), .B(G478), .ZN(n613) );
  XNOR2_X1 U592 ( .A(n493), .B(n492), .ZN(n497) );
  XNOR2_X1 U593 ( .A(G131), .B(KEYINPUT11), .ZN(n494) );
  XNOR2_X1 U594 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U595 ( .A(n497), .B(n496), .ZN(n501) );
  XOR2_X1 U596 ( .A(KEYINPUT101), .B(KEYINPUT12), .Z(n499) );
  NAND2_X1 U597 ( .A1(G214), .A2(n526), .ZN(n498) );
  XNOR2_X1 U598 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U599 ( .A(n501), .B(n500), .ZN(n505) );
  XNOR2_X1 U600 ( .A(G140), .B(KEYINPUT10), .ZN(n502) );
  XNOR2_X1 U601 ( .A(n502), .B(KEYINPUT71), .ZN(n504) );
  XNOR2_X1 U602 ( .A(n504), .B(n503), .ZN(n648) );
  XNOR2_X1 U603 ( .A(n505), .B(n648), .ZN(n672) );
  NAND2_X1 U604 ( .A1(n672), .A2(n390), .ZN(n509) );
  XOR2_X1 U605 ( .A(KEYINPUT104), .B(KEYINPUT13), .Z(n507) );
  XNOR2_X1 U606 ( .A(KEYINPUT103), .B(G475), .ZN(n506) );
  XOR2_X1 U607 ( .A(n507), .B(n506), .Z(n508) );
  XNOR2_X1 U608 ( .A(n509), .B(n508), .ZN(n563) );
  OR2_X1 U609 ( .A1(n613), .A2(n563), .ZN(n712) );
  NAND2_X1 U610 ( .A1(n627), .A2(G234), .ZN(n510) );
  XNOR2_X1 U611 ( .A(n510), .B(KEYINPUT20), .ZN(n538) );
  INV_X1 U612 ( .A(n538), .ZN(n512) );
  INV_X1 U613 ( .A(G221), .ZN(n511) );
  OR2_X1 U614 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U615 ( .A(n513), .B(KEYINPUT21), .ZN(n698) );
  NOR2_X1 U616 ( .A1(n712), .A2(n698), .ZN(n514) );
  XNOR2_X1 U617 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n515) );
  XNOR2_X1 U618 ( .A(KEYINPUT4), .B(G131), .ZN(n517) );
  XNOR2_X1 U619 ( .A(G137), .B(KEYINPUT72), .ZN(n516) );
  XNOR2_X1 U620 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X2 U621 ( .A(n519), .B(n518), .ZN(n649) );
  NAND2_X1 U622 ( .A1(n755), .A2(G227), .ZN(n520) );
  XNOR2_X1 U623 ( .A(n521), .B(n520), .ZN(n522) );
  INV_X1 U624 ( .A(G469), .ZN(n524) );
  NAND2_X1 U625 ( .A1(n526), .A2(G210), .ZN(n528) );
  XNOR2_X1 U626 ( .A(n528), .B(n527), .ZN(n530) );
  XNOR2_X1 U627 ( .A(n530), .B(n529), .ZN(n532) );
  XNOR2_X1 U628 ( .A(KEYINPUT98), .B(G472), .ZN(n533) );
  INV_X1 U629 ( .A(n648), .ZN(n536) );
  AND2_X1 U630 ( .A1(n538), .A2(G217), .ZN(n540) );
  XNOR2_X1 U631 ( .A(KEYINPUT77), .B(KEYINPUT25), .ZN(n539) );
  INV_X1 U632 ( .A(n699), .ZN(n542) );
  NAND2_X2 U633 ( .A1(n541), .A2(n699), .ZN(n646) );
  OR2_X1 U634 ( .A1(n604), .A2(n542), .ZN(n543) );
  NAND2_X1 U635 ( .A1(n547), .A2(n562), .ZN(n549) );
  INV_X1 U636 ( .A(KEYINPUT34), .ZN(n548) );
  XNOR2_X1 U637 ( .A(n549), .B(n548), .ZN(n551) );
  AND2_X1 U638 ( .A1(n613), .A2(n563), .ZN(n550) );
  NAND2_X1 U639 ( .A1(n551), .A2(n550), .ZN(n553) );
  XNOR2_X1 U640 ( .A(KEYINPUT88), .B(KEYINPUT35), .ZN(n552) );
  INV_X1 U641 ( .A(n604), .ZN(n554) );
  AND2_X1 U642 ( .A1(n554), .A2(n525), .ZN(n555) );
  NAND2_X1 U643 ( .A1(n556), .A2(n555), .ZN(n558) );
  NAND2_X1 U644 ( .A1(n706), .A2(n562), .ZN(n560) );
  XOR2_X1 U645 ( .A(KEYINPUT99), .B(KEYINPUT31), .Z(n559) );
  OR2_X1 U646 ( .A1(n584), .A2(n696), .ZN(n590) );
  NOR2_X1 U647 ( .A1(n590), .A2(n583), .ZN(n561) );
  AND2_X1 U648 ( .A1(n562), .A2(n561), .ZN(n733) );
  INV_X1 U649 ( .A(n563), .ZN(n612) );
  INV_X1 U650 ( .A(n613), .ZN(n564) );
  NOR2_X1 U651 ( .A1(n564), .A2(n563), .ZN(n744) );
  NOR2_X1 U652 ( .A1(n742), .A2(n744), .ZN(n713) );
  INV_X1 U653 ( .A(n713), .ZN(n608) );
  NAND2_X1 U654 ( .A1(n446), .A2(n366), .ZN(n569) );
  AND2_X1 U655 ( .A1(n657), .A2(n565), .ZN(n568) );
  INV_X1 U656 ( .A(KEYINPUT44), .ZN(n566) );
  AND2_X1 U657 ( .A1(n566), .A2(KEYINPUT64), .ZN(n567) );
  NAND2_X1 U658 ( .A1(n569), .A2(n365), .ZN(n572) );
  AND2_X1 U659 ( .A1(n646), .A2(n658), .ZN(n570) );
  NAND2_X1 U660 ( .A1(n572), .A2(n571), .ZN(n574) );
  XNOR2_X1 U661 ( .A(KEYINPUT87), .B(KEYINPUT45), .ZN(n573) );
  NOR2_X1 U662 ( .A1(G900), .A2(n575), .ZN(n576) );
  AND2_X1 U663 ( .A1(n576), .A2(G953), .ZN(n577) );
  NOR2_X1 U664 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U665 ( .A(n579), .B(KEYINPUT79), .ZN(n594) );
  INV_X1 U666 ( .A(n698), .ZN(n580) );
  AND2_X1 U667 ( .A1(n594), .A2(n580), .ZN(n581) );
  NAND2_X1 U668 ( .A1(n699), .A2(n581), .ZN(n601) );
  INV_X1 U669 ( .A(n601), .ZN(n582) );
  NOR2_X1 U670 ( .A1(n713), .A2(KEYINPUT47), .ZN(n586) );
  XNOR2_X1 U671 ( .A(KEYINPUT74), .B(n586), .ZN(n587) );
  XNOR2_X1 U672 ( .A(KEYINPUT30), .B(KEYINPUT109), .ZN(n588) );
  XNOR2_X1 U673 ( .A(n589), .B(n588), .ZN(n591) );
  NOR2_X1 U674 ( .A1(n591), .A2(n590), .ZN(n610) );
  INV_X1 U675 ( .A(KEYINPUT38), .ZN(n593) );
  BUF_X1 U676 ( .A(n592), .Z(n622) );
  XNOR2_X1 U677 ( .A(n593), .B(n622), .ZN(n710) );
  INV_X1 U678 ( .A(n594), .ZN(n611) );
  NOR2_X1 U679 ( .A1(n710), .A2(n611), .ZN(n595) );
  NAND2_X1 U680 ( .A1(n610), .A2(n595), .ZN(n596) );
  INV_X1 U681 ( .A(n764), .ZN(n600) );
  XNOR2_X1 U682 ( .A(n597), .B(KEYINPUT41), .ZN(n726) );
  NOR2_X1 U683 ( .A1(n601), .A2(n709), .ZN(n602) );
  AND2_X1 U684 ( .A1(n742), .A2(n602), .ZN(n603) );
  NAND2_X1 U685 ( .A1(n604), .A2(n603), .ZN(n619) );
  NOR2_X1 U686 ( .A1(n619), .A2(n622), .ZN(n605) );
  XOR2_X1 U687 ( .A(KEYINPUT36), .B(n605), .Z(n606) );
  NOR2_X1 U688 ( .A1(n606), .A2(n525), .ZN(n746) );
  NAND2_X1 U689 ( .A1(n609), .A2(KEYINPUT47), .ZN(n617) );
  NOR2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n614) );
  NAND2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U692 ( .A1(n615), .A2(n622), .ZN(n616) );
  NAND2_X1 U693 ( .A1(n610), .A2(n616), .ZN(n644) );
  NAND2_X1 U694 ( .A1(n617), .A2(n644), .ZN(n618) );
  XOR2_X1 U695 ( .A(n619), .B(KEYINPUT108), .Z(n620) );
  NAND2_X1 U696 ( .A1(n620), .A2(n525), .ZN(n621) );
  XNOR2_X1 U697 ( .A(n621), .B(KEYINPUT43), .ZN(n623) );
  NAND2_X1 U698 ( .A1(n623), .A2(n622), .ZN(n645) );
  NAND2_X1 U699 ( .A1(n624), .A2(n744), .ZN(n625) );
  XNOR2_X1 U700 ( .A(n625), .B(KEYINPUT112), .ZN(n765) );
  AND2_X1 U701 ( .A1(n645), .A2(n765), .ZN(n626) );
  XNOR2_X1 U702 ( .A(n627), .B(KEYINPUT86), .ZN(n629) );
  INV_X1 U703 ( .A(KEYINPUT2), .ZN(n628) );
  NAND2_X1 U704 ( .A1(n765), .A2(KEYINPUT2), .ZN(n630) );
  XOR2_X1 U705 ( .A(KEYINPUT80), .B(n630), .Z(n631) );
  AND2_X1 U706 ( .A1(n631), .A2(n645), .ZN(n632) );
  NAND2_X1 U707 ( .A1(n633), .A2(n632), .ZN(n636) );
  BUF_X1 U708 ( .A(n634), .Z(n635) );
  NOR2_X1 U709 ( .A1(n636), .A2(n635), .ZN(n694) );
  NAND2_X1 U710 ( .A1(n683), .A2(G472), .ZN(n640) );
  XOR2_X1 U711 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n637) );
  XNOR2_X1 U712 ( .A(n637), .B(KEYINPUT62), .ZN(n638) );
  INV_X1 U713 ( .A(n688), .ZN(n641) );
  NAND2_X1 U714 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U715 ( .A(n643), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U716 ( .A(n644), .B(G143), .ZN(G45) );
  XNOR2_X1 U717 ( .A(n645), .B(G140), .ZN(G42) );
  XNOR2_X1 U718 ( .A(n646), .B(G110), .ZN(G12) );
  XNOR2_X1 U719 ( .A(n649), .B(n648), .ZN(n651) );
  XNOR2_X1 U720 ( .A(n647), .B(n651), .ZN(n650) );
  NAND2_X1 U721 ( .A1(n650), .A2(n755), .ZN(n655) );
  XNOR2_X1 U722 ( .A(n651), .B(G227), .ZN(n652) );
  NAND2_X1 U723 ( .A1(G900), .A2(n652), .ZN(n653) );
  NAND2_X1 U724 ( .A1(n653), .A2(G953), .ZN(n654) );
  NAND2_X1 U725 ( .A1(n655), .A2(n654), .ZN(G72) );
  XOR2_X1 U726 ( .A(G101), .B(KEYINPUT115), .Z(n656) );
  XNOR2_X1 U727 ( .A(n657), .B(n656), .ZN(G3) );
  XNOR2_X1 U728 ( .A(n658), .B(G119), .ZN(G21) );
  NAND2_X1 U729 ( .A1(n683), .A2(G217), .ZN(n662) );
  BUF_X1 U730 ( .A(n659), .Z(n660) );
  XNOR2_X1 U731 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U732 ( .A(n664), .B(KEYINPUT126), .ZN(G66) );
  NAND2_X1 U733 ( .A1(n683), .A2(G478), .ZN(n667) );
  XNOR2_X1 U734 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U735 ( .A(n669), .B(KEYINPUT124), .ZN(G63) );
  NAND2_X1 U736 ( .A1(n683), .A2(G475), .ZN(n674) );
  XNOR2_X1 U737 ( .A(KEYINPUT66), .B(KEYINPUT92), .ZN(n670) );
  XNOR2_X1 U738 ( .A(n670), .B(KEYINPUT59), .ZN(n671) );
  XNOR2_X1 U739 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U740 ( .A(n676), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U741 ( .A1(n683), .A2(G469), .ZN(n681) );
  XOR2_X1 U742 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n678) );
  XNOR2_X1 U743 ( .A(n678), .B(KEYINPUT58), .ZN(n679) );
  XNOR2_X1 U744 ( .A(n677), .B(n679), .ZN(n680) );
  XNOR2_X1 U745 ( .A(n681), .B(n680), .ZN(n682) );
  NOR2_X1 U746 ( .A1(n682), .A2(n688), .ZN(G54) );
  NAND2_X1 U747 ( .A1(n683), .A2(G210), .ZN(n687) );
  XNOR2_X1 U748 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n684) );
  XNOR2_X1 U749 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X1 U750 ( .A(n687), .B(n686), .ZN(n689) );
  XOR2_X1 U751 ( .A(KEYINPUT89), .B(KEYINPUT56), .Z(n690) );
  XNOR2_X1 U752 ( .A(n691), .B(n690), .ZN(G51) );
  NOR2_X1 U753 ( .A1(n647), .A2(n635), .ZN(n692) );
  NOR2_X1 U754 ( .A1(n692), .A2(KEYINPUT2), .ZN(n693) );
  NOR2_X1 U755 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U756 ( .A(KEYINPUT85), .B(n695), .Z(n730) );
  NAND2_X1 U757 ( .A1(n525), .A2(n696), .ZN(n697) );
  XOR2_X1 U758 ( .A(KEYINPUT50), .B(n697), .Z(n704) );
  NAND2_X1 U759 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U760 ( .A(KEYINPUT49), .B(n700), .Z(n702) );
  NAND2_X1 U761 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U762 ( .A1(n704), .A2(n703), .ZN(n705) );
  OR2_X1 U763 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U764 ( .A(KEYINPUT51), .B(n707), .ZN(n708) );
  NOR2_X1 U765 ( .A1(n726), .A2(n708), .ZN(n720) );
  AND2_X1 U766 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U767 ( .A1(n712), .A2(n711), .ZN(n715) );
  NOR2_X1 U768 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U769 ( .A(n716), .B(KEYINPUT120), .ZN(n718) );
  NOR2_X1 U770 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U771 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U772 ( .A(n721), .B(KEYINPUT121), .ZN(n722) );
  XNOR2_X1 U773 ( .A(n722), .B(KEYINPUT52), .ZN(n724) );
  NAND2_X1 U774 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U775 ( .A1(n725), .A2(n755), .ZN(n728) );
  NOR2_X1 U776 ( .A1(n726), .A2(n717), .ZN(n727) );
  OR2_X1 U777 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U778 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U779 ( .A(n731), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U780 ( .A1(n733), .A2(n742), .ZN(n732) );
  XNOR2_X1 U781 ( .A(n732), .B(G104), .ZN(G6) );
  XNOR2_X1 U782 ( .A(n357), .B(KEYINPUT27), .ZN(n737) );
  XOR2_X1 U783 ( .A(KEYINPUT116), .B(KEYINPUT26), .Z(n735) );
  NAND2_X1 U784 ( .A1(n733), .A2(n744), .ZN(n734) );
  XNOR2_X1 U785 ( .A(n735), .B(n734), .ZN(n736) );
  XNOR2_X1 U786 ( .A(n737), .B(n736), .ZN(G9) );
  XOR2_X1 U787 ( .A(KEYINPUT117), .B(KEYINPUT29), .Z(n739) );
  XNOR2_X1 U788 ( .A(n739), .B(n738), .ZN(n740) );
  XOR2_X1 U789 ( .A(G128), .B(n740), .Z(G30) );
  XNOR2_X1 U790 ( .A(n741), .B(G146), .ZN(G48) );
  XNOR2_X1 U791 ( .A(n743), .B(G113), .ZN(G15) );
  XNOR2_X1 U792 ( .A(n745), .B(G116), .ZN(G18) );
  XNOR2_X1 U793 ( .A(n746), .B(KEYINPUT118), .ZN(n747) );
  XNOR2_X1 U794 ( .A(n747), .B(KEYINPUT37), .ZN(n748) );
  XNOR2_X1 U795 ( .A(G125), .B(n748), .ZN(G27) );
  XOR2_X1 U796 ( .A(G101), .B(KEYINPUT127), .Z(n749) );
  XNOR2_X1 U797 ( .A(n750), .B(n749), .ZN(n752) );
  XNOR2_X1 U798 ( .A(n752), .B(n751), .ZN(n754) );
  AND2_X1 U799 ( .A1(n754), .A2(n753), .ZN(n762) );
  INV_X1 U800 ( .A(n635), .ZN(n756) );
  NAND2_X1 U801 ( .A1(n756), .A2(n755), .ZN(n760) );
  NAND2_X1 U802 ( .A1(G953), .A2(G224), .ZN(n757) );
  XNOR2_X1 U803 ( .A(KEYINPUT61), .B(n757), .ZN(n758) );
  NAND2_X1 U804 ( .A1(n758), .A2(G898), .ZN(n759) );
  NAND2_X1 U805 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U806 ( .A(n762), .B(n761), .ZN(G69) );
  XOR2_X1 U807 ( .A(G137), .B(n763), .Z(G39) );
  XOR2_X1 U808 ( .A(G131), .B(n764), .Z(G33) );
  XOR2_X1 U809 ( .A(G134), .B(n765), .Z(n766) );
  XNOR2_X1 U810 ( .A(KEYINPUT119), .B(n766), .ZN(G36) );
endmodule

