//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 0 1 1 0 1 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1270, new_n1271, new_n1272, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1331, new_n1332, new_n1333;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(KEYINPUT64), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n201), .B(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT65), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n210), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  OR2_X1    g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  NOR2_X1   g0021(.A1(G58), .A2(G68), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n222), .A2(KEYINPUT66), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(KEYINPUT66), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n223), .A2(G50), .A3(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n227), .A2(new_n208), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n213), .A2(new_n221), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n220), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G68), .ZN(new_n245));
  INV_X1    g0045(.A(G68), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n243), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(KEYINPUT74), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT10), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n203), .A2(G20), .ZN(new_n254));
  INV_X1    g0054(.A(G150), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n208), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT8), .B(G58), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT69), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT69), .ZN(new_n260));
  INV_X1    g0060(.A(G58), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT8), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n208), .A2(G33), .ZN(new_n264));
  OAI221_X1 g0064(.A(new_n254), .B1(new_n255), .B2(new_n257), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n227), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(G50), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n267), .B1(new_n207), .B2(G20), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n270), .B1(new_n271), .B2(G50), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT9), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n275), .B(KEYINPUT73), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n268), .A2(new_n272), .ZN(new_n277));
  AOI22_X1  g0077(.A1(new_n277), .A2(KEYINPUT9), .B1(KEYINPUT74), .B2(KEYINPUT10), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT68), .ZN(new_n279));
  AND2_X1   g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n279), .B1(new_n280), .B2(new_n227), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n282), .A2(KEYINPUT68), .A3(G1), .A4(G13), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT3), .B(G33), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G223), .A3(G1698), .ZN(new_n286));
  INV_X1    g0086(.A(G77), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G222), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n286), .B1(new_n287), .B2(new_n285), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT67), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n284), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n293), .B1(new_n292), .B2(new_n291), .ZN(new_n294));
  INV_X1    g0094(.A(G41), .ZN(new_n295));
  INV_X1    g0095(.A(G45), .ZN(new_n296));
  AOI21_X1  g0096(.A(G1), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n282), .A2(G1), .A3(G13), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n297), .A2(new_n298), .A3(G274), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n280), .A2(new_n227), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(new_n297), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n299), .B1(G226), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n294), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G190), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(G200), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n278), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n252), .B(new_n253), .C1(new_n276), .C2(new_n307), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n278), .A2(new_n306), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT73), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n275), .B(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n252), .A2(new_n253), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n309), .A2(new_n311), .A3(new_n312), .A4(new_n305), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n263), .A2(new_n271), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n269), .B2(new_n263), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT16), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT3), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G33), .ZN(new_n321));
  AOI21_X1  g0121(.A(G20), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT77), .B1(new_n322), .B2(KEYINPUT7), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT77), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT7), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n324), .B(new_n325), .C1(new_n285), .C2(G20), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n319), .A2(new_n321), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n328), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT78), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n322), .A2(KEYINPUT78), .A3(KEYINPUT7), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n246), .B1(new_n327), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n261), .A2(new_n246), .ZN(new_n335));
  OAI21_X1  g0135(.A(G20), .B1(new_n335), .B2(new_n222), .ZN(new_n336));
  INV_X1    g0136(.A(G159), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n336), .B1(new_n337), .B2(new_n257), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n318), .B1(new_n334), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n267), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n325), .B1(new_n285), .B2(G20), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n329), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n338), .B1(new_n342), .B2(G68), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n340), .B1(new_n343), .B2(KEYINPUT16), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n317), .B1(new_n339), .B2(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n319), .A2(new_n321), .A3(G223), .A4(new_n288), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n319), .A2(new_n321), .A3(G226), .A4(G1698), .ZN(new_n347));
  NAND2_X1  g0147(.A1(G33), .A2(G87), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT79), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT79), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n346), .A2(new_n347), .A3(new_n351), .A4(new_n348), .ZN(new_n352));
  AND2_X1   g0152(.A1(new_n281), .A2(new_n283), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n350), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n299), .B1(G232), .B2(new_n301), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G169), .ZN(new_n357));
  XNOR2_X1  g0157(.A(KEYINPUT70), .B(G179), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n354), .A2(new_n359), .A3(new_n355), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT18), .B1(new_n345), .B2(new_n361), .ZN(new_n362));
  NOR4_X1   g0162(.A1(new_n285), .A2(new_n330), .A3(new_n325), .A4(G20), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT78), .B1(new_n322), .B2(KEYINPUT7), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n323), .B(new_n326), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n338), .B1(new_n365), .B2(G68), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n344), .B1(new_n366), .B2(KEYINPUT16), .ZN(new_n367));
  INV_X1    g0167(.A(new_n317), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT18), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n357), .A2(new_n360), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n362), .A2(new_n372), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n354), .A2(G190), .A3(new_n355), .ZN(new_n374));
  INV_X1    g0174(.A(G200), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n375), .B1(new_n354), .B2(new_n355), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n377), .A2(new_n367), .A3(new_n368), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT17), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n345), .A2(KEYINPUT17), .A3(new_n377), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n373), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n273), .B1(new_n304), .B2(G169), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n303), .A2(new_n359), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n269), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n287), .ZN(new_n388));
  INV_X1    g0188(.A(new_n271), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n388), .B1(new_n389), .B2(new_n287), .ZN(new_n390));
  OAI22_X1  g0190(.A1(new_n258), .A2(new_n257), .B1(new_n208), .B2(new_n287), .ZN(new_n391));
  XNOR2_X1  g0191(.A(KEYINPUT15), .B(G87), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n392), .A2(new_n264), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n267), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT71), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g0196(.A(KEYINPUT71), .B(new_n267), .C1(new_n391), .C2(new_n393), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n390), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n285), .A2(G232), .A3(new_n288), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n285), .A2(G238), .A3(G1698), .ZN(new_n400));
  INV_X1    g0200(.A(G107), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n399), .B(new_n400), .C1(new_n401), .C2(new_n285), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n353), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n299), .B1(G244), .B2(new_n301), .ZN(new_n404));
  AOI21_X1  g0204(.A(G169), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n398), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT72), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT72), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n398), .B2(new_n405), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n403), .A2(new_n404), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n358), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n407), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n410), .A2(G190), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n403), .A2(new_n404), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(G200), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n414), .A2(new_n398), .A3(new_n416), .ZN(new_n417));
  NOR3_X1   g0217(.A1(new_n386), .A2(new_n413), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n387), .A2(KEYINPUT12), .A3(new_n246), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT12), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n269), .B2(G68), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n419), .B(new_n421), .C1(new_n389), .C2(new_n246), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n422), .A2(KEYINPUT75), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(KEYINPUT75), .ZN(new_n424));
  OAI22_X1  g0224(.A1(new_n257), .A2(new_n244), .B1(new_n208), .B2(G68), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n264), .A2(new_n287), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n267), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n427), .B(KEYINPUT11), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n423), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G33), .A2(G97), .ZN(new_n430));
  INV_X1    g0230(.A(G226), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n430), .B1(new_n289), .B2(new_n431), .ZN(new_n432));
  NOR3_X1   g0232(.A1(new_n328), .A2(new_n233), .A3(new_n288), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n353), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n299), .B1(G238), .B2(new_n301), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT13), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT13), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n434), .A2(new_n438), .A3(new_n435), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(G179), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(KEYINPUT76), .A2(G169), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n441), .B1(new_n437), .B2(new_n439), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT14), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n440), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n441), .ZN(new_n445));
  INV_X1    g0245(.A(new_n439), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n438), .B1(new_n434), .B2(new_n435), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n443), .B(new_n445), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n429), .B1(new_n444), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n446), .A2(new_n447), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n429), .B1(new_n451), .B2(G190), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n375), .B2(new_n451), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n315), .A2(new_n383), .A3(new_n418), .A4(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n296), .A2(G1), .ZN(new_n458));
  XNOR2_X1  g0258(.A(KEYINPUT5), .B(G41), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n300), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n459), .A2(new_n458), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n298), .A2(G274), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n460), .A2(G257), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT80), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n319), .A2(new_n321), .A3(G244), .A4(new_n288), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT4), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G283), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G250), .A2(G1698), .ZN(new_n470));
  NAND2_X1  g0270(.A1(KEYINPUT4), .A2(G244), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n470), .B1(new_n471), .B2(G1698), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n469), .B1(new_n285), .B2(new_n472), .ZN(new_n473));
  AOI211_X1 g0273(.A(new_n464), .B(new_n284), .C1(new_n467), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n467), .A2(new_n473), .ZN(new_n475));
  AOI21_X1  g0275(.A(KEYINPUT80), .B1(new_n475), .B2(new_n353), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n463), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G200), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT81), .ZN(new_n479));
  INV_X1    g0279(.A(G97), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n387), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n207), .A2(G33), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n269), .A2(new_n482), .A3(new_n227), .A4(new_n266), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n481), .B1(new_n483), .B2(new_n480), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n365), .A2(G107), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT6), .ZN(new_n486));
  NOR3_X1   g0286(.A1(new_n486), .A2(new_n480), .A3(G107), .ZN(new_n487));
  XNOR2_X1  g0287(.A(G97), .B(G107), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n487), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  OAI22_X1  g0289(.A1(new_n489), .A2(new_n208), .B1(new_n287), .B2(new_n257), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n485), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n484), .B1(new_n492), .B2(new_n267), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT81), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n477), .A2(new_n494), .A3(G200), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n475), .A2(new_n353), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n496), .A2(new_n463), .A3(G190), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n479), .A2(new_n493), .A3(new_n495), .A4(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n392), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n499), .A2(new_n269), .ZN(new_n500));
  NOR2_X1   g0300(.A1(G97), .A2(G107), .ZN(new_n501));
  INV_X1    g0301(.A(G87), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n501), .A2(new_n502), .B1(new_n430), .B2(new_n208), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT19), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G97), .ZN(new_n505));
  OAI22_X1  g0305(.A1(new_n503), .A2(new_n504), .B1(new_n264), .B2(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n285), .A2(KEYINPUT82), .A3(new_n208), .A4(G68), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n319), .A2(new_n321), .A3(new_n208), .A4(G68), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT82), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n506), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n500), .B1(new_n511), .B2(new_n267), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n298), .A2(G274), .A3(new_n458), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n207), .A2(G45), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n514), .B(G250), .C1(new_n280), .C2(new_n227), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n319), .A2(new_n321), .A3(G244), .A4(G1698), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n319), .A2(new_n321), .A3(G238), .A4(new_n288), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G116), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n516), .B1(new_n520), .B2(new_n353), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G190), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n483), .A2(new_n502), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n512), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n520), .A2(new_n353), .ZN(new_n526));
  INV_X1    g0326(.A(new_n516), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G200), .ZN(new_n529));
  AOI211_X1 g0329(.A(new_n359), .B(new_n516), .C1(new_n353), .C2(new_n520), .ZN(new_n530));
  AOI21_X1  g0330(.A(G169), .B1(new_n526), .B2(new_n527), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n483), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n499), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n512), .A2(new_n534), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n525), .A2(new_n529), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n358), .B(new_n463), .C1(new_n474), .C2(new_n476), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n496), .A2(new_n463), .ZN(new_n538));
  INV_X1    g0338(.A(G169), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n484), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n490), .B1(new_n365), .B2(G107), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n543), .B1(new_n544), .B2(new_n340), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n498), .A2(new_n536), .A3(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT83), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n498), .A2(KEYINPUT83), .A3(new_n536), .A4(new_n546), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n319), .A2(new_n321), .A3(new_n208), .A4(G87), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT22), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT22), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n285), .A2(new_n554), .A3(new_n208), .A4(G87), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT24), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT23), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n208), .B2(G107), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n401), .A2(KEYINPUT23), .A3(G20), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT86), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n519), .B2(G20), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n208), .A2(KEYINPUT86), .A3(G33), .A4(G116), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n561), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n556), .A2(new_n557), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n557), .B1(new_n556), .B2(new_n565), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n267), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n387), .A2(KEYINPUT25), .A3(new_n401), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT25), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(new_n269), .B2(G107), .ZN(new_n571));
  AOI22_X1  g0371(.A1(G107), .A2(new_n533), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n319), .A2(new_n321), .A3(G257), .A4(G1698), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n319), .A2(new_n321), .A3(G250), .A4(new_n288), .ZN(new_n575));
  NAND2_X1  g0375(.A1(G33), .A2(G294), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n353), .A2(new_n577), .B1(new_n460), .B2(G264), .ZN(new_n578));
  INV_X1    g0378(.A(G179), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n461), .A2(new_n462), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n578), .A2(new_n580), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n539), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n573), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(G190), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n577), .A2(new_n353), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n460), .A2(G264), .ZN(new_n587));
  AND4_X1   g0387(.A1(new_n585), .A2(new_n586), .A3(new_n580), .A4(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(G200), .B1(new_n578), .B2(new_n580), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n568), .B(new_n572), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n533), .A2(KEYINPUT84), .A3(G116), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT84), .ZN(new_n594));
  INV_X1    g0394(.A(G116), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n594), .B1(new_n483), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n387), .A2(new_n595), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n266), .A2(new_n227), .B1(G20), .B2(new_n595), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n468), .B(new_n208), .C1(G33), .C2(new_n480), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT20), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n599), .A2(KEYINPUT20), .A3(new_n600), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n597), .A2(new_n598), .A3(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n285), .A2(G264), .A3(G1698), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n285), .A2(G257), .A3(new_n288), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n328), .A2(G303), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n353), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n460), .A2(G270), .B1(new_n461), .B2(new_n462), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(G200), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT85), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n607), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n375), .B1(new_n612), .B2(new_n613), .ZN(new_n618));
  OAI21_X1  g0418(.A(KEYINPUT85), .B1(new_n618), .B2(new_n606), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n612), .A2(new_n613), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G190), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n617), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n539), .B1(new_n612), .B2(new_n613), .ZN(new_n623));
  AOI21_X1  g0423(.A(KEYINPUT21), .B1(new_n623), .B2(new_n606), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n620), .A2(new_n606), .A3(G179), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n623), .A2(new_n606), .A3(KEYINPUT21), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n622), .A2(new_n628), .ZN(new_n629));
  AND4_X1   g0429(.A1(new_n457), .A2(new_n551), .A3(new_n592), .A4(new_n629), .ZN(G372));
  INV_X1    g0430(.A(KEYINPUT90), .ZN(new_n631));
  NOR3_X1   g0431(.A1(new_n345), .A2(new_n361), .A3(KEYINPUT18), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n370), .B1(new_n369), .B2(new_n371), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n362), .A2(KEYINPUT90), .A3(new_n372), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n450), .A2(new_n412), .ZN(new_n637));
  INV_X1    g0437(.A(new_n382), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(new_n638), .A3(new_n453), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n314), .B1(new_n636), .B2(new_n639), .ZN(new_n640));
  OR3_X1    g0440(.A1(new_n640), .A2(KEYINPUT91), .A3(new_n386), .ZN(new_n641));
  OAI21_X1  g0441(.A(KEYINPUT91), .B1(new_n640), .B2(new_n386), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT87), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n644), .B1(new_n528), .B2(G200), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n521), .A2(KEYINPUT87), .A3(new_n375), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n647), .A2(new_n525), .B1(new_n535), .B2(new_n532), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT88), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n541), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n537), .A2(KEYINPUT88), .A3(new_n540), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n648), .A2(new_n650), .A3(new_n545), .A4(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT26), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n536), .A2(new_n542), .A3(KEYINPUT26), .A4(new_n545), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT89), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n493), .A2(new_n541), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n658), .A2(KEYINPUT89), .A3(KEYINPUT26), .A4(new_n536), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n654), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n532), .A2(new_n535), .ZN(new_n661));
  INV_X1    g0461(.A(new_n584), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n590), .B(new_n648), .C1(new_n662), .C2(new_n628), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n498), .A2(new_n546), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n661), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n643), .B1(new_n456), .B2(new_n666), .ZN(G369));
  OR2_X1    g0467(.A1(new_n629), .A2(KEYINPUT92), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n629), .A2(KEYINPUT92), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n668), .B(new_n669), .C1(new_n607), .C2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n627), .A2(new_n626), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(new_n624), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n679), .A2(new_n606), .A3(new_n675), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G330), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n676), .B1(new_n568), .B2(new_n572), .ZN(new_n684));
  OAI22_X1  g0484(.A1(new_n591), .A2(new_n684), .B1(new_n584), .B2(new_n676), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n628), .A2(new_n676), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(new_n591), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n688), .B1(new_n662), .B2(new_n676), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n686), .A2(new_n689), .ZN(G399));
  INV_X1    g0490(.A(new_n211), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(G41), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n501), .A2(new_n502), .A3(new_n595), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n692), .A2(new_n693), .A3(new_n207), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(new_n226), .B2(new_n692), .ZN(new_n695));
  XOR2_X1   g0495(.A(new_n695), .B(KEYINPUT28), .Z(new_n696));
  INV_X1    g0496(.A(KEYINPUT94), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n629), .A2(new_n592), .A3(new_n676), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n698), .B1(new_n549), .B2(new_n550), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n614), .A2(new_n579), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n538), .A2(new_n528), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(new_n701), .A3(new_n578), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n701), .A2(new_n700), .A3(KEYINPUT30), .A4(new_n578), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n521), .A2(new_n359), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n614), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n477), .A2(new_n582), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT93), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n477), .A2(KEYINPUT93), .A3(new_n582), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n708), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n675), .B1(new_n706), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT31), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n714), .A2(new_n715), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n699), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n697), .B1(new_n719), .B2(new_n682), .ZN(new_n720));
  INV_X1    g0520(.A(new_n698), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n551), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n718), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n722), .A2(new_n716), .A3(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n724), .A2(KEYINPUT94), .A3(G330), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n720), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n652), .A2(KEYINPUT26), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n658), .A2(new_n653), .A3(new_n536), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n727), .A2(new_n661), .A3(new_n728), .ZN(new_n729));
  AOI211_X1 g0529(.A(new_n500), .B(new_n523), .C1(new_n511), .C2(new_n267), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n528), .A2(new_n644), .A3(G200), .ZN(new_n731));
  OAI21_X1  g0531(.A(KEYINPUT87), .B1(new_n521), .B2(new_n375), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n730), .A2(new_n731), .A3(new_n522), .A4(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n589), .A2(new_n588), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n733), .B(new_n661), .C1(new_n573), .C2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n735), .B1(new_n679), .B2(new_n584), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n543), .B(new_n497), .C1(new_n544), .C2(new_n340), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n494), .B1(new_n477), .B2(G200), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n739), .A2(new_n495), .B1(new_n542), .B2(new_n545), .ZN(new_n740));
  AND3_X1   g0540(.A1(new_n736), .A2(new_n740), .A3(KEYINPUT95), .ZN(new_n741));
  AOI21_X1  g0541(.A(KEYINPUT95), .B1(new_n736), .B2(new_n740), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n729), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n743), .A2(KEYINPUT29), .A3(new_n676), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n654), .A2(new_n657), .A3(new_n659), .ZN(new_n745));
  INV_X1    g0545(.A(new_n661), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(new_n736), .B2(new_n740), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n675), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n744), .B1(KEYINPUT29), .B2(new_n748), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n726), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n696), .B1(new_n750), .B2(G1), .ZN(G364));
  INV_X1    g0551(.A(new_n681), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G330), .ZN(new_n753));
  INV_X1    g0553(.A(G13), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n207), .B1(new_n755), .B2(G45), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n692), .A2(new_n757), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n753), .A2(new_n683), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT96), .ZN(new_n760));
  INV_X1    g0560(.A(new_n758), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n227), .B1(G20), .B2(new_n539), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n691), .A2(new_n328), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n767), .A2(G355), .B1(new_n595), .B2(new_n691), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT97), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n226), .A2(new_n296), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n691), .A2(new_n285), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n770), .B(new_n771), .C1(new_n250), .C2(new_n296), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n766), .B1(new_n773), .B2(KEYINPUT98), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n774), .B1(KEYINPUT98), .B2(new_n773), .ZN(new_n775));
  OR3_X1    g0575(.A1(new_n208), .A2(KEYINPUT99), .A3(G190), .ZN(new_n776));
  OAI21_X1  g0576(.A(KEYINPUT99), .B1(new_n208), .B2(G190), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n375), .A2(G179), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n401), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n778), .A2(G20), .A3(G190), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G87), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n358), .A2(new_n208), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G190), .A2(G200), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n285), .B(new_n783), .C1(new_n787), .C2(new_n287), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n585), .A2(G200), .ZN(new_n789));
  AND2_X1   g0589(.A1(new_n784), .A2(new_n789), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n780), .B(new_n788), .C1(G58), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n579), .A2(new_n375), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT100), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n793), .A2(new_n777), .A3(new_n776), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G159), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n793), .A2(G190), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n208), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n791), .B1(KEYINPUT32), .B2(new_n796), .C1(new_n480), .C2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n784), .A2(new_n585), .A3(G200), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n796), .A2(KEYINPUT32), .B1(new_n801), .B2(G68), .ZN(new_n802));
  NOR4_X1   g0602(.A1(new_n358), .A2(new_n208), .A3(new_n585), .A4(new_n375), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n802), .B1(new_n244), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(KEYINPUT33), .B(G317), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n801), .A2(new_n806), .B1(new_n790), .B2(G322), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT101), .Z(new_n808));
  INV_X1    g0608(.A(new_n798), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n809), .A2(G294), .B1(G326), .B2(new_n803), .ZN(new_n810));
  INV_X1    g0610(.A(new_n779), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G283), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n285), .B1(new_n782), .B2(G303), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n795), .A2(G329), .B1(G311), .B2(new_n786), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n810), .A2(new_n812), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n799), .A2(new_n805), .B1(new_n808), .B2(new_n815), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n761), .B(new_n775), .C1(new_n765), .C2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n764), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n752), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n760), .A2(new_n819), .ZN(G396));
  NAND2_X1  g0620(.A1(new_n720), .A2(new_n725), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n398), .A2(new_n676), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n412), .A2(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n406), .A2(KEYINPUT72), .B1(new_n358), .B2(new_n410), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n417), .B1(new_n824), .B2(new_n409), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n823), .B1(new_n825), .B2(new_n822), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT102), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(new_n748), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n828), .A2(KEYINPUT103), .ZN(new_n829));
  INV_X1    g0629(.A(new_n826), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n676), .B(new_n830), .C1(new_n660), .C2(new_n665), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n828), .A2(KEYINPUT103), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n829), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT104), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(new_n834), .B2(new_n821), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n833), .A2(new_n726), .A3(KEYINPUT104), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n761), .B1(new_n821), .B2(new_n834), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n765), .A2(new_n762), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n761), .B1(new_n287), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n765), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n285), .B1(new_n782), .B2(G107), .ZN(new_n842));
  INV_X1    g0642(.A(G311), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n842), .B1(new_n843), .B2(new_n794), .C1(new_n798), .C2(new_n480), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n811), .A2(G87), .ZN(new_n845));
  INV_X1    g0645(.A(new_n790), .ZN(new_n846));
  INV_X1    g0646(.A(G294), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n845), .B1(new_n846), .B2(new_n847), .C1(new_n595), .C2(new_n787), .ZN(new_n848));
  INV_X1    g0648(.A(G303), .ZN(new_n849));
  INV_X1    g0649(.A(G283), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n804), .A2(new_n849), .B1(new_n800), .B2(new_n850), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n844), .A2(new_n848), .A3(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(G143), .A2(new_n790), .B1(new_n786), .B2(G159), .ZN(new_n853));
  INV_X1    g0653(.A(G137), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n853), .B1(new_n854), .B2(new_n804), .C1(new_n255), .C2(new_n800), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT34), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n811), .A2(G68), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n328), .B1(new_n782), .B2(G50), .ZN(new_n858));
  INV_X1    g0658(.A(G132), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n857), .B(new_n858), .C1(new_n794), .C2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(new_n809), .B2(G58), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n852), .B1(new_n856), .B2(new_n861), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n840), .B1(new_n841), .B2(new_n862), .C1(new_n830), .C2(new_n763), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n838), .A2(new_n863), .ZN(G384));
  NOR2_X1   g0664(.A1(new_n755), .A2(new_n207), .ZN(new_n865));
  INV_X1    g0665(.A(new_n673), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n636), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n344), .B1(KEYINPUT16), .B2(new_n343), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n368), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n371), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n866), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n870), .A2(new_n871), .A3(new_n378), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT37), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n369), .A2(KEYINPUT107), .A3(new_n371), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n369), .A2(new_n866), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n874), .A2(new_n378), .A3(new_n875), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n367), .A2(new_n368), .B1(new_n360), .B2(new_n357), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n873), .B1(new_n877), .B2(KEYINPUT107), .ZN(new_n878));
  OAI22_X1  g0678(.A1(new_n872), .A2(new_n873), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n871), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n373), .B2(new_n382), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n879), .A2(new_n881), .A3(KEYINPUT38), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n884), .A2(KEYINPUT39), .A3(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT108), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n377), .A2(new_n367), .A3(new_n368), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n673), .B1(new_n367), .B2(new_n368), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n888), .A2(new_n877), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n887), .B1(new_n890), .B2(new_n873), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n369), .A2(new_n371), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT107), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT37), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n894), .A2(new_n378), .A3(new_n874), .A4(new_n875), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n892), .A2(new_n875), .A3(new_n378), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(KEYINPUT108), .A3(KEYINPUT37), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n891), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n875), .B1(new_n636), .B2(new_n638), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n883), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n885), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT39), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n886), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n450), .A2(new_n675), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n867), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n429), .A2(new_n675), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n450), .A2(new_n453), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n906), .B1(new_n450), .B2(new_n453), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT105), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n675), .B(new_n826), .C1(new_n745), .C2(new_n747), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n412), .A2(new_n675), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n912), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n831), .A2(KEYINPUT105), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n909), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT106), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n884), .A2(new_n885), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n916), .B2(new_n917), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n905), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  OR2_X1    g0722(.A1(new_n749), .A2(new_n456), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n643), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n922), .B(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n830), .B1(new_n907), .B2(new_n908), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n718), .B1(new_n551), .B2(new_n721), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT109), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT31), .B1(new_n714), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n928), .B2(new_n714), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n926), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n362), .A2(KEYINPUT90), .A3(new_n372), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT90), .B1(new_n362), .B2(new_n372), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n638), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n889), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n891), .A2(new_n895), .A3(new_n897), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT38), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n885), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n931), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT40), .B1(new_n884), .B2(new_n885), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n939), .A2(KEYINPUT40), .B1(new_n931), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n456), .B1(new_n927), .B2(new_n930), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n682), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n943), .B2(new_n942), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n865), .B1(new_n925), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n925), .B2(new_n945), .ZN(new_n947));
  INV_X1    g0747(.A(new_n489), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n948), .A2(KEYINPUT35), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(KEYINPUT35), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n949), .A2(G116), .A3(new_n228), .A4(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT36), .ZN(new_n952));
  OAI21_X1  g0752(.A(G77), .B1(new_n261), .B2(new_n246), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n245), .B1(new_n225), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(G1), .A3(new_n754), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n947), .A2(new_n952), .A3(new_n955), .ZN(G367));
  OAI21_X1  g0756(.A(new_n740), .B1(new_n493), .B2(new_n676), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n650), .A2(new_n545), .A3(new_n651), .A4(new_n675), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n688), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n960), .A2(KEYINPUT42), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n957), .A2(new_n958), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n546), .B1(new_n962), .B2(new_n584), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n676), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n960), .A2(KEYINPUT42), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n966), .A2(KEYINPUT110), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT110), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(new_n964), .B2(new_n965), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n961), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(KEYINPUT111), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT111), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n972), .B(new_n961), .C1(new_n967), .C2(new_n969), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n648), .B1(new_n730), .B2(new_n676), .ZN(new_n974));
  OR3_X1    g0774(.A1(new_n661), .A2(new_n730), .A3(new_n676), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT43), .Z(new_n977));
  NAND3_X1  g0777(.A1(new_n971), .A2(new_n973), .A3(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(new_n971), .B2(new_n973), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n979), .A2(new_n982), .B1(new_n686), .B2(new_n962), .ZN(new_n983));
  INV_X1    g0783(.A(new_n982), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n686), .A2(new_n962), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n984), .A2(new_n985), .A3(new_n978), .ZN(new_n986));
  INV_X1    g0786(.A(new_n750), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n689), .A2(new_n959), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT45), .Z(new_n989));
  NOR2_X1   g0789(.A1(new_n689), .A2(new_n959), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT44), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(new_n686), .ZN(new_n993));
  INV_X1    g0793(.A(new_n688), .ZN(new_n994));
  INV_X1    g0794(.A(new_n687), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n994), .B1(new_n685), .B2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n683), .B(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n987), .B1(new_n993), .B2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n692), .B(KEYINPUT41), .Z(new_n999));
  OAI21_X1  g0799(.A(new_n756), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n983), .A2(new_n986), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n771), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n766), .B1(new_n211), .B2(new_n392), .C1(new_n1002), .C2(new_n239), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n1003), .A2(new_n758), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n779), .A2(new_n287), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n809), .A2(G68), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n337), .B2(new_n800), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n846), .A2(new_n255), .B1(new_n854), .B2(new_n794), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n328), .B1(new_n782), .B2(G58), .ZN(new_n1009));
  INV_X1    g0809(.A(G143), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1009), .B1(new_n804), .B2(new_n1010), .C1(new_n787), .C2(new_n244), .ZN(new_n1011));
  OR4_X1    g0811(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .A4(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n795), .A2(G317), .B1(G97), .B2(new_n811), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n850), .B2(new_n787), .C1(new_n849), .C2(new_n846), .ZN(new_n1014));
  AOI21_X1  g0814(.A(KEYINPUT46), .B1(new_n782), .B2(G116), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n782), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n328), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1015), .B(new_n1017), .C1(G294), .C2(new_n801), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n401), .B2(new_n798), .C1(new_n843), .C2(new_n804), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1012), .B1(new_n1014), .B2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT47), .Z(new_n1021));
  OAI221_X1 g0821(.A(new_n1004), .B1(new_n818), .B2(new_n976), .C1(new_n1021), .C2(new_n841), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1001), .A2(new_n1022), .ZN(G387));
  NAND2_X1  g0823(.A1(new_n997), .A2(new_n757), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n767), .A2(new_n693), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(G107), .B2(new_n211), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1002), .B1(new_n236), .B2(G45), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n258), .A2(G50), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT50), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n296), .B1(new_n246), .B2(new_n287), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(new_n693), .B2(KEYINPUT112), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1029), .B(new_n1031), .C1(KEYINPUT112), .C2(new_n693), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1026), .B1(new_n1027), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n766), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n758), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n787), .A2(new_n246), .B1(new_n255), .B2(new_n794), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(G50), .B2(new_n790), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n782), .A2(G77), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1038), .B(new_n285), .C1(new_n480), .C2(new_n779), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n263), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1039), .B1(new_n1040), .B2(new_n801), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n809), .A2(new_n499), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n803), .A2(G159), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1037), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n285), .B1(new_n795), .B2(G326), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G303), .A2(new_n786), .B1(new_n790), .B2(G317), .ZN(new_n1046));
  XOR2_X1   g0846(.A(KEYINPUT113), .B(G322), .Z(new_n1047));
  NAND2_X1  g0847(.A1(new_n803), .A2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1046), .B(new_n1048), .C1(new_n843), .C2(new_n800), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT114), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1050), .A2(KEYINPUT48), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(KEYINPUT48), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n809), .A2(G283), .B1(G294), .B2(new_n782), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT49), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1045), .B1(new_n595), .B2(new_n779), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1054), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1057), .A2(KEYINPUT49), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1044), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1035), .B1(new_n1059), .B2(new_n765), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT115), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n685), .B2(new_n818), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n750), .A2(new_n997), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n692), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n750), .A2(new_n997), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1024), .B1(new_n1062), .B2(new_n1064), .C1(new_n1066), .C2(new_n1067), .ZN(G393));
  NAND2_X1  g0868(.A1(new_n993), .A2(new_n757), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n766), .B1(new_n480), .B2(new_n211), .C1(new_n1002), .C2(new_n243), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n758), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n790), .A2(G159), .B1(G150), .B2(new_n803), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT51), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n809), .A2(G77), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n244), .B2(new_n800), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n845), .B(new_n285), .C1(new_n246), .C2(new_n781), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n787), .A2(new_n258), .B1(new_n1010), .B2(new_n794), .ZN(new_n1077));
  OR4_X1    g0877(.A1(new_n1073), .A2(new_n1075), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n809), .A2(G116), .B1(G294), .B2(new_n786), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n849), .B2(new_n800), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT116), .Z(new_n1081));
  AOI22_X1  g0881(.A1(new_n790), .A2(G311), .B1(G317), .B2(new_n803), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT52), .Z(new_n1083));
  INV_X1    g0883(.A(new_n780), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n795), .A2(new_n1047), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n285), .B1(new_n782), .B2(G283), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .A4(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1078), .B1(new_n1081), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1071), .B1(new_n1088), .B2(new_n765), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n959), .B2(new_n818), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1069), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n993), .A2(new_n750), .A3(new_n997), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n686), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n992), .B(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n1065), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1092), .A2(new_n692), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT117), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1092), .A2(new_n1095), .A3(KEYINPUT117), .A4(new_n692), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1091), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(G390));
  INV_X1    g0901(.A(new_n909), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n910), .B(new_n912), .C1(new_n748), .C2(new_n830), .ZN(new_n1103));
  AOI21_X1  g0903(.A(KEYINPUT105), .B1(new_n831), .B2(new_n914), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1102), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n904), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n902), .B1(new_n937), .B2(new_n938), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n884), .A2(KEYINPUT39), .A3(new_n885), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1105), .A2(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1106), .B1(new_n937), .B2(new_n938), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n743), .A2(new_n676), .A3(new_n830), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n909), .B1(new_n1111), .B2(new_n914), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n826), .B(new_n909), .C1(new_n720), .C2(new_n725), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n1109), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n682), .B1(new_n927), .B2(new_n930), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n926), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n382), .B1(new_n634), .B2(new_n635), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n936), .B1(new_n875), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n938), .B1(new_n1120), .B2(new_n883), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1108), .B1(new_n1121), .B2(KEYINPUT39), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n916), .B2(new_n904), .ZN(new_n1123));
  OR2_X1    g0923(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1118), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1115), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n757), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n839), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n758), .B1(new_n1040), .B2(new_n1128), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n787), .A2(new_n480), .B1(new_n847), .B2(new_n794), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(G116), .B2(new_n790), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n857), .A2(new_n328), .A3(new_n783), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n801), .A2(G107), .B1(G283), .B2(new_n803), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1131), .A2(new_n1074), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n798), .A2(new_n337), .B1(new_n854), .B2(new_n800), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G128), .B2(new_n803), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n790), .A2(G132), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n781), .A2(new_n255), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT53), .ZN(new_n1139));
  XOR2_X1   g0939(.A(KEYINPUT54), .B(G143), .Z(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT119), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n786), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1136), .A2(new_n1137), .A3(new_n1139), .A4(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(G125), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n285), .B1(new_n244), .B2(new_n779), .C1(new_n794), .C2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT120), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1134), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1129), .B1(new_n1147), .B2(new_n765), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(new_n903), .B2(new_n763), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1127), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n826), .B1(new_n720), .B2(new_n725), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1118), .B1(new_n1151), .B2(new_n1102), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n913), .A2(new_n915), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n821), .A2(new_n830), .A3(new_n1102), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1111), .A2(new_n914), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1116), .A2(new_n827), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1156), .B1(new_n1157), .B2(new_n909), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1154), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n457), .A2(new_n1116), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n643), .A2(new_n923), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1117), .B(new_n1116), .C1(new_n1109), .C2(new_n1113), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n904), .B1(new_n1153), .B2(new_n1102), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1124), .B(new_n1155), .C1(new_n1165), .C2(new_n903), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1160), .A2(new_n1163), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n692), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1162), .B1(new_n1154), .B2(new_n1159), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1168), .B1(new_n1126), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1167), .B1(new_n1170), .B2(KEYINPUT118), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1113), .B1(new_n1173), .B2(new_n1122), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1166), .B1(new_n1174), .B2(new_n1118), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n692), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT118), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1150), .B1(new_n1171), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(G378));
  INV_X1    g0980(.A(new_n386), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n308), .A2(new_n313), .A3(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n277), .A2(new_n673), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1183), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n308), .A2(new_n313), .A3(new_n1181), .A4(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1184), .A2(new_n1186), .A3(new_n1188), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n1190), .A2(KEYINPUT121), .A3(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n941), .B2(new_n682), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1190), .A2(KEYINPUT121), .A3(new_n1191), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT40), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n901), .B2(new_n931), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n940), .A2(new_n931), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1194), .B(G330), .C1(new_n1196), .C2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1193), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n922), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT122), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1105), .A2(KEYINPUT106), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1202), .A2(new_n918), .A3(new_n920), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1193), .A2(new_n1203), .A3(new_n1198), .A4(new_n905), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1200), .A2(new_n1201), .A3(new_n1204), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1152), .A2(new_n1153), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1163), .B1(new_n1175), .B2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1199), .A2(new_n922), .A3(KEYINPUT122), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1205), .A2(new_n1207), .A3(KEYINPUT57), .A4(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n692), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(KEYINPUT123), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT123), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1209), .A2(new_n1212), .A3(new_n692), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1200), .A2(new_n1204), .ZN(new_n1214));
  AOI21_X1  g1014(.A(KEYINPUT57), .B1(new_n1207), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1211), .A2(new_n1213), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1214), .A2(new_n757), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1190), .A2(new_n762), .A3(new_n1191), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n285), .A2(G41), .ZN(new_n1220));
  AOI211_X1 g1020(.A(G50), .B(new_n1220), .C1(new_n256), .C2(new_n295), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n846), .A2(new_n401), .B1(new_n850), .B2(new_n794), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n499), .B2(new_n786), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1038), .A2(new_n1220), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n779), .A2(new_n261), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n801), .A2(G97), .B1(G116), .B2(new_n803), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1223), .A2(new_n1006), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT58), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1221), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n798), .A2(new_n255), .B1(new_n859), .B2(new_n800), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1141), .A2(new_n782), .B1(new_n790), .B2(G128), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n854), .B2(new_n787), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1231), .B(new_n1233), .C1(G125), .C2(new_n803), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1235), .A2(KEYINPUT59), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n256), .B(new_n295), .C1(new_n779), .C2(new_n337), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n795), .B2(G124), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT59), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1238), .B1(new_n1234), .B2(new_n1239), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n1230), .B1(new_n1229), .B2(new_n1228), .C1(new_n1236), .C2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n765), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n761), .B1(new_n244), .B2(new_n839), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1219), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1218), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1217), .A2(new_n1246), .ZN(G375));
  INV_X1    g1047(.A(new_n999), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1206), .A2(new_n1162), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1172), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n909), .A2(new_n762), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n758), .B1(G68), .B2(new_n1128), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n809), .A2(G50), .B1(new_n801), .B2(new_n1141), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n328), .B(new_n1225), .C1(G159), .C2(new_n782), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1253), .B(new_n1254), .C1(new_n859), .C2(new_n804), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n795), .A2(G128), .B1(G137), .B2(new_n790), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n255), .B2(new_n787), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n795), .A2(G303), .B1(G283), .B2(new_n790), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n401), .B2(new_n787), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n801), .A2(G116), .B1(G294), .B2(new_n803), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n285), .B(new_n1005), .C1(G97), .C2(new_n782), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1042), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n1255), .A2(new_n1257), .B1(new_n1259), .B2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1252), .B1(new_n1263), .B2(new_n765), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n1160), .A2(new_n757), .B1(new_n1251), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1250), .A2(new_n1265), .ZN(G381));
  NOR3_X1   g1066(.A1(G384), .A2(G393), .A3(G396), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1267), .A2(new_n1100), .A3(new_n1001), .A4(new_n1022), .ZN(new_n1268));
  OR4_X1    g1068(.A1(G378), .A2(G375), .A3(G381), .A4(new_n1268), .ZN(G407));
  NAND2_X1  g1069(.A1(new_n674), .A2(G213), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1179), .A2(new_n1271), .ZN(new_n1272));
  OAI211_X1 g1072(.A(G407), .B(G213), .C1(G375), .C2(new_n1272), .ZN(G409));
  INV_X1    g1073(.A(KEYINPUT124), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1215), .B1(new_n1210), .B2(KEYINPUT123), .ZN(new_n1275));
  AOI211_X1 g1075(.A(new_n1179), .B(new_n1245), .C1(new_n1275), .C2(new_n1213), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1205), .A2(new_n757), .A3(new_n1208), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1207), .A2(new_n1214), .A3(new_n1248), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1277), .A2(new_n1278), .A3(new_n1244), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(G378), .A2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1274), .B1(new_n1276), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT60), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1249), .B1(new_n1169), .B2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1206), .A2(KEYINPUT60), .A3(new_n1162), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1283), .A2(new_n692), .A3(new_n1284), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1285), .A2(new_n1265), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT125), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n838), .A2(new_n1288), .A3(new_n863), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1286), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1287), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1291), .B1(new_n1286), .B2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1217), .A2(G378), .A3(new_n1246), .ZN(new_n1295));
  OR2_X1    g1095(.A1(G378), .A2(new_n1279), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1295), .A2(KEYINPUT124), .A3(new_n1296), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1281), .A2(new_n1270), .A3(new_n1294), .A4(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT63), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(KEYINPUT126), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT126), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1298), .A2(new_n1302), .A3(new_n1299), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT127), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(G390), .A2(new_n1022), .A3(new_n1001), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(G387), .A2(new_n1100), .ZN(new_n1306));
  XOR2_X1   g1106(.A(G393), .B(G396), .Z(new_n1307));
  AND4_X1   g1107(.A1(new_n1304), .A2(new_n1305), .A3(new_n1306), .A4(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(KEYINPUT127), .B1(G387), .B2(new_n1100), .ZN(new_n1309));
  AOI22_X1  g1109(.A1(new_n1309), .A2(new_n1307), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1310));
  NOR3_X1   g1110(.A1(new_n1308), .A2(new_n1310), .A3(KEYINPUT61), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1293), .A2(new_n1299), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1312), .B(new_n1270), .C1(new_n1276), .C2(new_n1280), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1311), .A2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1281), .A2(new_n1270), .A3(new_n1297), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1271), .A2(G2897), .ZN(new_n1316));
  XNOR2_X1  g1116(.A(new_n1293), .B(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1314), .B1(new_n1315), .B2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1301), .A2(new_n1303), .A3(new_n1318), .ZN(new_n1319));
  OR2_X1    g1119(.A1(new_n1308), .A2(new_n1310), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1271), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT62), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1293), .A2(new_n1322), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1321), .A2(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1324), .B1(new_n1298), .B2(new_n1322), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT61), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1317), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1326), .B1(new_n1327), .B2(new_n1321), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1320), .B1(new_n1325), .B2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1319), .A2(new_n1329), .ZN(G405));
  XNOR2_X1  g1130(.A(new_n1320), .B(new_n1294), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(G375), .A2(new_n1179), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n1295), .ZN(new_n1333));
  XNOR2_X1  g1133(.A(new_n1331), .B(new_n1333), .ZN(G402));
endmodule


