//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n555, new_n556, new_n557, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n610, new_n612,
    new_n613, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT66), .Z(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT67), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n464), .A2(G137), .A3(new_n463), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n467), .A2(new_n472), .ZN(G160));
  OAI21_X1  g048(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(G112), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n474), .B1(new_n475), .B2(G2105), .ZN(new_n476));
  AND2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(new_n463), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n476), .B1(new_n480), .B2(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n479), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  OAI21_X1  g060(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n487), .B1(new_n463), .B2(G114), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n489), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n486), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  AND2_X1   g066(.A1(G126), .A2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n492), .B1(new_n477), .B2(new_n478), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(KEYINPUT68), .B(new_n492), .C1(new_n477), .C2(new_n478), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n491), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(G138), .B(new_n463), .C1(new_n477), .C2(new_n478), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n464), .A2(new_n500), .A3(G138), .A4(new_n463), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AND2_X1   g077(.A1(new_n497), .A2(new_n502), .ZN(G164));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT70), .A3(KEYINPUT5), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n509), .A2(G88), .A3(new_n511), .A4(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(G50), .A3(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n510), .B1(new_n506), .B2(new_n508), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n516), .B1(new_n517), .B2(G62), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n513), .B(new_n514), .C1(new_n518), .C2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  NAND2_X1  g096(.A1(new_n517), .A2(new_n512), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G89), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n525));
  XOR2_X1   g100(.A(KEYINPUT71), .B(KEYINPUT7), .Z(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n526), .B(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n512), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G51), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n524), .A2(new_n525), .A3(new_n528), .A4(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n522), .A2(new_n534), .B1(new_n535), .B2(new_n529), .ZN(new_n536));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n509), .A2(new_n511), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G651), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n536), .B1(new_n541), .B2(KEYINPUT72), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT72), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n540), .A2(new_n543), .A3(G651), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  AOI22_X1  g121(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(new_n519), .ZN(new_n548));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n522), .A2(new_n549), .B1(new_n550), .B2(new_n529), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(new_n557));
  XOR2_X1   g132(.A(new_n557), .B(KEYINPUT73), .Z(G188));
  INV_X1    g133(.A(KEYINPUT74), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n512), .A2(G53), .A3(G543), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n523), .A2(G91), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n517), .A2(G65), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n519), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n559), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n566), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n568), .A2(new_n561), .A3(KEYINPUT74), .A4(new_n562), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(G299));
  NAND2_X1  g146(.A1(new_n530), .A2(G49), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n573));
  INV_X1    g148(.A(G87), .ZN(new_n574));
  OAI211_X1 g149(.A(new_n572), .B(new_n573), .C1(new_n574), .C2(new_n522), .ZN(G288));
  NAND3_X1  g150(.A1(new_n509), .A2(G61), .A3(new_n511), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n519), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n509), .A2(G86), .A3(new_n511), .A4(new_n512), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n512), .A2(G48), .A3(G543), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n519), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  INV_X1    g161(.A(G47), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n522), .A2(new_n586), .B1(new_n587), .B2(new_n529), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT75), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n523), .A2(new_n592), .A3(G92), .ZN(new_n593));
  INV_X1    g168(.A(G92), .ZN(new_n594));
  OAI21_X1  g169(.A(KEYINPUT75), .B1(new_n522), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n593), .A2(KEYINPUT10), .A3(new_n595), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n538), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(G54), .B2(new_n530), .ZN(new_n603));
  AND3_X1   g178(.A1(new_n598), .A2(new_n599), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n591), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n591), .B1(new_n604), .B2(G868), .ZN(G321));
  NAND2_X1  g181(.A1(G286), .A2(G868), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(new_n570), .B2(G868), .ZN(G280));
  XOR2_X1   g183(.A(G280), .B(KEYINPUT76), .Z(G297));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n604), .B1(new_n610), .B2(G860), .ZN(G148));
  NAND2_X1  g186(.A1(new_n604), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g189(.A(KEYINPUT77), .B(KEYINPUT11), .ZN(new_n615));
  XNOR2_X1  g190(.A(G323), .B(new_n615), .ZN(G282));
  NAND2_X1  g191(.A1(new_n482), .A2(G135), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT78), .ZN(new_n618));
  OAI21_X1  g193(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n619));
  INV_X1    g194(.A(G111), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G2105), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(new_n480), .B2(G123), .ZN(new_n622));
  AND2_X1   g197(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n624), .A2(G2096), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n464), .A2(new_n470), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(G2100), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(G2100), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n624), .A2(G2096), .ZN(new_n632));
  NAND4_X1  g207(.A1(new_n625), .A2(new_n630), .A3(new_n631), .A4(new_n632), .ZN(G156));
  INV_X1    g208(.A(KEYINPUT14), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n634), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(new_n637), .B2(new_n636), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2451), .B(G2454), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n639), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  AND3_X1   g222(.A1(new_n646), .A2(G14), .A3(new_n647), .ZN(G401));
  XOR2_X1   g223(.A(G2072), .B(G2078), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT79), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT17), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2084), .B(G2090), .ZN(new_n653));
  NOR3_X1   g228(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n653), .B1(new_n650), .B2(new_n652), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n655), .B1(new_n651), .B2(new_n652), .ZN(new_n656));
  INV_X1    g231(.A(new_n652), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n657), .A2(new_n653), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n650), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT18), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n654), .A2(new_n656), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(G2096), .Z(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT80), .B(G2100), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1956), .B(G2474), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT20), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n668), .A2(new_n669), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n667), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n667), .B2(new_n673), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1991), .B(G1996), .Z(new_n677));
  XOR2_X1   g252(.A(new_n676), .B(new_n677), .Z(new_n678));
  XOR2_X1   g253(.A(KEYINPUT81), .B(KEYINPUT82), .Z(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1981), .B(G1986), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n678), .B(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(G229));
  INV_X1    g260(.A(G29), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G33), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT88), .B(KEYINPUT25), .Z(new_n688));
  NAND3_X1  g263(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(G139), .ZN(new_n691));
  INV_X1    g266(.A(new_n482), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  AOI22_X1  g268(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n694), .A2(new_n463), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n687), .B1(new_n696), .B2(new_n686), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT89), .ZN(new_n698));
  INV_X1    g273(.A(G2072), .ZN(new_n699));
  NOR2_X1   g274(.A1(G16), .A2(G19), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n552), .B2(G16), .ZN(new_n701));
  OAI22_X1  g276(.A1(new_n698), .A2(new_n699), .B1(G1341), .B2(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(G27), .A2(G29), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(G164), .B2(G29), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(G2078), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT30), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n706), .A2(G28), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n686), .B1(new_n706), .B2(G28), .ZN(new_n708));
  AND2_X1   g283(.A1(KEYINPUT31), .A2(G11), .ZN(new_n709));
  NOR2_X1   g284(.A1(KEYINPUT31), .A2(G11), .ZN(new_n710));
  OAI22_X1  g285(.A1(new_n707), .A2(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(new_n623), .B2(G29), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT24), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n686), .B1(new_n713), .B2(G34), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(KEYINPUT91), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n714), .A2(KEYINPUT91), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n713), .B2(G34), .ZN(new_n717));
  AOI22_X1  g292(.A1(G160), .A2(G29), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G2084), .ZN(new_n719));
  OR2_X1    g294(.A1(G104), .A2(G2105), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n720), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n721));
  OAI211_X1 g296(.A(G140), .B(new_n463), .C1(new_n477), .C2(new_n478), .ZN(new_n722));
  OAI211_X1 g297(.A(G128), .B(G2105), .C1(new_n477), .C2(new_n478), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G29), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n686), .A2(G26), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT28), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT87), .B(G2067), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n712), .A2(new_n719), .A3(new_n730), .ZN(new_n731));
  NOR3_X1   g306(.A1(new_n702), .A2(new_n705), .A3(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G16), .ZN(new_n733));
  OR3_X1    g308(.A1(G286), .A2(KEYINPUT95), .A3(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(G286), .A2(new_n733), .ZN(new_n735));
  OAI21_X1  g310(.A(KEYINPUT95), .B1(G16), .B2(G21), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n737), .A2(G1966), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G1341), .B2(new_n701), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n732), .B(new_n739), .C1(G1966), .C2(new_n737), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n470), .A2(G105), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT92), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G141), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(new_n692), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n480), .A2(G129), .ZN(new_n746));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(KEYINPUT26), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n747), .A2(KEYINPUT26), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n746), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n745), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT93), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(G29), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT94), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n754), .B(new_n755), .C1(G29), .C2(G32), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n755), .B2(new_n754), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT27), .B(G1996), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n686), .A2(G35), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT97), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G162), .B2(new_n686), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT29), .B(G2090), .Z(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(KEYINPUT96), .B1(new_n718), .B2(G2084), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR3_X1   g341(.A1(new_n718), .A2(KEYINPUT96), .A3(G2084), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n759), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n757), .A2(new_n758), .ZN(new_n770));
  NOR3_X1   g345(.A1(new_n740), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n604), .A2(G16), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G4), .B2(G16), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT86), .B(G1348), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n733), .A2(G20), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT23), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n570), .B2(new_n733), .ZN(new_n779));
  INV_X1    g354(.A(G1956), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n775), .A2(new_n776), .A3(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n698), .A2(new_n699), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT90), .Z(new_n785));
  NAND2_X1  g360(.A1(new_n733), .A2(G5), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G171), .B2(new_n733), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1961), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n771), .A2(new_n783), .A3(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(G6), .A2(G16), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n582), .B2(G16), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT32), .B(G1981), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n792), .B(new_n793), .Z(new_n794));
  AND2_X1   g369(.A1(new_n794), .A2(KEYINPUT85), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n794), .A2(KEYINPUT85), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n733), .A2(G22), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G166), .B2(new_n733), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G1971), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n733), .A2(G23), .ZN(new_n800));
  INV_X1    g375(.A(G288), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(new_n733), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT33), .B(G1976), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n802), .B(new_n803), .Z(new_n804));
  NOR4_X1   g379(.A1(new_n795), .A2(new_n796), .A3(new_n799), .A4(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT34), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  NOR2_X1   g383(.A1(G25), .A2(G29), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n480), .A2(G119), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n482), .A2(G131), .ZN(new_n811));
  OR2_X1    g386(.A1(G95), .A2(G2105), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n812), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n809), .B1(new_n815), .B2(G29), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT35), .B(G1991), .Z(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT83), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n816), .B(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n733), .A2(G24), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n589), .A2(KEYINPUT84), .ZN(new_n821));
  OAI21_X1  g396(.A(G16), .B1(new_n589), .B2(KEYINPUT84), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n819), .B1(new_n823), .B2(G1986), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G1986), .B2(new_n823), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n807), .A2(new_n808), .A3(new_n825), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n826), .A2(KEYINPUT36), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(KEYINPUT36), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n790), .B1(new_n827), .B2(new_n828), .ZN(G311));
  XNOR2_X1  g404(.A(new_n826), .B(KEYINPUT36), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n771), .A2(new_n789), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n830), .A2(new_n783), .A3(new_n831), .ZN(G150));
  AOI22_X1  g407(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n833), .A2(new_n519), .ZN(new_n834));
  INV_X1    g409(.A(G93), .ZN(new_n835));
  INV_X1    g410(.A(G55), .ZN(new_n836));
  OAI22_X1  g411(.A1(new_n522), .A2(new_n835), .B1(new_n836), .B2(new_n529), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n838));
  OR3_X1    g413(.A1(new_n834), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n834), .B2(new_n837), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n839), .A2(new_n552), .A3(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n834), .A2(new_n837), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n842), .B(new_n838), .C1(new_n548), .C2(new_n551), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n598), .A2(new_n599), .A3(new_n603), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n846), .A2(new_n610), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n845), .B(new_n847), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n850));
  NOR3_X1   g425(.A1(new_n849), .A2(new_n850), .A3(G860), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n842), .A2(G860), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT37), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n851), .A2(new_n853), .ZN(G145));
  INV_X1    g429(.A(KEYINPUT99), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n724), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n721), .A2(new_n722), .A3(new_n723), .A4(KEYINPUT99), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(G164), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n497), .A2(new_n502), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n860), .A2(new_n856), .A3(new_n857), .ZN(new_n861));
  AND3_X1   g436(.A1(new_n859), .A2(new_n751), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n751), .B1(new_n859), .B2(new_n861), .ZN(new_n863));
  OAI21_X1  g438(.A(KEYINPUT93), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n859), .A2(new_n861), .ZN(new_n865));
  INV_X1    g440(.A(new_n751), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n859), .A2(new_n751), .A3(new_n861), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n867), .A2(new_n752), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n864), .A2(new_n869), .A3(new_n696), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n862), .A2(new_n863), .ZN(new_n871));
  INV_X1    g446(.A(new_n696), .ZN(new_n872));
  AOI21_X1  g447(.A(KEYINPUT100), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n864), .A2(new_n869), .A3(KEYINPUT100), .A4(new_n696), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n480), .A2(G130), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n482), .A2(G142), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n463), .A2(G118), .ZN(new_n879));
  OAI21_X1  g454(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n877), .B(new_n878), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n881), .B(new_n627), .Z(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n815), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n876), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n874), .A2(new_n883), .A3(new_n875), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(KEYINPUT101), .A3(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n484), .B(G160), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n623), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n883), .B1(new_n874), .B2(new_n875), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(G37), .B1(new_n887), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n886), .A2(KEYINPUT102), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT102), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n874), .A2(new_n896), .A3(new_n883), .A4(new_n875), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n895), .A2(new_n885), .A3(new_n897), .A4(new_n890), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n891), .A2(new_n889), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n901), .A2(KEYINPUT103), .A3(new_n897), .A4(new_n895), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n894), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g479(.A(G868), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n842), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n612), .B(new_n844), .ZN(new_n907));
  NAND3_X1  g482(.A1(G299), .A2(KEYINPUT104), .A3(new_n846), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT104), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n570), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n567), .A2(KEYINPUT104), .A3(new_n569), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(new_n604), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n907), .A2(new_n908), .A3(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(KEYINPUT105), .ZN(new_n914));
  XNOR2_X1  g489(.A(G305), .B(new_n589), .ZN(new_n915));
  XNOR2_X1  g490(.A(G166), .B(G288), .ZN(new_n916));
  XOR2_X1   g491(.A(new_n915), .B(new_n916), .Z(new_n917));
  NAND2_X1  g492(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n920));
  XOR2_X1   g495(.A(new_n920), .B(KEYINPUT107), .Z(new_n921));
  XNOR2_X1  g496(.A(new_n919), .B(new_n921), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n567), .A2(KEYINPUT104), .A3(new_n569), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT104), .B1(new_n567), .B2(new_n569), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n923), .A2(new_n924), .A3(new_n846), .ZN(new_n925));
  NOR3_X1   g500(.A1(new_n604), .A2(new_n570), .A3(new_n909), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT41), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT41), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n912), .A2(new_n928), .A3(new_n908), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n914), .B(new_n922), .C1(new_n907), .C2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n922), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT105), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n913), .B(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n931), .A2(new_n907), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n932), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n906), .B1(new_n938), .B2(new_n905), .ZN(G295));
  OAI21_X1  g514(.A(new_n906), .B1(new_n938), .B2(new_n905), .ZN(G331));
  INV_X1    g515(.A(new_n917), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n912), .A2(new_n928), .A3(new_n908), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT109), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n528), .A2(new_n531), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n944), .A2(KEYINPUT108), .A3(new_n524), .A4(new_n525), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT108), .ZN(new_n946));
  NAND2_X1  g521(.A1(G286), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(G301), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(G168), .A2(new_n542), .A3(KEYINPUT108), .A4(new_n544), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n844), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n948), .A2(new_n949), .A3(new_n841), .A4(new_n843), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n943), .B(new_n953), .C1(new_n930), .C2(KEYINPUT109), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n912), .A2(new_n908), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n941), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n928), .B1(new_n912), .B2(new_n908), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n953), .B1(new_n942), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n960), .A2(new_n957), .A3(new_n941), .ZN(new_n961));
  INV_X1    g536(.A(G37), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT43), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n958), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n956), .B1(new_n930), .B2(new_n953), .ZN(new_n966));
  AOI21_X1  g541(.A(G37), .B1(new_n966), .B2(new_n941), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n941), .B1(new_n960), .B2(new_n957), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT43), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT44), .B1(new_n965), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n958), .A2(new_n963), .A3(KEYINPUT43), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n964), .B1(new_n967), .B2(new_n969), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n971), .A2(new_n975), .ZN(G397));
  INV_X1    g551(.A(G1384), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n860), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G125), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n466), .B1(new_n479), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(G2105), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n983), .A2(G40), .A3(new_n471), .A4(new_n468), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n986), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT46), .ZN(new_n988));
  INV_X1    g563(.A(G1996), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n988), .B1(new_n985), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G2067), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n724), .B(new_n991), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n751), .A2(new_n992), .ZN(new_n993));
  OAI22_X1  g568(.A1(new_n987), .A2(new_n990), .B1(new_n986), .B2(new_n993), .ZN(new_n994));
  XOR2_X1   g569(.A(new_n994), .B(KEYINPUT47), .Z(new_n995));
  NAND2_X1  g570(.A1(new_n753), .A2(new_n989), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n996), .B(new_n992), .C1(new_n989), .C2(new_n751), .ZN(new_n997));
  XOR2_X1   g572(.A(new_n814), .B(new_n817), .Z(new_n998));
  NOR2_X1   g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT48), .ZN(new_n1000));
  OR3_X1    g575(.A1(new_n986), .A2(G1986), .A3(G290), .ZN(new_n1001));
  OAI22_X1  g576(.A1(new_n999), .A2(new_n986), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1002), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n815), .A2(new_n817), .ZN(new_n1004));
  OAI22_X1  g579(.A1(new_n997), .A2(new_n1004), .B1(G2067), .B2(new_n724), .ZN(new_n1005));
  AOI211_X1 g580(.A(new_n995), .B(new_n1003), .C1(new_n985), .C2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n978), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n1008));
  AOI21_X1  g583(.A(G1384), .B1(new_n497), .B2(new_n502), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1008), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n984), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1007), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT120), .ZN(new_n1014));
  INV_X1    g589(.A(G1961), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT120), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1007), .A2(new_n1011), .A3(new_n1012), .A4(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1014), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n978), .A2(new_n979), .ZN(new_n1020));
  INV_X1    g595(.A(G40), .ZN(new_n1021));
  NOR3_X1   g596(.A1(new_n467), .A2(new_n472), .A3(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1022), .B1(new_n1009), .B2(KEYINPUT45), .ZN(new_n1023));
  OR4_X1    g598(.A1(new_n1019), .A2(new_n1020), .A3(new_n1023), .A4(G2078), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1018), .A2(KEYINPUT125), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n979), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1022), .B1(new_n1009), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT45), .ZN(new_n1028));
  AOI211_X1 g603(.A(new_n1028), .B(G1384), .C1(new_n497), .C2(new_n502), .ZN(new_n1029));
  OR2_X1    g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1019), .B1(new_n1030), .B2(G2078), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n1025), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT125), .B1(new_n1018), .B2(new_n1024), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(G301), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT49), .ZN(new_n1036));
  INV_X1    g611(.A(G1981), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n576), .A2(new_n577), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(G651), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n579), .A2(new_n580), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1037), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n578), .A2(new_n581), .A3(G1981), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1036), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G8), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1044), .B1(new_n1009), .B2(new_n1022), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1039), .A2(new_n1040), .A3(new_n1037), .ZN(new_n1047));
  OAI21_X1  g622(.A(G1981), .B1(new_n578), .B2(new_n581), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT113), .B1(new_n1049), .B2(new_n1036), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT113), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1047), .A2(new_n1048), .A3(new_n1051), .A4(KEYINPUT49), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1046), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n801), .A2(G1976), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n1045), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT52), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT112), .B(G1976), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT52), .B1(G288), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1054), .A2(new_n1045), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT116), .B1(new_n1053), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1046), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT52), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1065), .B1(new_n1054), .B2(new_n1045), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1055), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1066), .B1(new_n1067), .B2(new_n1058), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1064), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1061), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n509), .A2(G62), .A3(new_n511), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n519), .B1(new_n1072), .B2(new_n515), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n513), .A2(new_n514), .ZN(new_n1074));
  OAI211_X1 g649(.A(KEYINPUT55), .B(G8), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G2090), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1007), .A2(new_n1011), .A3(new_n1012), .A4(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G1971), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1082));
  AOI211_X1 g657(.A(new_n1044), .B(new_n1078), .C1(new_n1080), .C2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1022), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT115), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1087));
  OAI211_X1 g662(.A(KEYINPUT115), .B(new_n1022), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1086), .A2(new_n1087), .A3(new_n1079), .A4(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n1082), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(G8), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1083), .B1(new_n1091), .B2(new_n1078), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1071), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(G2084), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1007), .A2(new_n1011), .A3(new_n1012), .A4(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(G1966), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(new_n1097), .A3(G168), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(G8), .ZN(new_n1099));
  AOI21_X1  g674(.A(G168), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT51), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT62), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT51), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1098), .A2(new_n1103), .A3(G8), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1101), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT62), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1035), .A2(new_n1093), .A3(new_n1105), .A4(new_n1107), .ZN(new_n1108));
  AOI211_X1 g683(.A(new_n1044), .B(G286), .C1(new_n1095), .C2(new_n1097), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1071), .A2(new_n1092), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT63), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1044), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1113), .B(new_n1078), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1053), .A2(new_n1060), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1114), .A2(KEYINPUT63), .A3(new_n1115), .A4(new_n1109), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1042), .B(KEYINPUT114), .ZN(new_n1118));
  OR2_X1    g693(.A1(G288), .A2(G1976), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1118), .B1(new_n1053), .B2(new_n1119), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1120), .A2(new_n1045), .B1(new_n1115), .B2(new_n1083), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1108), .A2(new_n1117), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1093), .A2(new_n1106), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT61), .ZN(new_n1124));
  XOR2_X1   g699(.A(KEYINPUT56), .B(G2072), .Z(new_n1125));
  OAI21_X1  g700(.A(KEYINPUT117), .B1(new_n1030), .B2(new_n1125), .ZN(new_n1126));
  OR4_X1    g701(.A1(KEYINPUT117), .A2(new_n1027), .A3(new_n1029), .A4(new_n1125), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1126), .A2(new_n1127), .B1(new_n1128), .B2(new_n780), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n563), .A2(new_n566), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1130), .B(KEYINPUT57), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1124), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1128), .A2(new_n780), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT57), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1130), .B(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT121), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT121), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1131), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1135), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1009), .A2(new_n1022), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1143), .B(KEYINPUT118), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n991), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT119), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1014), .A2(new_n774), .A3(new_n1017), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1144), .A2(KEYINPUT119), .A3(new_n991), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT60), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n846), .A2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .A4(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n846), .A2(new_n1150), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n1132), .A2(new_n1142), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1133), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1124), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g732(.A(KEYINPUT58), .B(G1341), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1144), .A2(new_n1158), .ZN(new_n1159));
  XOR2_X1   g734(.A(KEYINPUT122), .B(G1996), .Z(new_n1160));
  NOR2_X1   g735(.A1(new_n1030), .A2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g736(.A(KEYINPUT123), .B(new_n552), .C1(new_n1159), .C2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT59), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1154), .A2(new_n1157), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1156), .A2(new_n846), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1167));
  AOI22_X1  g742(.A1(new_n1166), .A2(new_n1167), .B1(new_n1135), .B2(new_n1141), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1123), .B1(new_n1165), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT126), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1018), .A2(new_n1170), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1014), .A2(KEYINPUT126), .A3(new_n1015), .A4(new_n1017), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1030), .A2(G2078), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1174), .B(new_n1019), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(KEYINPUT127), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT127), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1173), .A2(new_n1178), .A3(new_n1175), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1177), .A2(G171), .A3(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT54), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1025), .A2(new_n1031), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1182), .A2(new_n1033), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1181), .B1(new_n1183), .B2(G301), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1173), .A2(G301), .A3(new_n1175), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1185), .B1(new_n1183), .B2(G301), .ZN(new_n1186));
  XOR2_X1   g761(.A(KEYINPUT124), .B(KEYINPUT54), .Z(new_n1187));
  AOI22_X1  g762(.A1(new_n1180), .A2(new_n1184), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1122), .B1(new_n1169), .B2(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n589), .B(G1986), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n986), .B1(new_n999), .B2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1006), .B1(new_n1189), .B2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g767(.A1(new_n461), .A2(G401), .ZN(new_n1194));
  NAND3_X1  g768(.A1(new_n664), .A2(new_n684), .A3(new_n1194), .ZN(new_n1195));
  NOR3_X1   g769(.A1(new_n942), .A2(new_n959), .A3(KEYINPUT109), .ZN(new_n1196));
  INV_X1    g770(.A(KEYINPUT109), .ZN(new_n1197));
  OAI21_X1  g771(.A(new_n953), .B1(new_n929), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g772(.A(new_n957), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g773(.A1(new_n1199), .A2(new_n917), .ZN(new_n1200));
  NAND3_X1  g774(.A1(new_n1200), .A2(new_n967), .A3(new_n964), .ZN(new_n1201));
  OAI21_X1  g775(.A(KEYINPUT43), .B1(new_n963), .B2(new_n968), .ZN(new_n1202));
  AOI21_X1  g776(.A(new_n1195), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  AND2_X1   g777(.A1(new_n1203), .A2(new_n903), .ZN(G308));
  NAND2_X1  g778(.A1(new_n1203), .A2(new_n903), .ZN(G225));
endmodule


