//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 1 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008;
  INV_X1    g000(.A(KEYINPUT23), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G128), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT23), .A3(G119), .ZN(new_n191));
  OAI211_X1 g005(.A(new_n189), .B(new_n191), .C1(G119), .C2(new_n190), .ZN(new_n192));
  XNOR2_X1  g006(.A(G119), .B(G128), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT24), .B(G110), .Z(new_n194));
  AOI22_X1  g008(.A1(new_n192), .A2(G110), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G125), .ZN(new_n196));
  NOR3_X1   g010(.A1(new_n196), .A2(KEYINPUT16), .A3(G140), .ZN(new_n197));
  XNOR2_X1  g011(.A(G125), .B(G140), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(KEYINPUT16), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(G146), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  AOI211_X1 g015(.A(new_n201), .B(new_n197), .C1(KEYINPUT16), .C2(new_n198), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n195), .B1(new_n200), .B2(new_n202), .ZN(new_n203));
  OAI22_X1  g017(.A1(new_n192), .A2(G110), .B1(new_n193), .B2(new_n194), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n199), .A2(G146), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT64), .B(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(new_n198), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n203), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G137), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT70), .ZN(new_n211));
  NAND2_X1  g025(.A1(G221), .A2(G234), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n211), .B1(new_n212), .B2(G953), .ZN(new_n213));
  INV_X1    g027(.A(G953), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n214), .A2(KEYINPUT70), .A3(G221), .A4(G234), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT22), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n216), .A2(KEYINPUT22), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n210), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n219), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(G137), .A3(new_n217), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n209), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n203), .A2(new_n220), .A3(new_n222), .A4(new_n208), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT25), .B1(new_n226), .B2(G902), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT25), .ZN(new_n228));
  INV_X1    g042(.A(G902), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n224), .A2(new_n228), .A3(new_n229), .A4(new_n225), .ZN(new_n230));
  NAND2_X1  g044(.A1(G217), .A2(G902), .ZN(new_n231));
  INV_X1    g045(.A(G217), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(G234), .ZN(new_n233));
  XOR2_X1   g047(.A(new_n233), .B(KEYINPUT69), .Z(new_n234));
  NAND3_X1  g048(.A1(new_n227), .A2(new_n230), .A3(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n234), .A2(G902), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n235), .B1(new_n226), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT30), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT11), .ZN(new_n240));
  INV_X1    g054(.A(G134), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n240), .B1(new_n241), .B2(G137), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(G137), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n210), .A2(KEYINPUT11), .A3(G134), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G131), .ZN(new_n246));
  INV_X1    g060(.A(G131), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n242), .A2(new_n244), .A3(new_n247), .A4(new_n243), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT64), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G146), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n251), .A2(new_n253), .A3(G143), .ZN(new_n254));
  INV_X1    g068(.A(G143), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G146), .ZN(new_n256));
  AND2_X1   g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n254), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n255), .A2(G146), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n251), .A2(new_n253), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n259), .B1(new_n260), .B2(new_n255), .ZN(new_n261));
  NOR2_X1   g075(.A1(KEYINPUT0), .A2(G128), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n258), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n250), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(G134), .B(G137), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT65), .B1(new_n267), .B2(new_n247), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n210), .A2(G134), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n243), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT65), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n271), .A3(G131), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n268), .A2(new_n272), .A3(new_n248), .ZN(new_n273));
  INV_X1    g087(.A(new_n259), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n274), .B1(new_n206), .B2(G143), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT1), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n276), .B1(new_n206), .B2(G143), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n275), .B1(new_n277), .B2(new_n190), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n254), .A2(new_n276), .A3(G128), .A4(new_n256), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n273), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n239), .B1(new_n266), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n190), .B1(new_n254), .B2(KEYINPUT1), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n279), .B1(new_n282), .B2(new_n261), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n283), .A2(new_n248), .A3(new_n268), .A4(new_n272), .ZN(new_n284));
  INV_X1    g098(.A(new_n265), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n249), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n284), .A2(new_n286), .A3(KEYINPUT30), .ZN(new_n287));
  XNOR2_X1  g101(.A(KEYINPUT2), .B(G113), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT66), .ZN(new_n290));
  XNOR2_X1  g104(.A(G116), .B(G119), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n291), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(KEYINPUT66), .A3(new_n288), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n281), .A2(new_n287), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT67), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n292), .A2(new_n294), .A3(KEYINPUT67), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n300), .A2(new_n284), .A3(new_n286), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT26), .B(G101), .ZN(new_n302));
  NOR2_X1   g116(.A1(G237), .A2(G953), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G210), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n302), .B(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n305), .B(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n296), .A2(new_n301), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT31), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT28), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n301), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n284), .A2(new_n286), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n295), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n300), .A2(new_n284), .A3(new_n286), .A4(KEYINPUT28), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n312), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n307), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT31), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n296), .A2(new_n318), .A3(new_n301), .A4(new_n308), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n310), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(G472), .A2(G902), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(KEYINPUT32), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT32), .B1(new_n320), .B2(new_n321), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n316), .A2(new_n307), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n308), .B1(new_n296), .B2(new_n301), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT29), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n313), .A2(new_n299), .A3(new_n298), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n312), .A2(new_n329), .A3(new_n315), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n308), .A2(KEYINPUT29), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n229), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(G472), .B1(new_n328), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n238), .B1(new_n325), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT9), .B(G234), .ZN(new_n335));
  OAI21_X1  g149(.A(G221), .B1(new_n335), .B2(G902), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G469), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(new_n229), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT3), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT71), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n340), .A2(KEYINPUT71), .ZN(new_n342));
  INV_X1    g156(.A(G107), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G104), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n341), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT73), .B(G101), .ZN(new_n346));
  INV_X1    g160(.A(G104), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G107), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n340), .A2(new_n343), .A3(KEYINPUT71), .A4(G104), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n345), .A2(new_n346), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT74), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n351), .B1(new_n343), .B2(G104), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n344), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n348), .A2(new_n351), .ZN(new_n354));
  OAI21_X1  g168(.A(G101), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n254), .A2(new_n256), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n190), .B1(new_n274), .B2(KEYINPUT1), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n279), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n350), .A2(new_n355), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n362), .A2(new_n361), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n360), .A2(new_n361), .B1(new_n363), .B2(new_n283), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT71), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n365), .A2(KEYINPUT3), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n347), .A2(G107), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(KEYINPUT3), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n349), .A2(new_n348), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT72), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT72), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n345), .A2(new_n372), .A3(new_n348), .A4(new_n349), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(G101), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(KEYINPUT4), .A3(new_n350), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT4), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n371), .A2(new_n373), .A3(new_n376), .A4(G101), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n375), .A2(new_n285), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n364), .A2(new_n250), .A3(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(G110), .B(G140), .ZN(new_n380));
  INV_X1    g194(.A(G227), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(G953), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n380), .B(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT75), .B1(new_n356), .B2(new_n283), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT75), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n362), .A2(new_n278), .A3(new_n387), .A4(new_n279), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n360), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(KEYINPUT12), .A3(new_n249), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT12), .B1(new_n389), .B2(new_n249), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT76), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n362), .A2(new_n278), .A3(new_n279), .ZN(new_n394));
  AOI22_X1  g208(.A1(new_n394), .A2(KEYINPUT75), .B1(new_n356), .B2(new_n359), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n250), .B1(new_n395), .B2(new_n388), .ZN(new_n396));
  NOR3_X1   g210(.A1(new_n396), .A2(KEYINPUT76), .A3(KEYINPUT12), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n385), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n364), .A2(new_n378), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n249), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n384), .B1(new_n400), .B2(new_n379), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(G902), .B1(new_n398), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n339), .B1(new_n403), .B2(new_n338), .ZN(new_n404));
  INV_X1    g218(.A(new_n379), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n250), .B1(new_n364), .B2(new_n378), .ZN(new_n406));
  NOR3_X1   g220(.A1(new_n405), .A2(new_n383), .A3(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n379), .B1(new_n393), .B2(new_n397), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n407), .B1(new_n408), .B2(new_n383), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G469), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n337), .B1(new_n404), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G122), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G116), .ZN(new_n413));
  INV_X1    g227(.A(G116), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G122), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n416), .A2(G107), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n255), .A2(G128), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n190), .A2(G143), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(new_n241), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n419), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G134), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n417), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT88), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n413), .B1(new_n415), .B2(KEYINPUT14), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT87), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n412), .A2(G116), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT14), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n415), .A2(KEYINPUT87), .A3(KEYINPUT14), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n425), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n424), .B1(new_n431), .B2(new_n343), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NOR3_X1   g247(.A1(new_n431), .A2(new_n424), .A3(new_n343), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n423), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n343), .B1(new_n413), .B2(new_n415), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n420), .B1(new_n417), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT13), .B1(new_n255), .B2(G128), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(KEYINPUT86), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT13), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n439), .B(new_n419), .C1(new_n440), .C2(new_n418), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n437), .B1(new_n441), .B2(G134), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT89), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n435), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n423), .ZN(new_n446));
  INV_X1    g260(.A(new_n431), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(KEYINPUT88), .A3(G107), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n446), .B1(new_n448), .B2(new_n432), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT89), .B1(new_n449), .B2(new_n442), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n335), .A2(new_n232), .A3(G953), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n445), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n451), .B1(new_n445), .B2(new_n450), .ZN(new_n453));
  OAI211_X1 g267(.A(KEYINPUT91), .B(new_n229), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G478), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT15), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n455), .B1(KEYINPUT90), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n457), .B1(KEYINPUT90), .B2(new_n456), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n454), .B(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n303), .A2(G143), .A3(G214), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(G143), .B1(new_n303), .B2(G214), .ZN(new_n463));
  OAI21_X1  g277(.A(G131), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n303), .A2(G214), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n255), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n247), .A3(new_n461), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT17), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n464), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT84), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n200), .A2(new_n202), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT84), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n464), .A2(new_n467), .A3(new_n472), .A4(new_n468), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n466), .A2(new_n461), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(KEYINPUT17), .A3(G131), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n470), .A2(new_n471), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(KEYINPUT18), .A2(G131), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n474), .B(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n207), .B1(new_n201), .B2(new_n198), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(G113), .B(G122), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT83), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n482), .B(new_n347), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n476), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT85), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n476), .A2(KEYINPUT85), .A3(new_n480), .A4(new_n483), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n476), .A2(new_n480), .ZN(new_n488));
  INV_X1    g302(.A(new_n483), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n486), .A2(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(G475), .B1(new_n490), .B2(G902), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT20), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n486), .A2(new_n487), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n464), .A2(new_n467), .ZN(new_n494));
  AND2_X1   g308(.A1(KEYINPUT82), .A2(KEYINPUT19), .ZN(new_n495));
  NOR2_X1   g309(.A1(KEYINPUT82), .A2(KEYINPUT19), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n198), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n497), .B1(new_n198), .B2(new_n496), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n494), .B(new_n205), .C1(new_n498), .C2(new_n260), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n480), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n489), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n493), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(G475), .A2(G902), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n492), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n486), .A2(new_n487), .B1(new_n489), .B2(new_n500), .ZN(new_n505));
  INV_X1    g319(.A(new_n503), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n505), .A2(KEYINPUT20), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n491), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(G234), .A2(G237), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(G952), .A3(new_n214), .ZN(new_n510));
  XOR2_X1   g324(.A(KEYINPUT21), .B(G898), .Z(new_n511));
  NAND3_X1  g325(.A1(new_n509), .A2(G902), .A3(G953), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(KEYINPUT92), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n460), .A2(new_n508), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(G214), .B1(G237), .B2(G902), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n371), .A2(G101), .A3(new_n373), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n350), .A2(KEYINPUT4), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n295), .B(new_n377), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n291), .A2(KEYINPUT5), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT5), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n523), .A2(new_n188), .A3(G116), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G113), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n293), .A2(new_n288), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n356), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n521), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(G110), .B(G122), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n521), .A2(new_n529), .A3(new_n531), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(KEYINPUT6), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT77), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n285), .A2(G125), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n283), .A2(new_n196), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT79), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n214), .A2(G224), .ZN(new_n542));
  XOR2_X1   g356(.A(new_n542), .B(KEYINPUT78), .Z(new_n543));
  INV_X1    g357(.A(KEYINPUT79), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n538), .A2(new_n539), .A3(new_n544), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n541), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n543), .B1(new_n541), .B2(new_n545), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n533), .A2(KEYINPUT77), .A3(KEYINPUT6), .A4(new_n534), .ZN(new_n549));
  OR2_X1    g363(.A1(new_n533), .A2(KEYINPUT6), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n537), .A2(new_n548), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n540), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n543), .A2(KEYINPUT7), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT81), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n543), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  OAI211_X1 g370(.A(KEYINPUT7), .B(new_n543), .C1(new_n540), .C2(new_n554), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n524), .A2(KEYINPUT80), .A3(G113), .ZN(new_n558));
  AOI21_X1  g372(.A(KEYINPUT80), .B1(new_n524), .B2(G113), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n522), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n356), .B1(new_n560), .B2(new_n527), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n528), .A2(new_n362), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n531), .B(KEYINPUT8), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n556), .A2(new_n557), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(G902), .B1(new_n565), .B2(new_n534), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n551), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(G210), .B1(G237), .B2(G902), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n551), .A2(new_n568), .A3(new_n566), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n518), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n334), .A2(new_n411), .A3(new_n516), .A4(new_n572), .ZN(new_n573));
  XOR2_X1   g387(.A(new_n573), .B(new_n346), .Z(G3));
  INV_X1    g388(.A(KEYINPUT33), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n575), .B1(new_n452), .B2(new_n453), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n445), .A2(new_n450), .ZN(new_n577));
  INV_X1    g391(.A(new_n451), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n445), .A2(new_n450), .A3(new_n451), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(KEYINPUT33), .A3(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n455), .A2(G902), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n576), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n229), .B1(new_n452), .B2(new_n453), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n455), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n508), .A2(new_n586), .A3(new_n514), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n551), .A2(new_n568), .A3(new_n566), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n568), .B1(new_n551), .B2(new_n566), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n517), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(KEYINPUT93), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT93), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n592), .B(new_n517), .C1(new_n588), .C2(new_n589), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n587), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n339), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n398), .A2(new_n402), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n596), .A2(new_n338), .A3(new_n229), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n410), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n320), .A2(new_n321), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(G472), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n601), .B1(new_n320), .B2(new_n229), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n600), .A2(new_n602), .A3(new_n238), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n598), .A2(new_n603), .A3(new_n336), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n594), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(KEYINPUT34), .B(G104), .Z(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G6));
  XNOR2_X1  g421(.A(new_n491), .B(KEYINPUT94), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n502), .A2(new_n492), .A3(new_n503), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT20), .B1(new_n505), .B2(new_n506), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n608), .A2(new_n460), .A3(new_n611), .A4(new_n514), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(new_n591), .B2(new_n593), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n604), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT35), .B(G107), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G9));
  OR3_X1    g430(.A1(new_n209), .A2(new_n223), .A3(KEYINPUT36), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n209), .B1(new_n223), .B2(KEYINPUT36), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n617), .A2(new_n236), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT95), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n617), .A2(new_n618), .A3(KEYINPUT95), .A4(new_n236), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n235), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT96), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n235), .A2(new_n621), .A3(KEYINPUT96), .A4(new_n622), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n627), .A2(new_n600), .A3(new_n602), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n411), .A2(new_n572), .A3(new_n516), .A4(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT37), .B(G110), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G12));
  NAND2_X1  g445(.A1(new_n591), .A2(new_n593), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT32), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n599), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n634), .A2(new_n333), .A3(new_n322), .ZN(new_n635));
  INV_X1    g449(.A(new_n627), .ZN(new_n636));
  AND4_X1   g450(.A1(new_n635), .A2(new_n598), .A3(new_n336), .A4(new_n636), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n632), .A2(new_n637), .ZN(new_n638));
  OR2_X1    g452(.A1(new_n512), .A2(G900), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n510), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n608), .A2(new_n460), .A3(new_n611), .A4(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G128), .ZN(G30));
  NOR2_X1   g458(.A1(new_n588), .A2(new_n589), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT97), .ZN(new_n646));
  OR2_X1    g460(.A1(new_n646), .A2(KEYINPUT38), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(KEYINPUT38), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n640), .B(KEYINPUT39), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n411), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT40), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n308), .B1(new_n329), .B2(new_n301), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n296), .A2(new_n301), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n654), .B1(new_n655), .B2(new_n308), .ZN(new_n656));
  OAI21_X1  g470(.A(G472), .B1(new_n656), .B2(G902), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n634), .A2(new_n322), .A3(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n460), .A2(new_n508), .ZN(new_n660));
  NOR4_X1   g474(.A1(new_n659), .A2(new_n660), .A3(new_n518), .A4(new_n623), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n650), .A2(new_n653), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G143), .ZN(G45));
  NAND3_X1  g477(.A1(new_n508), .A2(new_n586), .A3(new_n640), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n638), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G146), .ZN(G48));
  OAI21_X1  g481(.A(KEYINPUT76), .B1(new_n396), .B2(KEYINPUT12), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n391), .A2(new_n392), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n668), .A2(new_n669), .A3(new_n390), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n401), .B1(new_n670), .B2(new_n385), .ZN(new_n671));
  OAI21_X1  g485(.A(G469), .B1(new_n671), .B2(G902), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n672), .A2(new_n597), .A3(new_n336), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(KEYINPUT98), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT98), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n672), .A2(new_n597), .A3(new_n675), .A4(new_n336), .ZN(new_n676));
  AND3_X1   g490(.A1(new_n334), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n594), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT41), .B(G113), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G15));
  NAND2_X1  g494(.A1(new_n677), .A2(new_n613), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G116), .ZN(G18));
  AOI21_X1  g496(.A(new_n673), .B1(new_n591), .B2(new_n593), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n516), .A2(new_n635), .A3(new_n636), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G119), .ZN(G21));
  AOI21_X1  g500(.A(new_n660), .B1(new_n591), .B2(new_n593), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n330), .A2(new_n307), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n310), .A2(new_n688), .A3(new_n319), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n321), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT99), .B(G472), .Z(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(new_n320), .B2(new_n229), .ZN(new_n694));
  NOR4_X1   g508(.A1(new_n691), .A2(new_n694), .A3(new_n238), .A4(new_n515), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n674), .A2(new_n676), .A3(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT100), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n687), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n697), .B1(new_n687), .B2(new_n696), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n412), .ZN(G24));
  AND2_X1   g515(.A1(new_n320), .A2(new_n229), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n623), .B(new_n690), .C1(new_n702), .C2(new_n693), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n664), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n683), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G125), .ZN(G27));
  NAND3_X1  g520(.A1(new_n570), .A2(new_n517), .A3(new_n571), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT101), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT101), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n570), .A2(new_n709), .A3(new_n517), .A4(new_n571), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n708), .A2(new_n411), .A3(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT42), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(KEYINPUT102), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n711), .A2(new_n334), .A3(new_n665), .A4(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n713), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n708), .A2(new_n334), .A3(new_n411), .A4(new_n710), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n715), .B1(new_n716), .B2(new_n664), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G131), .ZN(G33));
  NAND3_X1  g533(.A1(new_n711), .A2(new_n334), .A3(new_n642), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G134), .ZN(G36));
  NAND2_X1  g535(.A1(new_n409), .A2(KEYINPUT45), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n384), .B1(new_n670), .B2(new_n379), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n723), .B1(new_n724), .B2(new_n407), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n722), .A2(new_n725), .A3(G469), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n595), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT46), .ZN(new_n728));
  AOI22_X1  g542(.A1(new_n727), .A2(new_n728), .B1(new_n338), .B2(new_n403), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n726), .A2(KEYINPUT46), .A3(new_n595), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(new_n336), .A3(new_n651), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT103), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n337), .B1(new_n729), .B2(new_n730), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(KEYINPUT103), .A3(new_n651), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT105), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n488), .A2(new_n489), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n493), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n229), .ZN(new_n741));
  AOI22_X1  g555(.A1(new_n609), .A2(new_n610), .B1(new_n741), .B2(G475), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT104), .ZN(new_n743));
  OR2_X1    g557(.A1(new_n743), .A2(KEYINPUT43), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n742), .A2(new_n586), .A3(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  XOR2_X1   g560(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n748), .B1(new_n742), .B2(new_n586), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n738), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n742), .A2(new_n586), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n745), .B(KEYINPUT105), .C1(new_n751), .C2(new_n748), .ZN(new_n752));
  INV_X1    g566(.A(new_n623), .ZN(new_n753));
  INV_X1    g567(.A(new_n602), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n753), .B1(new_n754), .B2(new_n599), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n750), .A2(new_n752), .A3(KEYINPUT44), .A4(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT106), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n708), .A2(new_n710), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n757), .B1(new_n756), .B2(new_n758), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n750), .A2(new_n752), .A3(new_n755), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n763), .A2(KEYINPUT44), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n737), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(new_n210), .ZN(G39));
  INV_X1    g580(.A(new_n238), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n635), .A2(new_n664), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n758), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n731), .A2(new_n336), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT107), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT107), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n735), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n771), .A2(KEYINPUT47), .A3(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT47), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n735), .A2(new_n772), .ZN(new_n776));
  AOI211_X1 g590(.A(KEYINPUT107), .B(new_n337), .C1(new_n729), .C2(new_n730), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n769), .B1(new_n774), .B2(new_n778), .ZN(new_n779));
  XOR2_X1   g593(.A(new_n779), .B(G140), .Z(G42));
  NAND4_X1  g594(.A1(new_n751), .A2(new_n767), .A3(new_n336), .A4(new_n517), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n672), .A2(new_n597), .ZN(new_n782));
  AOI211_X1 g596(.A(new_n658), .B(new_n781), .C1(KEYINPUT49), .C2(new_n782), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n649), .B(new_n783), .C1(KEYINPUT49), .C2(new_n782), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n454), .B(new_n458), .ZN(new_n785));
  AND4_X1   g599(.A1(new_n785), .A2(new_n608), .A3(new_n611), .A4(new_n640), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n708), .A3(new_n710), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(KEYINPUT110), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT110), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n786), .A2(new_n708), .A3(new_n789), .A4(new_n710), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n788), .A2(new_n637), .A3(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n708), .A2(new_n704), .A3(new_n411), .A4(new_n710), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n792), .B1(new_n716), .B2(new_n641), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n718), .A2(new_n791), .A3(new_n794), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n632), .B(new_n637), .C1(new_n642), .C2(new_n665), .ZN(new_n796));
  INV_X1    g610(.A(new_n660), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n640), .B(KEYINPUT111), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n658), .A2(new_n753), .A3(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n632), .A2(new_n411), .A3(new_n797), .A4(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n796), .A2(new_n705), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n796), .A2(new_n705), .A3(new_n800), .A4(KEYINPUT52), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n785), .A2(new_n508), .A3(new_n515), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n411), .A2(new_n572), .A3(new_n806), .A4(new_n603), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n629), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n678), .A2(new_n681), .A3(new_n808), .A4(new_n685), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n700), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(KEYINPUT108), .B1(new_n590), .B2(new_n587), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT108), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n508), .A2(new_n514), .A3(new_n586), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n572), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n604), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n573), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT109), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT109), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n815), .A2(new_n818), .A3(new_n573), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n795), .A2(new_n805), .A3(new_n810), .A4(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n801), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT52), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n801), .A2(new_n824), .A3(new_n802), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n817), .A2(new_n819), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n829), .A2(new_n700), .A3(new_n809), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n828), .A2(KEYINPUT53), .A3(new_n830), .A4(new_n795), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n823), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n794), .A2(new_n791), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n810), .A2(new_n718), .A3(new_n820), .A4(new_n834), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n801), .A2(new_n824), .A3(new_n802), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n802), .B1(new_n801), .B2(new_n824), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n822), .B1(new_n835), .B2(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n830), .A2(KEYINPUT53), .A3(new_n795), .A4(new_n805), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n832), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT113), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n833), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI211_X1 g657(.A(KEYINPUT113), .B(new_n832), .C1(new_n839), .C2(new_n840), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT114), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n718), .A2(new_n791), .A3(new_n794), .ZN(new_n846));
  NOR4_X1   g660(.A1(new_n846), .A2(new_n829), .A3(new_n700), .A4(new_n809), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT53), .B1(new_n847), .B2(new_n828), .ZN(new_n848));
  INV_X1    g662(.A(new_n840), .ZN(new_n849));
  OAI21_X1  g663(.A(KEYINPUT54), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT113), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n841), .A2(new_n842), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n851), .A2(new_n852), .A3(new_n853), .A4(new_n833), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n749), .B1(new_n751), .B2(new_n744), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n855), .A2(new_n510), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n767), .B(new_n690), .C1(new_n702), .C2(new_n693), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n860), .A2(new_n758), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n774), .A2(new_n778), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT115), .ZN(new_n863));
  OAI22_X1  g677(.A1(new_n862), .A2(new_n863), .B1(new_n336), .B2(new_n782), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT115), .B1(new_n774), .B2(new_n778), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n861), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT50), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n673), .A2(new_n517), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n860), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n867), .B1(new_n650), .B2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n649), .A2(KEYINPUT50), .A3(new_n860), .A4(new_n868), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n673), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n758), .A2(new_n873), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n658), .A2(new_n238), .A3(new_n510), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OR2_X1    g690(.A1(new_n876), .A2(KEYINPUT116), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(KEYINPUT116), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n508), .A2(new_n586), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n874), .A2(new_n856), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n881), .A2(new_n703), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n872), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT51), .B1(new_n866), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n782), .A2(new_n336), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n861), .B1(new_n862), .B2(new_n885), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n883), .A2(KEYINPUT51), .A3(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n508), .A2(new_n586), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n877), .A2(new_n888), .A3(new_n878), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n874), .A2(new_n334), .A3(new_n856), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT48), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n214), .A2(G952), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(new_n860), .B2(new_n683), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n889), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n884), .A2(new_n887), .A3(new_n894), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n845), .A2(new_n854), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(G952), .A2(G953), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n784), .B1(new_n896), .B2(new_n897), .ZN(G75));
  INV_X1    g712(.A(KEYINPUT118), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n229), .B1(new_n823), .B2(new_n831), .ZN(new_n900));
  AOI211_X1 g714(.A(new_n899), .B(KEYINPUT56), .C1(new_n900), .C2(G210), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n537), .A2(new_n549), .A3(new_n550), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(new_n548), .Z(new_n903));
  XNOR2_X1  g717(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n903), .B(new_n904), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n901), .A2(new_n905), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n214), .A2(G952), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(G51));
  NAND2_X1  g723(.A1(new_n823), .A2(new_n831), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT54), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n833), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n339), .B(KEYINPUT57), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n596), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n900), .A2(G469), .A3(new_n722), .A4(new_n725), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n908), .B1(new_n915), .B2(new_n916), .ZN(G54));
  NAND3_X1  g731(.A1(new_n900), .A2(KEYINPUT58), .A3(G475), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n918), .A2(new_n505), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n919), .A2(KEYINPUT119), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(KEYINPUT119), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n908), .B1(new_n918), .B2(new_n505), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(G60));
  NAND2_X1  g737(.A1(G478), .A2(G902), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT59), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n912), .A2(new_n576), .A3(new_n581), .A4(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(G952), .B2(new_n214), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n823), .A2(new_n832), .A3(new_n831), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n928), .B1(new_n850), .B2(KEYINPUT113), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n852), .B1(new_n929), .B2(new_n853), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n843), .A2(KEYINPUT114), .A3(new_n844), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n925), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n576), .A2(new_n581), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n927), .B1(new_n932), .B2(new_n933), .ZN(G63));
  XNOR2_X1  g748(.A(new_n231), .B(KEYINPUT120), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT60), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n910), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n908), .B1(new_n937), .B2(new_n226), .ZN(new_n938));
  INV_X1    g752(.A(new_n937), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT121), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n617), .A2(new_n618), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n940), .B1(new_n939), .B2(new_n941), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n938), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI211_X1 g760(.A(KEYINPUT61), .B(new_n938), .C1(new_n942), .C2(new_n943), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(G66));
  NAND3_X1  g762(.A1(new_n511), .A2(G224), .A3(G953), .ZN(new_n949));
  INV_X1    g763(.A(new_n830), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n949), .B1(new_n950), .B2(G953), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n902), .B1(G898), .B2(new_n214), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n951), .B(new_n952), .Z(G69));
  NOR2_X1   g767(.A1(new_n214), .A2(G900), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n954), .B1(new_n381), .B2(G953), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT124), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n281), .A2(new_n287), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT122), .Z(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(new_n498), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n961));
  INV_X1    g775(.A(new_n769), .ZN(new_n962));
  INV_X1    g776(.A(new_n737), .ZN(new_n963));
  INV_X1    g777(.A(new_n761), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n764), .B1(new_n964), .B2(new_n759), .ZN(new_n965));
  AOI22_X1  g779(.A1(new_n862), .A2(new_n962), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n734), .A2(new_n334), .A3(new_n687), .A4(new_n736), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n796), .A2(new_n705), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n968), .A2(new_n720), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n967), .A2(new_n718), .A3(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(G953), .B1(new_n966), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n961), .B1(new_n972), .B2(new_n954), .ZN(new_n973));
  INV_X1    g787(.A(new_n954), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n970), .A2(new_n765), .A3(new_n779), .ZN(new_n975));
  OAI211_X1 g789(.A(KEYINPUT125), .B(new_n974), .C1(new_n975), .C2(G953), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n960), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n888), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(new_n785), .B2(new_n508), .ZN(new_n979));
  AND4_X1   g793(.A1(new_n334), .A2(new_n758), .A3(new_n652), .A4(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n662), .A2(new_n968), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT62), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n662), .A2(KEYINPUT62), .A3(new_n968), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n980), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(G953), .B1(new_n985), .B2(new_n966), .ZN(new_n986));
  INV_X1    g800(.A(new_n960), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n957), .B1(new_n977), .B2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT126), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI211_X1 g805(.A(KEYINPUT126), .B(new_n957), .C1(new_n977), .C2(new_n988), .ZN(new_n992));
  INV_X1    g806(.A(new_n977), .ZN(new_n993));
  OR3_X1    g807(.A1(new_n986), .A2(KEYINPUT123), .A3(new_n987), .ZN(new_n994));
  OAI21_X1  g808(.A(KEYINPUT123), .B1(new_n986), .B2(new_n987), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n993), .A2(new_n994), .A3(new_n956), .A4(new_n995), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n991), .A2(new_n992), .A3(new_n996), .ZN(G72));
  NAND2_X1  g811(.A1(G472), .A2(G902), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT63), .Z(new_n999));
  INV_X1    g813(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n1000), .B1(new_n975), .B2(new_n830), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n655), .B(KEYINPUT127), .ZN(new_n1002));
  NOR3_X1   g816(.A1(new_n1001), .A2(new_n308), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n308), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n985), .A2(new_n830), .A3(new_n966), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1004), .B1(new_n1005), .B2(new_n999), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n655), .B(new_n307), .ZN(new_n1007));
  AOI211_X1 g821(.A(new_n1000), .B(new_n1007), .C1(new_n839), .C2(new_n840), .ZN(new_n1008));
  NOR4_X1   g822(.A1(new_n1003), .A2(new_n1006), .A3(new_n908), .A4(new_n1008), .ZN(G57));
endmodule


