//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n614, new_n615, new_n616,
    new_n618, new_n619, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n778, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896;
  INV_X1    g000(.A(G113gat), .ZN(new_n202));
  INV_X1    g001(.A(G120gat), .ZN(new_n203));
  AOI21_X1  g002(.A(KEYINPUT1), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(new_n202), .B2(new_n203), .ZN(new_n205));
  INV_X1    g004(.A(G127gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(G134gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n205), .B1(KEYINPUT72), .B2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G127gat), .B(G134gat), .Z(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G155gat), .ZN(new_n212));
  INV_X1    g011(.A(G162gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n212), .A2(new_n213), .A3(KEYINPUT79), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT79), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n215), .B1(G155gat), .B2(G162gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n214), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G148gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G141gat), .ZN(new_n220));
  INV_X1    g019(.A(G141gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G148gat), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT2), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n212), .A2(new_n213), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n217), .B1(new_n225), .B2(KEYINPUT2), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT80), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n220), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(new_n222), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n220), .A2(new_n227), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n226), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n224), .A2(new_n231), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n232), .A2(KEYINPUT3), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(KEYINPUT3), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n211), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT4), .ZN(new_n236));
  INV_X1    g035(.A(new_n232), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n210), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n235), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n232), .B(KEYINPUT81), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT4), .B1(new_n240), .B2(new_n210), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT5), .ZN(new_n243));
  NAND2_X1  g042(.A1(G225gat), .A2(G233gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n238), .A2(KEYINPUT4), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n236), .B1(new_n240), .B2(new_n210), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT82), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n249), .B1(new_n248), .B2(new_n247), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(new_n244), .A3(new_n235), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n210), .B(new_n237), .ZN(new_n252));
  INV_X1    g051(.A(new_n244), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n252), .A2(KEYINPUT83), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT83), .B1(new_n252), .B2(new_n253), .ZN(new_n255));
  NOR3_X1   g054(.A1(new_n254), .A2(new_n255), .A3(new_n243), .ZN(new_n256));
  AND3_X1   g055(.A1(new_n251), .A2(KEYINPUT84), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT84), .B1(new_n251), .B2(new_n256), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n245), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G1gat), .B(G29gat), .ZN(new_n260));
  INV_X1    g059(.A(G85gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT0), .B(G57gat), .ZN(new_n263));
  XOR2_X1   g062(.A(new_n262), .B(new_n263), .Z(new_n264));
  OR2_X1    g063(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT6), .B1(new_n259), .B2(new_n264), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n259), .A2(KEYINPUT6), .A3(new_n264), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT90), .ZN(new_n269));
  AND2_X1   g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G8gat), .B(G36gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(G64gat), .B(G92gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n275), .B(KEYINPUT66), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT26), .ZN(new_n277));
  INV_X1    g076(.A(G169gat), .ZN(new_n278));
  INV_X1    g077(.A(G176gat), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .A4(KEYINPUT70), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n279), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT26), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n276), .A2(new_n280), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(G183gat), .A2(G190gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  XOR2_X1   g085(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n287));
  INV_X1    g086(.A(KEYINPUT67), .ZN(new_n288));
  INV_X1    g087(.A(G183gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n289), .A2(KEYINPUT27), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT27), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n291), .A2(G183gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n288), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(G183gat), .ZN(new_n294));
  AOI21_X1  g093(.A(G190gat), .B1(new_n294), .B2(KEYINPUT67), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n287), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT27), .B(G183gat), .ZN(new_n297));
  INV_X1    g096(.A(G190gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(KEYINPUT28), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT69), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n289), .A2(KEYINPUT27), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT67), .B1(new_n294), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT67), .B1(new_n289), .B2(KEYINPUT27), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(new_n298), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n302), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT69), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n308), .A3(new_n299), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n286), .B1(new_n301), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n281), .B(KEYINPUT23), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n311), .A2(new_n276), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT24), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n285), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n315), .A2(KEYINPUT65), .ZN(new_n316));
  NAND3_X1  g115(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT65), .ZN(new_n318));
  OAI221_X1 g117(.A(new_n317), .B1(G183gat), .B2(G190gat), .C1(new_n314), .C2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n312), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT25), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n314), .B(new_n317), .C1(G183gat), .C2(G190gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n312), .A2(new_n323), .A3(KEYINPUT25), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n310), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  AND2_X1   g124(.A1(G226gat), .A2(G233gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n322), .A2(new_n324), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n301), .A2(new_n309), .ZN(new_n329));
  INV_X1    g128(.A(new_n286), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT71), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT71), .ZN(new_n332));
  AOI211_X1 g131(.A(new_n332), .B(new_n286), .C1(new_n301), .C2(new_n309), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n328), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n326), .A2(KEYINPUT29), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n327), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G197gat), .B(G204gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT77), .B(KEYINPUT22), .ZN(new_n340));
  INV_X1    g139(.A(G211gat), .ZN(new_n341));
  INV_X1    g140(.A(G218gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n339), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  XOR2_X1   g143(.A(G211gat), .B(G218gat), .Z(new_n345));
  XOR2_X1   g144(.A(new_n344), .B(new_n345), .Z(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  OR2_X1    g146(.A1(new_n338), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n325), .A2(new_n337), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n349), .B1(new_n335), .B2(new_n326), .ZN(new_n350));
  OR2_X1    g149(.A1(new_n350), .A2(new_n346), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT37), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n348), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  OR2_X1    g152(.A1(new_n353), .A2(KEYINPUT89), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(KEYINPUT89), .ZN(new_n355));
  AOI211_X1 g154(.A(KEYINPUT38), .B(new_n274), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  OR2_X1    g155(.A1(new_n350), .A2(new_n347), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n357), .B(KEYINPUT37), .C1(new_n346), .C2(new_n338), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(KEYINPUT88), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n348), .A2(new_n351), .A3(new_n274), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT78), .ZN(new_n361));
  OR2_X1    g160(.A1(new_n360), .A2(KEYINPUT78), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n356), .A2(new_n359), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT90), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n259), .A2(new_n364), .A3(KEYINPUT6), .A4(new_n264), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n354), .A2(new_n355), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n348), .A2(new_n351), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n274), .B1(new_n367), .B2(KEYINPUT37), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT38), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n270), .A2(new_n363), .A3(new_n365), .A4(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G78gat), .B(G106gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n372), .B(G50gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n373), .B(KEYINPUT31), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT29), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n233), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n346), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT3), .B1(new_n347), .B2(new_n376), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n378), .B1(new_n237), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n380), .A2(G228gat), .A3(G233gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(G228gat), .A2(G233gat), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n378), .B(new_n382), .C1(new_n240), .C2(new_n379), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT87), .B1(new_n384), .B2(G22gat), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT86), .ZN(new_n386));
  INV_X1    g185(.A(G22gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n381), .A2(new_n387), .A3(new_n383), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n385), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n386), .B1(new_n385), .B2(new_n388), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n375), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n391), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n393), .A2(new_n389), .A3(new_n374), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n242), .A2(new_n244), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n397), .B(KEYINPUT39), .C1(new_n253), .C2(new_n252), .ZN(new_n398));
  INV_X1    g197(.A(new_n264), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n398), .B(new_n399), .C1(KEYINPUT39), .C2(new_n397), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT40), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n400), .A2(new_n401), .ZN(new_n403));
  AOI211_X1 g202(.A(new_n402), .B(new_n403), .C1(new_n264), .C2(new_n259), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT30), .B1(new_n362), .B2(new_n361), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n367), .A2(new_n273), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT30), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n406), .B1(new_n407), .B2(new_n360), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n395), .B1(new_n404), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT85), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n265), .A2(new_n412), .A3(new_n266), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n259), .B(new_n264), .C1(KEYINPUT85), .C2(KEYINPUT6), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n409), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n371), .A2(new_n411), .B1(new_n416), .B2(new_n395), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n210), .B(new_n328), .C1(new_n331), .C2(new_n333), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT73), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n334), .A2(new_n211), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n307), .A2(new_n308), .A3(new_n299), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n308), .B1(new_n307), .B2(new_n299), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n330), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n332), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n310), .A2(KEYINPUT71), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT73), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n426), .A2(new_n427), .A3(new_n210), .A4(new_n328), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n419), .A2(new_n420), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(G227gat), .A2(G233gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(KEYINPUT64), .ZN(new_n431));
  OR2_X1    g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(KEYINPUT34), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n429), .A2(new_n431), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT33), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XOR2_X1   g235(.A(G15gat), .B(G43gat), .Z(new_n437));
  XNOR2_X1  g236(.A(G71gat), .B(G99gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT74), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT32), .ZN(new_n442));
  AOI211_X1 g241(.A(new_n441), .B(new_n442), .C1(new_n429), .C2(new_n431), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT74), .B1(new_n434), .B2(KEYINPUT32), .ZN(new_n444));
  NOR3_X1   g243(.A1(new_n440), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n439), .A2(KEYINPUT33), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n434), .A2(KEYINPUT32), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT75), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n442), .B1(new_n429), .B2(new_n431), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT75), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(new_n450), .A3(new_n446), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n433), .B1(new_n445), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT76), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n449), .A2(new_n450), .A3(new_n446), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n450), .B1(new_n449), .B2(new_n446), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n434), .A2(KEYINPUT32), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n441), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n449), .A2(KEYINPUT74), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n459), .A2(new_n460), .A3(new_n439), .A4(new_n436), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT34), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n432), .B(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n457), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n453), .A2(new_n454), .A3(new_n464), .ZN(new_n465));
  OAI211_X1 g264(.A(KEYINPUT76), .B(new_n433), .C1(new_n445), .C2(new_n452), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n467), .A2(KEYINPUT36), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n453), .A2(new_n464), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n469), .A2(KEYINPUT36), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n417), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT35), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT91), .ZN(new_n475));
  INV_X1    g274(.A(new_n395), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n475), .B1(new_n467), .B2(new_n476), .ZN(new_n477));
  AOI211_X1 g276(.A(KEYINPUT91), .B(new_n395), .C1(new_n465), .C2(new_n466), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n410), .B1(new_n414), .B2(new_n413), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n474), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n267), .A2(new_n365), .A3(new_n269), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n405), .A2(new_n408), .A3(KEYINPUT35), .ZN(new_n483));
  AND4_X1   g282(.A1(new_n469), .A2(new_n482), .A3(new_n476), .A4(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n473), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G15gat), .B(G22gat), .ZN(new_n486));
  OR2_X1    g285(.A1(new_n486), .A2(G1gat), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT92), .ZN(new_n488));
  AOI21_X1  g287(.A(G8gat), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT16), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n486), .B1(new_n490), .B2(G1gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n489), .B(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(G57gat), .B(G64gat), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  XOR2_X1   g295(.A(G71gat), .B(G78gat), .Z(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT21), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n493), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(KEYINPUT97), .ZN(new_n501));
  XOR2_X1   g300(.A(KEYINPUT95), .B(KEYINPUT21), .Z(new_n502));
  NOR2_X1   g301(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n501), .B(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(G231gat), .A2(G233gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G127gat), .B(G155gat), .ZN(new_n507));
  XOR2_X1   g306(.A(new_n507), .B(KEYINPUT20), .Z(new_n508));
  XOR2_X1   g307(.A(KEYINPUT96), .B(KEYINPUT19), .Z(new_n509));
  XNOR2_X1  g308(.A(G183gat), .B(G211gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n508), .B(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n506), .A2(new_n513), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G43gat), .B(G50gat), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT14), .ZN(new_n518));
  INV_X1    g317(.A(G29gat), .ZN(new_n519));
  INV_X1    g318(.A(G36gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n521), .A2(new_n522), .B1(G29gat), .B2(G36gat), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n523), .A2(KEYINPUT15), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(KEYINPUT15), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n517), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n526), .B1(new_n524), .B2(new_n517), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT17), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(KEYINPUT93), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n527), .A2(KEYINPUT17), .ZN(new_n530));
  NAND2_X1  g329(.A1(G85gat), .A2(G92gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT98), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND2_X1  g332(.A1(G99gat), .A2(G106gat), .ZN(new_n534));
  INV_X1    g333(.A(G92gat), .ZN(new_n535));
  AOI22_X1  g334(.A1(KEYINPUT8), .A2(new_n534), .B1(new_n261), .B2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT99), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  XOR2_X1   g337(.A(G99gat), .B(G106gat), .Z(new_n539));
  OR2_X1    g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n539), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n529), .A2(new_n530), .A3(new_n542), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n527), .ZN(new_n544));
  AND2_X1   g343(.A1(G232gat), .A2(G233gat), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n544), .B1(KEYINPUT41), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G134gat), .B(G162gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n545), .A2(KEYINPUT41), .ZN(new_n550));
  XNOR2_X1  g349(.A(G190gat), .B(G218gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n549), .A2(new_n552), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n516), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n493), .A2(new_n527), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n530), .A2(new_n493), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n557), .B1(new_n529), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G229gat), .A2(G233gat), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT18), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n493), .B(new_n527), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n560), .B(KEYINPUT13), .Z(new_n563));
  AOI21_X1  g362(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n559), .A2(KEYINPUT18), .A3(new_n560), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G113gat), .B(G141gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(G197gat), .ZN(new_n568));
  XOR2_X1   g367(.A(KEYINPUT11), .B(G169gat), .Z(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT12), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n564), .A2(new_n565), .A3(new_n571), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n573), .A2(KEYINPUT94), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT94), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n566), .A2(new_n576), .A3(new_n572), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G120gat), .B(G148gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(G176gat), .B(G204gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n542), .B(new_n498), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT10), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n540), .A2(KEYINPUT10), .A3(new_n498), .A4(new_n541), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G230gat), .A2(G233gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT100), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n582), .ZN(new_n590));
  INV_X1    g389(.A(new_n587), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n581), .B1(new_n589), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n581), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n586), .A2(new_n587), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NOR3_X1   g397(.A1(new_n556), .A2(new_n578), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n485), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n415), .B(KEYINPUT101), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g403(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n605));
  NAND2_X1  g404(.A1(new_n601), .A2(new_n410), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n605), .B1(new_n606), .B2(G8gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT16), .B(G8gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT103), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT42), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  OAI22_X1  g411(.A1(new_n607), .A2(new_n610), .B1(new_n606), .B2(new_n612), .ZN(G1325gat));
  INV_X1    g412(.A(G15gat), .ZN(new_n614));
  NOR3_X1   g413(.A1(new_n600), .A2(new_n614), .A3(new_n472), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n601), .A2(new_n469), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n615), .B1(new_n614), .B2(new_n616), .ZN(G1326gat));
  NOR2_X1   g416(.A1(new_n600), .A2(new_n476), .ZN(new_n618));
  XOR2_X1   g417(.A(KEYINPUT43), .B(G22gat), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(G1327gat));
  INV_X1    g419(.A(new_n473), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT105), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n622), .B1(new_n481), .B2(new_n484), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n467), .A2(new_n476), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT91), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n467), .A2(new_n475), .A3(new_n476), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n625), .A2(new_n626), .A3(new_n480), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT35), .ZN(new_n628));
  INV_X1    g427(.A(new_n484), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n628), .A2(KEYINPUT105), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n621), .B1(new_n623), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT106), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n555), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n553), .A2(KEYINPUT106), .A3(new_n554), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n636), .A2(KEYINPUT44), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(KEYINPUT107), .B1(new_n631), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT105), .B1(new_n628), .B2(new_n629), .ZN(new_n640));
  AOI211_X1 g439(.A(new_n622), .B(new_n484), .C1(new_n627), .C2(KEYINPUT35), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n473), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT107), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n642), .A2(new_n643), .A3(new_n637), .ZN(new_n644));
  INV_X1    g443(.A(new_n555), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n485), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(KEYINPUT44), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n639), .A2(new_n644), .A3(new_n647), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n578), .A2(new_n516), .A3(new_n598), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n649), .B(KEYINPUT104), .Z(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n602), .ZN(new_n652));
  OAI21_X1  g451(.A(G29gat), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n485), .A2(new_n645), .A3(new_n649), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n654), .A2(G29gat), .A3(new_n652), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n655), .B(KEYINPUT45), .Z(new_n656));
  NAND2_X1  g455(.A1(new_n653), .A2(new_n656), .ZN(G1328gat));
  OAI21_X1  g456(.A(G36gat), .B1(new_n651), .B2(new_n409), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n654), .A2(G36gat), .A3(new_n409), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT46), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(G1329gat));
  NAND3_X1  g460(.A1(new_n648), .A2(new_n471), .A3(new_n650), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(G43gat), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(KEYINPUT108), .ZN(new_n664));
  INV_X1    g463(.A(new_n469), .ZN(new_n665));
  OR3_X1    g464(.A1(new_n654), .A2(G43gat), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT47), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n664), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n663), .B(new_n666), .C1(KEYINPUT108), .C2(KEYINPUT47), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(G1330gat));
  OAI21_X1  g470(.A(G50gat), .B1(new_n651), .B2(new_n476), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n654), .A2(G50gat), .A3(new_n476), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT48), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n672), .A2(KEYINPUT48), .A3(new_n674), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(G1331gat));
  NAND2_X1  g478(.A1(new_n578), .A2(new_n598), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n631), .A2(new_n556), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n602), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g482(.A(new_n409), .B(KEYINPUT109), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n685), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT110), .B(KEYINPUT111), .ZN(new_n688));
  NOR2_X1   g487(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n687), .B(new_n690), .ZN(G1333gat));
  AOI21_X1  g490(.A(G71gat), .B1(new_n681), .B2(new_n469), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n471), .A2(G71gat), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n692), .B1(new_n681), .B2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1334gat));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n395), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g497(.A1(new_n680), .A2(new_n516), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n648), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(G85gat), .B1(new_n700), .B2(new_n652), .ZN(new_n701));
  INV_X1    g500(.A(new_n578), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n702), .A2(new_n516), .A3(new_n555), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n642), .A2(KEYINPUT51), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT51), .B1(new_n642), .B2(new_n703), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n602), .A2(new_n261), .A3(new_n598), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n701), .B1(new_n706), .B2(new_n707), .ZN(G1336gat));
  AND2_X1   g507(.A1(new_n648), .A2(new_n699), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n535), .B1(new_n709), .B2(new_n410), .ZN(new_n710));
  INV_X1    g509(.A(new_n598), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n685), .A2(G92gat), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(new_n704), .B2(new_n705), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT113), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT113), .ZN(new_n715));
  OAI211_X1 g514(.A(new_n715), .B(new_n712), .C1(new_n704), .C2(new_n705), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT52), .B1(new_n710), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(G92gat), .B1(new_n700), .B2(new_n685), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT114), .ZN(new_n720));
  AOI21_X1  g519(.A(KEYINPUT52), .B1(new_n713), .B2(new_n720), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n719), .B(new_n721), .C1(new_n720), .C2(new_n713), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n718), .A2(new_n722), .ZN(G1337gat));
  OAI21_X1  g522(.A(G99gat), .B1(new_n700), .B2(new_n472), .ZN(new_n724));
  OR3_X1    g523(.A1(new_n665), .A2(G99gat), .A3(new_n711), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(new_n706), .B2(new_n725), .ZN(G1338gat));
  NAND3_X1  g525(.A1(new_n648), .A2(new_n395), .A3(new_n699), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(G106gat), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT115), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n476), .A2(G106gat), .A3(new_n711), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n704), .B2(new_n705), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n729), .A2(new_n732), .A3(KEYINPUT53), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT53), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n728), .B(new_n731), .C1(KEYINPUT115), .C2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(G1339gat));
  INV_X1    g535(.A(new_n581), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT54), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(new_n589), .B2(new_n738), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n596), .B(KEYINPUT54), .C1(new_n586), .C2(new_n588), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT55), .ZN(new_n742));
  AOI22_X1  g541(.A1(new_n741), .A2(new_n742), .B1(new_n596), .B2(new_n595), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n739), .A2(KEYINPUT55), .A3(new_n740), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n743), .A2(new_n577), .A3(new_n575), .A4(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n559), .A2(new_n560), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n562), .A2(new_n563), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n570), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n574), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n598), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n635), .B1(new_n745), .B2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n743), .A2(new_n744), .A3(new_n749), .ZN(new_n753));
  OR2_X1    g552(.A1(new_n636), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n752), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n516), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n636), .A2(new_n753), .ZN(new_n758));
  OAI21_X1  g557(.A(KEYINPUT116), .B1(new_n758), .B2(new_n751), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n756), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n578), .A2(new_n516), .A3(new_n555), .A4(new_n711), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT117), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n760), .A2(KEYINPUT117), .A3(new_n761), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n766), .A2(new_n652), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n479), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n768), .A2(new_n684), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n769), .A2(new_n202), .A3(new_n702), .ZN(new_n770));
  AND4_X1   g569(.A1(new_n602), .A2(new_n764), .A3(new_n685), .A4(new_n765), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n771), .A2(new_n469), .A3(new_n476), .ZN(new_n772));
  OAI21_X1  g571(.A(G113gat), .B1(new_n772), .B2(new_n578), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n770), .A2(new_n773), .ZN(G1340gat));
  NAND3_X1  g573(.A1(new_n769), .A2(new_n203), .A3(new_n598), .ZN(new_n775));
  OAI21_X1  g574(.A(G120gat), .B1(new_n772), .B2(new_n711), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(G1341gat));
  NOR3_X1   g576(.A1(new_n772), .A2(new_n206), .A3(new_n757), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n769), .A2(new_n516), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n778), .B1(new_n779), .B2(new_n206), .ZN(G1342gat));
  OAI21_X1  g579(.A(G134gat), .B1(new_n772), .B2(new_n555), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT118), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n410), .A2(new_n555), .ZN(new_n785));
  INV_X1    g584(.A(G134gat), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT56), .B1(new_n768), .B2(new_n787), .ZN(new_n788));
  OR3_X1    g587(.A1(new_n768), .A2(KEYINPUT56), .A3(new_n787), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n783), .A2(new_n784), .A3(new_n788), .A4(new_n789), .ZN(G1343gat));
  INV_X1    g589(.A(KEYINPUT57), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n764), .A2(new_n791), .A3(new_n395), .A4(new_n765), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n472), .A2(new_n602), .A3(new_n685), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n645), .B1(new_n745), .B2(new_n750), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n757), .B1(new_n758), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n761), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n395), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n793), .B1(new_n797), .B2(KEYINPUT57), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n792), .A2(new_n702), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(G141gat), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n471), .A2(new_n476), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(KEYINPUT119), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n771), .A2(new_n221), .A3(new_n702), .A4(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT121), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n800), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n804), .B1(new_n800), .B2(new_n803), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT58), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT120), .B1(new_n799), .B2(G141gat), .ZN(new_n808));
  OAI22_X1  g607(.A1(new_n805), .A2(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n800), .A2(new_n803), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT121), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT120), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n807), .B1(new_n800), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n800), .A2(new_n803), .A3(new_n804), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n811), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n809), .A2(new_n815), .ZN(G1344gat));
  AND2_X1   g615(.A1(new_n771), .A2(new_n802), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(new_n219), .A3(new_n598), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT59), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n753), .A2(new_n555), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n757), .B1(new_n794), .B2(new_n820), .ZN(new_n821));
  AOI211_X1 g620(.A(KEYINPUT57), .B(new_n476), .C1(new_n821), .C2(new_n761), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n764), .A2(new_n395), .A3(new_n765), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n822), .B1(new_n823), .B2(KEYINPUT57), .ZN(new_n824));
  INV_X1    g623(.A(new_n793), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n824), .A2(new_n598), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n819), .B1(new_n826), .B2(G148gat), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n792), .A2(new_n798), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(new_n711), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n829), .A2(KEYINPUT59), .A3(new_n219), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n818), .B1(new_n827), .B2(new_n830), .ZN(G1345gat));
  AOI21_X1  g630(.A(G155gat), .B1(new_n817), .B2(new_n516), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n828), .A2(new_n212), .A3(new_n757), .ZN(new_n833));
  OR3_X1    g632(.A1(new_n832), .A2(KEYINPUT122), .A3(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT122), .B1(new_n832), .B2(new_n833), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(G1346gat));
  OAI21_X1  g635(.A(G162gat), .B1(new_n828), .B2(new_n636), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n767), .A2(new_n213), .A3(new_n785), .A4(new_n802), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1347gat));
  NOR3_X1   g638(.A1(new_n665), .A2(new_n395), .A3(new_n409), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n764), .A2(new_n652), .A3(new_n765), .A4(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(G169gat), .B1(new_n841), .B2(new_n578), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n766), .A2(new_n602), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n685), .A2(new_n477), .A3(new_n478), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n702), .A2(new_n278), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n842), .B1(new_n845), .B2(new_n846), .ZN(G1348gat));
  NOR3_X1   g646(.A1(new_n841), .A2(new_n279), .A3(new_n711), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n843), .A2(new_n598), .A3(new_n844), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n848), .B1(new_n849), .B2(new_n279), .ZN(G1349gat));
  NAND4_X1  g649(.A1(new_n843), .A2(new_n297), .A3(new_n516), .A4(new_n844), .ZN(new_n851));
  OAI21_X1  g650(.A(G183gat), .B1(new_n841), .B2(new_n757), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT60), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n854), .A2(KEYINPUT124), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n854), .A2(KEYINPUT124), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT123), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n851), .A2(new_n852), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n857), .B1(new_n858), .B2(KEYINPUT60), .ZN(new_n859));
  AOI211_X1 g658(.A(KEYINPUT123), .B(new_n853), .C1(new_n851), .C2(new_n852), .ZN(new_n860));
  OAI22_X1  g659(.A1(new_n855), .A2(new_n856), .B1(new_n859), .B2(new_n860), .ZN(G1350gat));
  OR2_X1    g660(.A1(new_n841), .A2(new_n555), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT61), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n863), .A3(G190gat), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n863), .B1(new_n862), .B2(G190gat), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n635), .A2(new_n298), .ZN(new_n867));
  OAI22_X1  g666(.A1(new_n865), .A2(new_n866), .B1(new_n845), .B2(new_n867), .ZN(G1351gat));
  NAND2_X1  g667(.A1(new_n801), .A2(new_n684), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT125), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n869), .A2(KEYINPUT125), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n843), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(G197gat), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n872), .A2(new_n873), .A3(new_n702), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n471), .A2(new_n602), .A3(new_n409), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n824), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(G197gat), .B1(new_n876), .B2(new_n578), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT126), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT126), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n874), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(G1352gat));
  NAND3_X1  g681(.A1(new_n824), .A2(new_n598), .A3(new_n875), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(G204gat), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n711), .A2(G204gat), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n843), .A2(new_n870), .A3(new_n871), .A4(new_n885), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n886), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n887));
  AOI21_X1  g686(.A(KEYINPUT127), .B1(new_n886), .B2(KEYINPUT62), .ZN(new_n888));
  OAI221_X1 g687(.A(new_n884), .B1(KEYINPUT62), .B2(new_n886), .C1(new_n887), .C2(new_n888), .ZN(G1353gat));
  NAND3_X1  g688(.A1(new_n872), .A2(new_n341), .A3(new_n516), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n824), .A2(new_n516), .A3(new_n875), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n891), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT63), .B1(new_n891), .B2(G211gat), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n890), .B1(new_n892), .B2(new_n893), .ZN(G1354gat));
  AOI21_X1  g693(.A(G218gat), .B1(new_n872), .B2(new_n635), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n876), .A2(new_n342), .A3(new_n555), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n895), .A2(new_n896), .ZN(G1355gat));
endmodule


