//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 1 1 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1238, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT65), .Z(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(new_n201), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT1), .ZN(new_n220));
  INV_X1    g0020(.A(new_n209), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI21_X1  g0023(.A(KEYINPUT66), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n222), .A2(new_n223), .A3(KEYINPUT66), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n221), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n212), .B(new_n219), .C1(new_n220), .C2(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n230), .A2(new_n220), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT67), .Z(new_n233));
  NOR2_X1   g0033(.A1(new_n231), .A2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  AND2_X1   g0050(.A1(new_n250), .A2(new_n216), .ZN(new_n251));
  INV_X1    g0051(.A(G13), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G1), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G20), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT71), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NOR3_X1   g0057(.A1(new_n252), .A2(new_n217), .A3(G1), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n250), .A2(new_n216), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT71), .ZN(new_n261));
  INV_X1    g0061(.A(G1), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n257), .A2(new_n261), .B1(new_n262), .B2(G20), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G50), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n203), .A2(G20), .ZN(new_n265));
  INV_X1    g0065(.A(G150), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G20), .A2(G33), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n217), .A2(G33), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT8), .B(G58), .ZN(new_n270));
  OAI221_X1 g0070(.A(new_n265), .B1(new_n266), .B2(new_n268), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n271), .A2(new_n259), .B1(new_n202), .B2(new_n258), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n264), .A2(KEYINPUT9), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT74), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n273), .B(new_n274), .ZN(new_n275));
  AND2_X1   g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  OAI21_X1  g0076(.A(KEYINPUT69), .B1(new_n276), .B2(new_n216), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT68), .ZN(new_n278));
  INV_X1    g0078(.A(G41), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G45), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT68), .A2(G41), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  AND2_X1   g0083(.A1(G1), .A2(G13), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT69), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G41), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n262), .A2(G274), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n277), .A2(new_n283), .A3(new_n287), .A4(new_n289), .ZN(new_n290));
  NOR3_X1   g0090(.A1(new_n276), .A2(KEYINPUT69), .A3(new_n216), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n285), .B1(new_n284), .B2(new_n286), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n262), .B1(G41), .B2(G45), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(G226), .A3(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(KEYINPUT3), .B(G33), .ZN(new_n296));
  INV_X1    g0096(.A(G1698), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G222), .ZN(new_n299));
  INV_X1    g0099(.A(G77), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n298), .A2(new_n299), .B1(new_n300), .B2(new_n296), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT3), .ZN(new_n302));
  INV_X1    g0102(.A(G33), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(KEYINPUT3), .A2(G33), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n297), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT70), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n301), .B1(new_n307), .B2(G223), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n276), .A2(new_n216), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n290), .B(new_n295), .C1(new_n308), .C2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G190), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n264), .A2(new_n272), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT9), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n311), .A2(G200), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n275), .A2(new_n313), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT10), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT10), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n275), .A2(new_n319), .A3(new_n313), .A4(new_n316), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n312), .A2(G169), .ZN(new_n322));
  INV_X1    g0122(.A(new_n314), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n311), .A2(G179), .ZN(new_n324));
  NOR3_X1   g0124(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n321), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n277), .A2(new_n287), .A3(G238), .A4(new_n294), .ZN(new_n328));
  NAND2_X1  g0128(.A1(G33), .A2(G97), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n329), .B(KEYINPUT75), .ZN(new_n330));
  NOR2_X1   g0130(.A1(G226), .A2(G1698), .ZN(new_n331));
  INV_X1    g0131(.A(G232), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n331), .B1(new_n332), .B2(G1698), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n330), .B1(new_n296), .B2(new_n333), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n290), .B(new_n328), .C1(new_n334), .C2(new_n310), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT13), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n333), .A2(new_n296), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n309), .B1(new_n338), .B2(new_n330), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT13), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n339), .A2(new_n340), .A3(new_n290), .A4(new_n328), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n336), .A2(G179), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT77), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT77), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n336), .A2(new_n341), .A3(new_n344), .A4(G179), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G169), .ZN(new_n347));
  AOI211_X1 g0147(.A(KEYINPUT14), .B(new_n347), .C1(new_n336), .C2(new_n341), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n336), .A2(new_n341), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G169), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT14), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n346), .A2(new_n349), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G68), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n258), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT12), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n267), .A2(G50), .B1(G20), .B2(new_n354), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n300), .B2(new_n269), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(KEYINPUT11), .A3(new_n259), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n260), .B(G68), .C1(G1), .C2(new_n217), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n356), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT11), .B1(new_n358), .B2(new_n259), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g0163(.A(new_n363), .B(KEYINPUT78), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n353), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT76), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n336), .A2(G190), .A3(new_n341), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n363), .ZN(new_n369));
  INV_X1    g0169(.A(G200), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n370), .B1(new_n336), .B2(new_n341), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n367), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n371), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n373), .A2(KEYINPUT76), .A3(new_n368), .A4(new_n363), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(G77), .B1(new_n217), .B2(G1), .ZN(new_n376));
  OAI22_X1  g0176(.A1(new_n255), .A2(new_n376), .B1(G77), .B2(new_n254), .ZN(new_n377));
  XNOR2_X1  g0177(.A(KEYINPUT15), .B(G87), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n378), .B(KEYINPUT73), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n303), .A2(G20), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n270), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n382), .A2(new_n267), .B1(G20), .B2(G77), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n377), .B1(new_n384), .B2(new_n259), .ZN(new_n385));
  XNOR2_X1  g0185(.A(KEYINPUT72), .B(G107), .ZN(new_n386));
  OAI22_X1  g0186(.A1(new_n298), .A2(new_n332), .B1(new_n296), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n307), .B2(G238), .ZN(new_n388));
  OR2_X1    g0188(.A1(new_n388), .A2(new_n310), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n293), .A2(G244), .A3(new_n294), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n390), .A2(new_n290), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n385), .B1(new_n392), .B2(new_n347), .ZN(new_n393));
  INV_X1    g0193(.A(G179), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n389), .A2(new_n394), .A3(new_n391), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n370), .B1(new_n389), .B2(new_n391), .ZN(new_n397));
  OAI211_X1 g0197(.A(G190), .B(new_n391), .C1(new_n388), .C2(new_n310), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n385), .ZN(new_n399));
  OR2_X1    g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n366), .A2(new_n375), .A3(new_n396), .A4(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT17), .ZN(new_n402));
  AND2_X1   g0202(.A1(KEYINPUT3), .A2(G33), .ZN(new_n403));
  NOR2_X1   g0203(.A1(KEYINPUT3), .A2(G33), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT7), .B1(new_n405), .B2(new_n217), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n304), .A2(KEYINPUT7), .A3(new_n217), .A4(new_n305), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(G68), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(G58), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n410), .A2(new_n354), .ZN(new_n411));
  OAI21_X1  g0211(.A(G20), .B1(new_n411), .B2(new_n201), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n267), .A2(G159), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n409), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT79), .ZN(new_n417));
  AOI21_X1  g0217(.A(KEYINPUT16), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n304), .A2(new_n217), .A3(new_n305), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT7), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n354), .B1(new_n421), .B2(new_n407), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n417), .B(KEYINPUT16), .C1(new_n422), .C2(new_n414), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n259), .B1(new_n418), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n382), .A2(new_n254), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n426), .B1(new_n263), .B2(new_n382), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n277), .A2(new_n287), .A3(G232), .A4(new_n294), .ZN(new_n429));
  NOR2_X1   g0229(.A1(G223), .A2(G1698), .ZN(new_n430));
  INV_X1    g0230(.A(G226), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n430), .B1(new_n431), .B2(G1698), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n432), .A2(new_n296), .B1(G33), .B2(G87), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n290), .B(new_n429), .C1(new_n433), .C2(new_n310), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n370), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n431), .A2(G1698), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(G223), .B2(G1698), .ZN(new_n437));
  INV_X1    g0237(.A(G87), .ZN(new_n438));
  OAI22_X1  g0238(.A1(new_n437), .A2(new_n405), .B1(new_n303), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n309), .ZN(new_n440));
  INV_X1    g0240(.A(G190), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n440), .A2(new_n441), .A3(new_n290), .A4(new_n429), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n435), .A2(KEYINPUT80), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(KEYINPUT80), .B1(new_n435), .B2(new_n442), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n402), .B1(new_n428), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT18), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n434), .A2(G179), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n448), .B1(new_n347), .B2(new_n434), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n428), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n417), .B1(new_n422), .B2(new_n414), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT16), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n251), .B1(new_n453), .B2(new_n423), .ZN(new_n454));
  INV_X1    g0254(.A(new_n427), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n449), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT18), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n453), .A2(new_n423), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n455), .B1(new_n458), .B2(new_n259), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n435), .A2(new_n442), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT80), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n435), .A2(KEYINPUT80), .A3(new_n442), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n459), .A2(new_n464), .A3(KEYINPUT17), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n446), .A2(new_n450), .A3(new_n457), .A4(new_n465), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n327), .A2(new_n401), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n296), .A2(new_n217), .A3(G87), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT22), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT22), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n296), .A2(new_n470), .A3(new_n217), .A4(G87), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT24), .ZN(new_n473));
  INV_X1    g0273(.A(G107), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G20), .ZN(new_n475));
  INV_X1    g0275(.A(G116), .ZN(new_n476));
  OAI22_X1  g0276(.A1(KEYINPUT23), .A2(new_n475), .B1(new_n269), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n386), .A2(G20), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n477), .B1(new_n478), .B2(KEYINPUT23), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n472), .A2(new_n473), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n473), .B1(new_n472), .B2(new_n479), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n259), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n253), .A2(G20), .A3(new_n474), .ZN(new_n483));
  XNOR2_X1  g0283(.A(new_n483), .B(KEYINPUT25), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n262), .A2(G33), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n251), .A2(new_n254), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n484), .B1(G107), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n482), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(G257), .B(G1698), .C1(new_n403), .C2(new_n404), .ZN(new_n490));
  OAI211_X1 g0290(.A(G250), .B(new_n297), .C1(new_n403), .C2(new_n404), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G33), .A2(G294), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n309), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT5), .ZN(new_n495));
  AND2_X1   g0295(.A1(KEYINPUT68), .A2(G41), .ZN(new_n496));
  NOR2_X1   g0296(.A1(KEYINPUT68), .A2(G41), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n281), .A2(G1), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n279), .A2(KEYINPUT5), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n293), .A2(new_n501), .A3(G264), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n494), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT88), .ZN(new_n504));
  INV_X1    g0304(.A(G274), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n505), .B1(KEYINPUT5), .B2(new_n279), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n277), .A2(new_n287), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(KEYINPUT5), .B1(new_n280), .B2(new_n282), .ZN(new_n508));
  INV_X1    g0308(.A(new_n499), .ZN(new_n509));
  OAI21_X1  g0309(.A(KEYINPUT82), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT82), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n498), .A2(new_n511), .A3(new_n499), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n507), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT88), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n494), .A2(new_n502), .A3(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n504), .A2(G179), .A3(new_n513), .A4(new_n515), .ZN(new_n516));
  OR2_X1    g0316(.A1(new_n516), .A2(KEYINPUT89), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(KEYINPUT89), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n513), .A2(new_n502), .A3(new_n494), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G169), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n494), .A2(new_n502), .A3(new_n514), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n514), .B1(new_n494), .B2(new_n502), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n507), .A2(new_n510), .A3(new_n512), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  OAI22_X1  g0325(.A1(new_n525), .A2(G200), .B1(G190), .B2(new_n519), .ZN(new_n526));
  AND2_X1   g0326(.A1(new_n482), .A2(new_n488), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(new_n527), .A3(KEYINPUT90), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT90), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n519), .A2(G190), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n504), .A2(new_n513), .A3(new_n515), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n530), .B1(new_n531), .B2(new_n370), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n529), .B1(new_n532), .B2(new_n489), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n489), .A2(new_n521), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT21), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n535), .A2(new_n347), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n486), .A2(G116), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n254), .A2(new_n476), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G33), .A2(G283), .ZN(new_n541));
  INV_X1    g0341(.A(G97), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n541), .B(new_n217), .C1(G33), .C2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n476), .A2(G20), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(new_n259), .A3(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT20), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n543), .A2(KEYINPUT20), .A3(new_n259), .A4(new_n544), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n537), .B1(new_n540), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n293), .A2(new_n501), .A3(G270), .ZN(new_n551));
  OAI211_X1 g0351(.A(G264), .B(G1698), .C1(new_n403), .C2(new_n404), .ZN(new_n552));
  OAI211_X1 g0352(.A(G257), .B(new_n297), .C1(new_n403), .C2(new_n404), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n304), .A2(G303), .A3(new_n305), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n309), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n513), .A2(new_n551), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n550), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT87), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT87), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n550), .A2(new_n560), .A3(new_n557), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n540), .A2(new_n549), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n557), .A2(new_n563), .A3(G169), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n394), .B1(new_n555), .B2(new_n309), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n565), .A2(new_n513), .A3(new_n551), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n564), .A2(new_n535), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n563), .B1(new_n557), .B2(G200), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n441), .B2(new_n557), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n562), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n379), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n258), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n379), .A2(new_n487), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n380), .A2(G97), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT19), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n296), .A2(new_n217), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n576), .B1(new_n577), .B2(new_n354), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT85), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n474), .A2(KEYINPUT72), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT72), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G107), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n438), .A2(new_n542), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n579), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n386), .A2(KEYINPUT85), .A3(new_n438), .A4(new_n542), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT75), .ZN(new_n588));
  XNOR2_X1  g0388(.A(new_n329), .B(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n217), .B1(new_n589), .B2(new_n575), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n578), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n572), .B(new_n573), .C1(new_n591), .C2(new_n251), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT86), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n330), .A2(KEYINPUT19), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n595), .A2(new_n217), .B1(new_n585), .B2(new_n586), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n259), .B1(new_n596), .B2(new_n578), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n597), .A2(KEYINPUT86), .A3(new_n572), .A4(new_n573), .ZN(new_n598));
  OAI211_X1 g0398(.A(G238), .B(new_n297), .C1(new_n403), .C2(new_n404), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT84), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT84), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n296), .A2(new_n601), .A3(G238), .A4(new_n297), .ZN(new_n602));
  NAND2_X1  g0402(.A1(G33), .A2(G116), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n296), .A2(G244), .A3(G1698), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n600), .A2(new_n602), .A3(new_n603), .A4(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n309), .ZN(new_n606));
  INV_X1    g0406(.A(G250), .ZN(new_n607));
  OAI22_X1  g0407(.A1(new_n499), .A2(new_n607), .B1(new_n288), .B2(new_n281), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n608), .A2(new_n277), .A3(new_n287), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n606), .A2(G179), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n609), .B1(new_n605), .B2(new_n309), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n611), .B1(new_n347), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n594), .A2(new_n598), .A3(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n612), .A2(new_n370), .ZN(new_n615));
  AOI211_X1 g0415(.A(new_n441), .B(new_n609), .C1(new_n605), .C2(new_n309), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n487), .A2(G87), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n597), .A2(new_n572), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n614), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n293), .A2(new_n501), .A3(G257), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n513), .A2(new_n622), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n306), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n624));
  OAI211_X1 g0424(.A(G244), .B(new_n297), .C1(new_n403), .C2(new_n404), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT4), .ZN(new_n626));
  OAI21_X1  g0426(.A(KEYINPUT81), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(G244), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(new_n304), .B2(new_n305), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT81), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n629), .A2(new_n630), .A3(KEYINPUT4), .A4(new_n297), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n625), .A2(new_n626), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n624), .A2(new_n627), .A3(new_n631), .A4(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n309), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n623), .A2(G190), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n258), .A2(new_n542), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n636), .B1(new_n486), .B2(new_n542), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT6), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n542), .A2(new_n474), .ZN(new_n639));
  NOR2_X1   g0439(.A1(G97), .A2(G107), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n474), .A2(KEYINPUT6), .A3(G97), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n643), .A2(G20), .B1(G77), .B2(new_n267), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n583), .B1(new_n406), .B2(new_n408), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n637), .B1(new_n646), .B2(new_n259), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n635), .A2(new_n647), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n513), .A2(KEYINPUT83), .A3(new_n622), .ZN(new_n649));
  AOI21_X1  g0449(.A(KEYINPUT83), .B1(new_n513), .B2(new_n622), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n634), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(G200), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n623), .A2(new_n634), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n647), .B1(new_n653), .B2(new_n347), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n394), .B(new_n634), .C1(new_n649), .C2(new_n650), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n648), .A2(new_n652), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n570), .A2(new_n621), .A3(new_n656), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n467), .A2(new_n534), .A3(new_n657), .ZN(G372));
  AND2_X1   g0458(.A1(new_n372), .A2(new_n374), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(new_n396), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT14), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(new_n350), .B2(G169), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(new_n348), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n364), .B1(new_n663), .B2(new_n346), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n446), .A2(new_n465), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n457), .B(new_n450), .C1(new_n665), .C2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n325), .B1(new_n667), .B2(new_n321), .ZN(new_n668));
  INV_X1    g0468(.A(new_n467), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n516), .A2(KEYINPUT89), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n520), .B1(new_n516), .B2(KEYINPUT89), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n489), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n560), .B1(new_n550), .B2(new_n557), .ZN(new_n673));
  INV_X1    g0473(.A(new_n561), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n567), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n648), .A2(new_n652), .ZN(new_n678));
  AOI22_X1  g0478(.A1(new_n617), .A2(new_n619), .B1(new_n613), .B2(new_n592), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n653), .A2(new_n347), .ZN(new_n680));
  INV_X1    g0480(.A(new_n647), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(new_n655), .A3(new_n681), .ZN(new_n682));
  AND3_X1   g0482(.A1(new_n678), .A2(new_n679), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n528), .A2(new_n533), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n677), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n613), .A2(new_n592), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n614), .A2(new_n620), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT26), .ZN(new_n689));
  NOR3_X1   g0489(.A1(new_n688), .A2(new_n689), .A3(new_n682), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT91), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n682), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n654), .A2(KEYINPUT91), .A3(new_n655), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(new_n679), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n690), .B1(new_n689), .B2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n687), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n668), .B1(new_n669), .B2(new_n696), .ZN(G369));
  NAND2_X1  g0497(.A1(new_n253), .A2(new_n217), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n698), .A2(KEYINPUT27), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(KEYINPUT27), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(G213), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G343), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n672), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n521), .A2(new_n489), .A3(new_n703), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT92), .ZN(new_n706));
  INV_X1    g0506(.A(new_n703), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n534), .B1(new_n527), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n676), .A2(new_n703), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n704), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n563), .A2(new_n703), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n570), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n676), .B2(new_n712), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n709), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n711), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT93), .ZN(G399));
  INV_X1    g0519(.A(new_n210), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n496), .A2(new_n497), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n587), .A2(G116), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(G1), .A3(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n727), .A2(KEYINPUT94), .B1(new_n215), .B2(new_n723), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(KEYINPUT94), .B2(new_n727), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT28), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n692), .A2(KEYINPUT26), .A3(new_n679), .A4(new_n693), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n689), .B1(new_n688), .B2(new_n682), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n685), .A2(new_n733), .A3(new_n686), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(KEYINPUT29), .A3(new_n707), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n696), .A2(new_n703), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n735), .B1(new_n736), .B2(KEYINPUT29), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT30), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n566), .A2(new_n504), .A3(new_n515), .A4(new_n612), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n738), .B1(new_n739), .B2(new_n653), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n623), .A2(KEYINPUT30), .A3(new_n634), .ZN(new_n741));
  OAI21_X1  g0541(.A(KEYINPUT95), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n623), .A2(KEYINPUT30), .A3(new_n634), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT95), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n522), .A2(new_n523), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n606), .A2(new_n610), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n565), .A2(new_n513), .A3(new_n551), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n743), .A2(new_n744), .A3(new_n745), .A4(new_n748), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n746), .A2(new_n394), .A3(new_n557), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n750), .A2(new_n651), .A3(new_n531), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n740), .A2(new_n742), .A3(new_n749), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(new_n703), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT31), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n752), .A2(KEYINPUT31), .A3(new_n703), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n684), .A2(new_n672), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n570), .A2(new_n621), .A3(new_n656), .A4(new_n707), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n755), .B(new_n756), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G330), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n737), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n730), .B1(new_n762), .B2(G1), .ZN(G364));
  NOR2_X1   g0563(.A1(new_n252), .A2(G20), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n262), .B1(new_n764), .B2(G45), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n724), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n716), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(G330), .B2(new_n714), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n210), .A2(new_n296), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n769), .A2(new_n206), .B1(G116), .B2(new_n210), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n210), .A2(new_n405), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT96), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n214), .A2(G45), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(new_n248), .B2(G45), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n770), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n216), .B1(G20), .B2(new_n347), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT98), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G13), .A2(G33), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT97), .Z(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n766), .B1(new_n775), .B2(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n441), .A2(G179), .A3(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n217), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n542), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n217), .A2(new_n394), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G190), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G200), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n217), .A2(G179), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G190), .A2(G200), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G159), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XOR2_X1   g0596(.A(KEYINPUT99), .B(KEYINPUT32), .Z(new_n797));
  OAI22_X1  g0597(.A1(new_n791), .A2(new_n410), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n789), .A2(new_n370), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n787), .B(new_n798), .C1(G50), .C2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n792), .A2(new_n441), .A3(G200), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G107), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n792), .A2(G190), .A3(G200), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G87), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n803), .A2(new_n806), .A3(new_n296), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT100), .Z(new_n808));
  NAND3_X1  g0608(.A1(new_n788), .A2(new_n441), .A3(G200), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n788), .A2(new_n793), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n809), .A2(new_n354), .B1(new_n810), .B2(new_n300), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(new_n796), .B2(new_n797), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n800), .A2(new_n808), .A3(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(G294), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n786), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n810), .ZN(new_n816));
  INV_X1    g0616(.A(new_n794), .ZN(new_n817));
  AOI22_X1  g0617(.A1(G311), .A2(new_n816), .B1(new_n817), .B2(G329), .ZN(new_n818));
  INV_X1    g0618(.A(G283), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n818), .B1(new_n819), .B2(new_n801), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n815), .B(new_n820), .C1(G326), .C2(new_n799), .ZN(new_n821));
  INV_X1    g0621(.A(G303), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n405), .B1(new_n804), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT101), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n821), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(G322), .ZN(new_n828));
  XOR2_X1   g0628(.A(KEYINPUT33), .B(G317), .Z(new_n829));
  OAI22_X1  g0629(.A1(new_n791), .A2(new_n828), .B1(new_n809), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT102), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n813), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n784), .B1(new_n832), .B2(new_n778), .ZN(new_n833));
  INV_X1    g0633(.A(new_n781), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n833), .B1(new_n714), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n768), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G396));
  AOI21_X1  g0637(.A(KEYINPUT91), .B1(new_n654), .B2(new_n655), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n620), .A2(new_n686), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(KEYINPUT26), .B1(new_n840), .B2(new_n693), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n685), .B(new_n686), .C1(new_n841), .C2(new_n690), .ZN(new_n842));
  AND3_X1   g0642(.A1(new_n396), .A2(new_n400), .A3(new_n707), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n397), .A2(new_n399), .B1(new_n385), .B2(new_n707), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n396), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n393), .A2(new_n395), .A3(new_n707), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n844), .B1(new_n736), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n766), .B1(new_n850), .B2(new_n760), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n760), .B2(new_n850), .ZN(new_n852));
  INV_X1    g0652(.A(new_n780), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n778), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n766), .B1(G77), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n801), .A2(new_n354), .ZN(new_n858));
  INV_X1    g0658(.A(G132), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n296), .B1(new_n794), .B2(new_n859), .C1(new_n202), .C2(new_n804), .ZN(new_n860));
  INV_X1    g0660(.A(new_n786), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n858), .B(new_n860), .C1(G58), .C2(new_n861), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT105), .ZN(new_n863));
  INV_X1    g0663(.A(new_n809), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n864), .A2(G150), .B1(new_n816), .B2(G159), .ZN(new_n865));
  XOR2_X1   g0665(.A(KEYINPUT104), .B(G143), .Z(new_n866));
  INV_X1    g0666(.A(G137), .ZN(new_n867));
  INV_X1    g0667(.A(new_n799), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n865), .B1(new_n791), .B2(new_n866), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n869), .B(KEYINPUT34), .ZN(new_n870));
  OAI22_X1  g0670(.A1(new_n791), .A2(new_n814), .B1(new_n868), .B2(new_n822), .ZN(new_n871));
  OAI22_X1  g0671(.A1(new_n438), .A2(new_n801), .B1(new_n804), .B2(new_n474), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n296), .B(new_n787), .C1(G311), .C2(new_n817), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n809), .A2(new_n819), .B1(new_n810), .B2(new_n476), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT103), .ZN(new_n876));
  OR2_X1    g0676(.A1(new_n875), .A2(KEYINPUT103), .ZN(new_n877));
  AND3_X1   g0677(.A1(new_n874), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n863), .A2(new_n870), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  OAI221_X1 g0679(.A(new_n857), .B1(new_n777), .B2(new_n879), .C1(new_n849), .C2(new_n780), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n852), .A2(new_n880), .ZN(G384));
  NOR2_X1   g0681(.A1(new_n764), .A2(new_n262), .ZN(new_n882));
  INV_X1    g0682(.A(new_n701), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n454), .B2(new_n455), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n466), .A2(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n425), .B(new_n427), .C1(new_n444), .C2(new_n443), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n887), .A2(new_n456), .A3(new_n884), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT37), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT37), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n887), .A2(new_n890), .A3(new_n456), .A4(new_n884), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n886), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(KEYINPUT38), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n886), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n894), .A2(KEYINPUT39), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT107), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT108), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n886), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n893), .A2(new_n900), .A3(new_n895), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT39), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n886), .B(new_n892), .C1(new_n899), .C2(KEYINPUT38), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT107), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n894), .A2(new_n905), .A3(KEYINPUT39), .A4(new_n896), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n898), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n366), .A2(new_n703), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n883), .B1(new_n450), .B2(new_n457), .ZN(new_n910));
  INV_X1    g0710(.A(new_n847), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n842), .B2(new_n843), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n364), .A2(new_n707), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n659), .B2(new_n664), .ZN(new_n914));
  INV_X1    g0714(.A(new_n913), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n366), .A2(new_n375), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n912), .A2(new_n918), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n894), .A2(new_n896), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n910), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n909), .A2(new_n921), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n467), .B(new_n735), .C1(new_n736), .C2(KEYINPUT29), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n668), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n922), .B(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n901), .A2(new_n903), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n848), .B1(new_n914), .B2(new_n916), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n927), .A2(new_n759), .A3(KEYINPUT40), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n894), .A2(new_n927), .A3(new_n759), .A4(new_n896), .ZN(new_n929));
  XNOR2_X1  g0729(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n926), .A2(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n467), .A2(new_n759), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  INV_X1    g0734(.A(G330), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n882), .B1(new_n925), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n925), .B2(new_n937), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n643), .A2(KEYINPUT35), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n643), .A2(KEYINPUT35), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n940), .A2(G116), .A3(new_n218), .A4(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT36), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n214), .A2(new_n300), .A3(new_n411), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT106), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n944), .A2(new_n945), .B1(new_n202), .B2(G68), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n945), .B2(new_n944), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n947), .A2(G1), .A3(new_n252), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n939), .A2(new_n943), .A3(new_n948), .ZN(G367));
  NOR2_X1   g0749(.A1(new_n619), .A2(new_n707), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n950), .A2(new_n592), .A3(new_n613), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n839), .B2(new_n950), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n709), .A2(new_n710), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n656), .B1(new_n647), .B2(new_n707), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n654), .A2(new_n655), .A3(new_n703), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(KEYINPUT42), .B1(new_n954), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n682), .B1(new_n955), .B2(new_n672), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n707), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n954), .A2(KEYINPUT42), .A3(new_n958), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n953), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n965), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n967), .B(new_n953), .C1(new_n962), .C2(new_n963), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n717), .A2(new_n958), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n969), .B(new_n970), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n723), .B(KEYINPUT41), .Z(new_n972));
  INV_X1    g0772(.A(KEYINPUT45), .ZN(new_n973));
  INV_X1    g0773(.A(new_n711), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n973), .B1(new_n974), .B2(new_n958), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n711), .A2(KEYINPUT45), .A3(new_n957), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n974), .A2(KEYINPUT44), .A3(new_n958), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT44), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n711), .B2(new_n957), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n717), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n710), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n709), .B(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(new_n716), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n987), .A2(new_n761), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n977), .A2(new_n717), .A3(new_n981), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n984), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n972), .B1(new_n990), .B2(new_n762), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n765), .B(KEYINPUT110), .Z(new_n992));
  OAI21_X1  g0792(.A(new_n971), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n772), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n994), .A2(new_n241), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n782), .B1(new_n210), .B2(new_n571), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n766), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n868), .A2(new_n866), .B1(new_n804), .B2(new_n410), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n810), .A2(new_n202), .B1(new_n794), .B2(new_n867), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n405), .B(new_n999), .C1(G159), .C2(new_n864), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n354), .B2(new_n786), .C1(new_n300), .C2(new_n801), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n998), .B(new_n1001), .C1(G150), .C2(new_n790), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1002), .A2(KEYINPUT111), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(KEYINPUT111), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n801), .A2(new_n542), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n791), .A2(new_n822), .B1(new_n386), .B2(new_n786), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(G311), .C2(new_n799), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n405), .B1(new_n810), .B2(new_n819), .ZN(new_n1008));
  INV_X1    g0808(.A(G317), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n809), .A2(new_n814), .B1(new_n794), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n804), .A2(new_n476), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n1008), .B(new_n1010), .C1(KEYINPUT46), .C2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1007), .B(new_n1012), .C1(KEYINPUT46), .C2(new_n1011), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1003), .A2(new_n1004), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT47), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1016), .A2(new_n777), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n997), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n834), .B2(new_n952), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n993), .A2(new_n1020), .ZN(G387));
  INV_X1    g0821(.A(new_n987), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n706), .A2(new_n708), .A3(new_n781), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n772), .B1(new_n281), .B2(new_n238), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n725), .B2(new_n769), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n281), .B1(new_n354), .B2(new_n300), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n382), .A2(new_n202), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1026), .B1(new_n1027), .B2(KEYINPUT50), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n725), .B(new_n1028), .C1(KEYINPUT50), .C2(new_n1027), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n1025), .A2(new_n1029), .B1(new_n474), .B2(new_n720), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n766), .B1(new_n1030), .B2(new_n783), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n810), .A2(new_n354), .B1(new_n794), .B2(new_n266), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n405), .B(new_n1032), .C1(new_n382), .C2(new_n864), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1005), .B1(G50), .B2(new_n790), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n804), .A2(new_n300), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(G159), .B2(new_n799), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n379), .A2(new_n861), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1033), .A2(new_n1034), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n861), .A2(G283), .B1(new_n805), .B2(G294), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n864), .A2(G311), .B1(new_n816), .B2(G303), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n791), .B2(new_n1009), .C1(new_n828), .C2(new_n868), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT48), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1039), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT112), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1044), .A2(KEYINPUT49), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n296), .B1(new_n817), .B2(G326), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1046), .B(new_n1047), .C1(new_n476), .C2(new_n801), .ZN(new_n1048));
  AOI21_X1  g0848(.A(KEYINPUT49), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1038), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1031), .B1(new_n1050), .B2(new_n778), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1022), .A2(new_n992), .B1(new_n1023), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n723), .B1(new_n987), .B2(new_n761), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1022), .A2(new_n762), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(G393));
  INV_X1    g0855(.A(new_n989), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n717), .B1(new_n977), .B2(new_n981), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n1056), .A2(new_n1057), .B1(new_n761), .B2(new_n987), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1058), .A2(new_n723), .A3(new_n990), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n772), .A2(new_n245), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n782), .B1(new_n542), .B2(new_n210), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n790), .A2(G311), .B1(new_n799), .B2(G317), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT52), .Z(new_n1063));
  OAI221_X1 g0863(.A(new_n803), .B1(new_n819), .B2(new_n804), .C1(new_n476), .C2(new_n786), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n405), .B1(new_n809), .B2(new_n822), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n810), .A2(new_n814), .B1(new_n794), .B2(new_n828), .ZN(new_n1066));
  NOR3_X1   g0866(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n790), .A2(G159), .B1(new_n799), .B2(G150), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT51), .Z(new_n1069));
  NAND2_X1  g0869(.A1(new_n861), .A2(G77), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1070), .B1(new_n354), .B2(new_n804), .C1(new_n438), .C2(new_n801), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n296), .B1(new_n809), .B2(new_n202), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n866), .A2(new_n794), .B1(new_n810), .B2(new_n270), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n1063), .A2(new_n1067), .B1(new_n1069), .B2(new_n1074), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n766), .B1(new_n1060), .B2(new_n1061), .C1(new_n1075), .C2(new_n777), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n958), .B2(new_n781), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1077), .B1(new_n1078), .B2(new_n992), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1059), .A2(new_n1079), .ZN(G390));
  AND3_X1   g0880(.A1(new_n752), .A2(KEYINPUT31), .A3(new_n703), .ZN(new_n1081));
  AOI21_X1  g0881(.A(KEYINPUT31), .B1(new_n752), .B2(new_n703), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n657), .A2(new_n534), .A3(new_n707), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n935), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n467), .A2(new_n1085), .ZN(new_n1086));
  AND3_X1   g0886(.A1(new_n923), .A2(new_n668), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n844), .A2(new_n847), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n917), .B1(new_n1085), .B2(new_n849), .ZN(new_n1089));
  AND4_X1   g0889(.A1(G330), .A2(new_n759), .A3(new_n849), .A4(new_n917), .ZN(new_n1090));
  OAI211_X1 g0890(.A(KEYINPUT113), .B(new_n1088), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n918), .B1(new_n760), .B2(new_n848), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n734), .A2(new_n707), .A3(new_n846), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1093), .A2(new_n847), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1085), .A2(new_n849), .A3(new_n917), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1092), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1091), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1098));
  AOI21_X1  g0898(.A(KEYINPUT113), .B1(new_n1098), .B2(new_n1088), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1087), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n908), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n912), .B2(new_n918), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1102), .A2(new_n898), .A3(new_n904), .A4(new_n906), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n908), .B1(new_n901), .B2(new_n903), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n1094), .B2(new_n918), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1095), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n1103), .A2(new_n1105), .A3(new_n1095), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1100), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n908), .B1(new_n1088), .B2(new_n917), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1105), .B1(new_n907), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n1090), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT113), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1114), .A2(new_n1096), .A3(new_n1091), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1103), .A2(new_n1105), .A3(new_n1095), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1111), .A2(new_n1115), .A3(new_n1116), .A4(new_n1087), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1108), .A2(new_n1117), .A3(new_n723), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1107), .A2(new_n1106), .ZN(new_n1119));
  OR2_X1    g0919(.A1(new_n907), .A2(new_n780), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n766), .B1(new_n382), .B2(new_n855), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT114), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n861), .A2(G159), .B1(new_n802), .B2(G50), .ZN(new_n1123));
  INV_X1    g0923(.A(G128), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n1123), .B1(new_n1124), .B2(new_n868), .C1(new_n859), .C2(new_n791), .ZN(new_n1125));
  XOR2_X1   g0925(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n1126));
  OR3_X1    g0926(.A1(new_n1126), .A2(new_n804), .A3(new_n266), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT54), .B(G143), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n816), .A2(new_n1129), .B1(new_n817), .B2(G125), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n405), .B1(new_n864), .B2(G137), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1126), .B1(new_n804), .B2(new_n266), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1127), .A2(new_n1130), .A3(new_n1131), .A4(new_n1132), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n1070), .B1(new_n791), .B2(new_n476), .C1(new_n819), .C2(new_n868), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(G97), .A2(new_n816), .B1(new_n817), .B2(G294), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n296), .B1(new_n864), .B2(new_n583), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n858), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1135), .A2(new_n1136), .A3(new_n806), .A4(new_n1137), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n1125), .A2(new_n1133), .B1(new_n1134), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1122), .B1(new_n778), .B2(new_n1139), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1119), .A2(new_n992), .B1(new_n1120), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1118), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(KEYINPUT116), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT116), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1118), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n1143), .A2(new_n1145), .ZN(G378));
  NAND2_X1  g0946(.A1(new_n928), .A2(new_n926), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n929), .A2(new_n930), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1147), .A2(new_n1148), .A3(G330), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n323), .A2(new_n701), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n321), .B2(new_n326), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1150), .B(new_n325), .C1(new_n318), .C2(new_n320), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  OR3_X1    g0955(.A1(new_n1152), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1155), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1149), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n931), .A2(G330), .A3(new_n1158), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n922), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1160), .A2(new_n1161), .A3(new_n909), .A4(new_n921), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n992), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n766), .B1(G50), .B2(new_n855), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n296), .B(new_n722), .C1(G283), .C2(new_n817), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n542), .B2(new_n809), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1035), .B(new_n1169), .C1(G68), .C2(new_n861), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n791), .A2(new_n474), .B1(new_n801), .B2(new_n410), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G116), .B2(new_n799), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1170), .B(new_n1172), .C1(new_n571), .C2(new_n810), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT58), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n809), .A2(new_n859), .B1(new_n810), .B2(new_n867), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(G150), .A2(new_n861), .B1(new_n799), .B2(G125), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n1124), .B2(new_n791), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1176), .B(new_n1178), .C1(new_n805), .C2(new_n1129), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT59), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(G33), .A2(G41), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT117), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n801), .A2(new_n795), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n1184), .B(new_n1185), .C1(G124), .C2(new_n817), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1181), .A2(new_n1182), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1184), .B(new_n202), .C1(new_n296), .C2(new_n722), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n1189), .B(KEYINPUT118), .Z(new_n1190));
  NAND4_X1  g0990(.A1(new_n1175), .A2(new_n1187), .A3(new_n1188), .A4(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  OR2_X1    g0992(.A1(new_n1192), .A2(KEYINPUT119), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n777), .B1(new_n1192), .B2(KEYINPUT119), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1167), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n1158), .B2(new_n780), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1166), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1111), .A2(new_n1116), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1087), .B1(new_n1198), .B2(new_n1100), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n1165), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT57), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1201), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n724), .B1(new_n1199), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1197), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(G375));
  INV_X1    g1006(.A(new_n1097), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n923), .A2(new_n668), .A3(new_n1086), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1207), .A2(new_n1208), .A3(new_n1114), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n972), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1209), .A2(new_n1210), .A3(new_n1100), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n918), .A2(new_n853), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n766), .B1(G68), .B2(new_n855), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n799), .A2(G132), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT121), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n296), .B1(new_n810), .B2(new_n266), .C1(new_n809), .C2(new_n1128), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n786), .A2(new_n202), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n791), .A2(new_n867), .B1(new_n801), .B2(new_n410), .ZN(new_n1218));
  OR4_X1    g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n804), .A2(new_n795), .B1(new_n794), .B2(new_n1124), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT122), .Z(new_n1221));
  OAI22_X1  g1021(.A1(new_n868), .A2(new_n814), .B1(new_n801), .B2(new_n300), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(G283), .B2(new_n790), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n864), .A2(G116), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n296), .B1(new_n816), .B2(new_n583), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1223), .A2(new_n1037), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n804), .A2(new_n542), .B1(new_n794), .B2(new_n822), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT120), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n1219), .A2(new_n1221), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1213), .B1(new_n1229), .B2(new_n778), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1115), .A2(new_n992), .B1(new_n1212), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1211), .A2(new_n1231), .ZN(G381));
  NOR4_X1   g1032(.A1(G393), .A2(G381), .A3(G396), .A4(G384), .ZN(new_n1233));
  INV_X1    g1033(.A(G390), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1142), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  OR3_X1    g1036(.A1(new_n1236), .A2(G375), .A3(G387), .ZN(G407));
  NAND3_X1  g1037(.A1(new_n1205), .A2(new_n702), .A3(new_n1235), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(G407), .A2(G213), .A3(new_n1238), .ZN(G409));
  NAND3_X1  g1039(.A1(new_n993), .A2(new_n1020), .A3(G390), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(G393), .B(G396), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(G390), .B1(new_n993), .B2(new_n1020), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1242), .B1(KEYINPUT125), .B2(new_n1243), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1243), .A2(KEYINPUT125), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1241), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT124), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1243), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n1240), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1243), .A2(new_n1248), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1247), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1246), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(G213), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1254), .A2(G343), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1199), .A2(new_n1203), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1117), .A2(new_n1087), .B1(new_n1164), .B2(new_n1163), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1256), .B(new_n723), .C1(new_n1257), .C2(KEYINPUT57), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1197), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1258), .A2(new_n1143), .A3(new_n1145), .A4(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1200), .A2(new_n972), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1235), .B1(new_n1261), .B2(new_n1197), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1255), .B1(new_n1260), .B2(new_n1262), .ZN(new_n1263));
  XOR2_X1   g1063(.A(KEYINPUT123), .B(KEYINPUT60), .Z(new_n1264));
  NAND2_X1  g1064(.A1(new_n1209), .A2(new_n1264), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1207), .A2(KEYINPUT60), .A3(new_n1208), .A4(new_n1114), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1265), .A2(new_n723), .A3(new_n1100), .A4(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(G384), .A3(new_n1231), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(G384), .B1(new_n1267), .B2(new_n1231), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1263), .A2(KEYINPUT63), .A3(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1255), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1273), .A2(new_n1274), .A3(new_n1271), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT63), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1255), .A2(G2897), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1265), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1266), .A2(new_n723), .A3(new_n1100), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1231), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(G384), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1286), .A2(new_n1268), .A3(new_n1279), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1281), .A2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(KEYINPUT61), .B1(new_n1278), .B2(new_n1288), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1253), .A2(new_n1272), .A3(new_n1277), .A4(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(G387), .A2(new_n1234), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(KEYINPUT124), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(new_n1249), .A3(new_n1240), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n1247), .A2(new_n1293), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT61), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1281), .A2(new_n1287), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1295), .B1(new_n1263), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT62), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1275), .A2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1263), .A2(KEYINPUT62), .A3(new_n1271), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1297), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1294), .B1(new_n1301), .B2(KEYINPUT126), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1300), .ZN(new_n1303));
  AOI21_X1  g1103(.A(KEYINPUT62), .B1(new_n1263), .B2(new_n1271), .ZN(new_n1304));
  OAI211_X1 g1104(.A(KEYINPUT126), .B(new_n1289), .C1(new_n1303), .C2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1290), .B1(new_n1302), .B2(new_n1306), .ZN(G405));
  NAND2_X1  g1107(.A1(G375), .A2(new_n1235), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT127), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1308), .A2(new_n1309), .A3(new_n1260), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1309), .B1(new_n1308), .B2(new_n1260), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1271), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1312), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1271), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1314), .A2(new_n1315), .A3(new_n1310), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1313), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n1253), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1294), .A2(new_n1313), .A3(new_n1316), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(G402));
endmodule


