//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n566, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n639, new_n640, new_n641, new_n642, new_n643, new_n646,
    new_n648, new_n649, new_n650, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1256;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT65), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(KEYINPUT66), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n465), .A2(new_n470), .A3(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n461), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n467), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n468), .A2(new_n469), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n461), .ZN(new_n477));
  INV_X1    g052(.A(G137), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n473), .A2(new_n479), .ZN(G160));
  NOR2_X1   g055(.A1(new_n463), .A2(new_n464), .ZN(new_n481));
  OR3_X1    g056(.A1(new_n481), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n477), .A2(KEYINPUT67), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G112), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(G2105), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n481), .A2(new_n461), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G124), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n461), .B2(G114), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n495), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G102), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(new_n461), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n494), .A2(new_n496), .A3(G2104), .A4(new_n498), .ZN(new_n499));
  OAI211_X1 g074(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n499), .A2(KEYINPUT69), .A3(new_n500), .ZN(new_n504));
  INV_X1    g079(.A(G138), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n505), .A2(G2105), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n506), .B1(new_n463), .B2(new_n464), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT70), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n509));
  OAI211_X1 g084(.A(new_n506), .B(new_n509), .C1(new_n464), .C2(new_n463), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n508), .A2(KEYINPUT4), .A3(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT4), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n465), .A2(new_n470), .A3(new_n512), .A4(new_n506), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n503), .A2(new_n504), .B1(new_n511), .B2(new_n513), .ZN(G164));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  NAND3_X1  g090(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g092(.A(G543), .B1(KEYINPUT72), .B2(KEYINPUT5), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G62), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n515), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n517), .A2(new_n518), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n521), .A2(G651), .B1(new_n525), .B2(G88), .ZN(new_n526));
  OAI21_X1  g101(.A(G543), .B1(new_n522), .B2(new_n523), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n528), .A2(KEYINPUT71), .A3(G50), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n530));
  INV_X1    g105(.A(G50), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n526), .A2(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  NAND2_X1  g110(.A1(new_n525), .A2(G89), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n528), .A2(G51), .ZN(new_n538));
  NAND2_X1  g113(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n539));
  INV_X1    g114(.A(G543), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(new_n516), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n542), .A2(G63), .A3(G651), .ZN(new_n543));
  NAND3_X1  g118(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT7), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n538), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n537), .A2(new_n546), .ZN(G168));
  AOI22_X1  g122(.A1(new_n542), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G651), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G90), .ZN(new_n551));
  INV_X1    g126(.A(G52), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n524), .A2(new_n551), .B1(new_n527), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(G171));
  AOI22_X1  g129(.A1(new_n542), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(new_n549), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(G81), .ZN(new_n558));
  INV_X1    g133(.A(G43), .ZN(new_n559));
  OAI22_X1  g134(.A1(new_n524), .A2(new_n558), .B1(new_n527), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT73), .ZN(G188));
  NAND2_X1  g144(.A1(new_n525), .A2(G91), .ZN(new_n570));
  INV_X1    g145(.A(G53), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT74), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n571), .B1(new_n572), .B2(KEYINPUT9), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n528), .B(new_n573), .C1(new_n572), .C2(KEYINPUT9), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  OAI211_X1 g150(.A(KEYINPUT74), .B(new_n575), .C1(new_n527), .C2(new_n571), .ZN(new_n576));
  AND3_X1   g151(.A1(new_n570), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(G65), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n519), .A2(KEYINPUT76), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n542), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n578), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(G78), .A2(G543), .ZN(new_n583));
  XOR2_X1   g158(.A(new_n583), .B(KEYINPUT75), .Z(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n577), .A2(new_n585), .ZN(G299));
  INV_X1    g161(.A(G171), .ZN(G301));
  INV_X1    g162(.A(G168), .ZN(G286));
  OAI211_X1 g163(.A(G49), .B(G543), .C1(new_n522), .C2(new_n523), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT77), .Z(new_n590));
  OR3_X1    g165(.A1(new_n517), .A2(G74), .A3(new_n518), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n525), .A2(G87), .B1(new_n591), .B2(G651), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n590), .A2(new_n592), .ZN(G288));
  NAND2_X1  g168(.A1(new_n542), .A2(G61), .ZN(new_n594));
  NAND2_X1  g169(.A1(G73), .A2(G543), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n549), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(G86), .ZN(new_n597));
  INV_X1    g172(.A(G48), .ZN(new_n598));
  OAI22_X1  g173(.A1(new_n524), .A2(new_n597), .B1(new_n527), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(KEYINPUT78), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT78), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(new_n596), .B2(new_n599), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G305));
  INV_X1    g180(.A(G85), .ZN(new_n606));
  INV_X1    g181(.A(G47), .ZN(new_n607));
  OAI22_X1  g182(.A1(new_n524), .A2(new_n606), .B1(new_n527), .B2(new_n607), .ZN(new_n608));
  AND2_X1   g183(.A1(new_n542), .A2(G60), .ZN(new_n609));
  AND2_X1   g184(.A1(G72), .A2(G543), .ZN(new_n610));
  OAI21_X1  g185(.A(G651), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT79), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n608), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT80), .ZN(new_n614));
  OAI211_X1 g189(.A(KEYINPUT79), .B(G651), .C1(new_n609), .C2(new_n610), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n614), .B1(new_n613), .B2(new_n615), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(G290));
  NAND2_X1  g195(.A1(G301), .A2(G868), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT10), .ZN(new_n622));
  INV_X1    g197(.A(G92), .ZN(new_n623));
  OAI21_X1  g198(.A(KEYINPUT81), .B1(new_n524), .B2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  NOR3_X1   g200(.A1(new_n524), .A2(KEYINPUT81), .A3(new_n623), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n622), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(new_n626), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n628), .A2(KEYINPUT10), .A3(new_n624), .ZN(new_n629));
  INV_X1    g204(.A(G66), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n630), .B1(new_n579), .B2(new_n581), .ZN(new_n631));
  AND2_X1   g206(.A1(G79), .A2(G543), .ZN(new_n632));
  OAI21_X1  g207(.A(G651), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n528), .A2(G54), .ZN(new_n634));
  NAND4_X1  g209(.A1(new_n627), .A2(new_n629), .A3(new_n633), .A4(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n621), .B1(new_n636), .B2(G868), .ZN(G321));
  XOR2_X1   g212(.A(G321), .B(KEYINPUT82), .Z(G284));
  NAND3_X1  g213(.A1(G286), .A2(KEYINPUT83), .A3(G868), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT83), .ZN(new_n640));
  INV_X1    g215(.A(G868), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n640), .B1(G168), .B2(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(G299), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n639), .B(new_n642), .C1(new_n643), .C2(G868), .ZN(G297));
  XOR2_X1   g219(.A(G297), .B(KEYINPUT84), .Z(G280));
  INV_X1    g220(.A(G559), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n636), .B1(new_n646), .B2(G860), .ZN(G148));
  OR3_X1    g222(.A1(new_n635), .A2(KEYINPUT85), .A3(G559), .ZN(new_n648));
  OAI21_X1  g223(.A(KEYINPUT85), .B1(new_n635), .B2(G559), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  MUX2_X1   g225(.A(new_n562), .B(new_n650), .S(G868), .Z(G323));
  XNOR2_X1  g226(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g227(.A1(new_n489), .A2(G123), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT86), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n484), .A2(G135), .ZN(new_n655));
  OAI21_X1  g230(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT88), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  OR3_X1    g234(.A1(new_n461), .A2(KEYINPUT87), .A3(G111), .ZN(new_n660));
  OAI21_X1  g235(.A(KEYINPUT87), .B1(new_n461), .B2(G111), .ZN(new_n661));
  NAND4_X1  g236(.A1(new_n658), .A2(new_n659), .A3(new_n660), .A4(new_n661), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n654), .A2(new_n655), .A3(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(G2096), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n465), .A2(new_n470), .A3(new_n474), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT12), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT13), .ZN(new_n668));
  INV_X1    g243(.A(G2100), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n665), .A2(new_n670), .A3(new_n671), .ZN(G156));
  XOR2_X1   g247(.A(KEYINPUT15), .B(G2435), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G2438), .ZN(new_n674));
  XOR2_X1   g249(.A(G2427), .B(G2430), .Z(new_n675));
  OR2_X1    g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT89), .B(KEYINPUT14), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n675), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2451), .B(G2454), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT16), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n679), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2443), .B(G2446), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1341), .B(G1348), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT90), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n684), .A2(new_n685), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n688), .A2(G14), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G401));
  INV_X1    g266(.A(KEYINPUT18), .ZN(new_n692));
  XOR2_X1   g267(.A(G2084), .B(G2090), .Z(new_n693));
  XNOR2_X1  g268(.A(G2067), .B(G2678), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(KEYINPUT17), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n693), .A2(new_n694), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n692), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(new_n669), .ZN(new_n699));
  XOR2_X1   g274(.A(G2072), .B(G2078), .Z(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n695), .B2(KEYINPUT18), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(new_n664), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n699), .B(new_n702), .ZN(G227));
  XNOR2_X1  g278(.A(G1981), .B(G1986), .ZN(new_n704));
  XOR2_X1   g279(.A(G1991), .B(G1996), .Z(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1956), .B(G2474), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n708), .A2(KEYINPUT91), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(KEYINPUT91), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1961), .B(G1966), .ZN(new_n711));
  OR3_X1    g286(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1971), .B(G1976), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT19), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT20), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n711), .B1(new_n709), .B2(new_n710), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n717), .A2(new_n714), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT92), .Z(new_n719));
  NOR2_X1   g294(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n712), .A2(new_n717), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT93), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(new_n714), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n707), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n720), .A2(new_n723), .A3(new_n707), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n706), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n725), .A2(new_n706), .A3(new_n726), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n704), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n729), .ZN(new_n731));
  INV_X1    g306(.A(new_n704), .ZN(new_n732));
  NOR3_X1   g307(.A1(new_n731), .A2(new_n727), .A3(new_n732), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(G229));
  INV_X1    g310(.A(G16), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G20), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT23), .Z(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G299), .B2(G16), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1956), .ZN(new_n740));
  INV_X1    g315(.A(G29), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G35), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G162), .B2(new_n741), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT29), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G2090), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n740), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT104), .ZN(new_n748));
  NOR2_X1   g323(.A1(G4), .A2(G16), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT96), .Z(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n635), .B2(new_n736), .ZN(new_n751));
  INV_X1    g326(.A(G1348), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n484), .A2(G141), .ZN(new_n754));
  NAND3_X1  g329(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT101), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT26), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n489), .A2(G129), .B1(G105), .B2(new_n474), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n756), .A2(new_n757), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AND3_X1   g336(.A1(new_n754), .A2(new_n758), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G29), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n763), .B(KEYINPUT102), .C1(G29), .C2(G32), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(KEYINPUT102), .B2(new_n763), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT27), .B(G1996), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n563), .A2(G16), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G16), .B2(G19), .ZN(new_n769));
  INV_X1    g344(.A(G1341), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n741), .A2(G27), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G164), .B2(new_n741), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G2078), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n736), .A2(G21), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G168), .B2(new_n736), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G1966), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT31), .B(G11), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT103), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT30), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n780), .A2(G28), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n741), .B1(new_n780), .B2(G28), .ZN(new_n782));
  OAI221_X1 g357(.A(new_n779), .B1(new_n781), .B2(new_n782), .C1(new_n663), .C2(new_n741), .ZN(new_n783));
  NOR4_X1   g358(.A1(new_n771), .A2(new_n774), .A3(new_n777), .A4(new_n783), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n751), .A2(new_n752), .ZN(new_n785));
  AND4_X1   g360(.A1(new_n753), .A2(new_n767), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n741), .A2(G26), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT100), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT28), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n489), .A2(G128), .ZN(new_n790));
  NOR2_X1   g365(.A1(G104), .A2(G2105), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT98), .ZN(new_n792));
  OAI21_X1  g367(.A(G2104), .B1(new_n461), .B2(G116), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n484), .A2(G140), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT97), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(KEYINPUT97), .B1(new_n484), .B2(G140), .ZN(new_n797));
  OAI221_X1 g372(.A(new_n790), .B1(new_n792), .B2(new_n793), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(G29), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n799), .A2(KEYINPUT99), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n799), .A2(KEYINPUT99), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n789), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(G2067), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(G34), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n805), .A2(KEYINPUT24), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n805), .A2(KEYINPUT24), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n741), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G160), .B2(new_n741), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(G2084), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n736), .A2(G5), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G171), .B2(new_n736), .ZN(new_n812));
  INV_X1    g387(.A(G1961), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n810), .B(new_n814), .C1(new_n770), .C2(new_n769), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n484), .A2(G139), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT25), .Z(new_n818));
  AND2_X1   g393(.A1(new_n465), .A2(new_n470), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n819), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n816), .B(new_n818), .C1(new_n461), .C2(new_n820), .ZN(new_n821));
  MUX2_X1   g396(.A(G33), .B(new_n821), .S(G29), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G2072), .ZN(new_n823));
  AOI211_X1 g398(.A(new_n815), .B(new_n823), .C1(new_n746), .C2(new_n745), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n748), .A2(new_n786), .A3(new_n804), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n736), .A2(G6), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n604), .B2(new_n736), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT32), .B(G1981), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n736), .A2(G22), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(G166), .B2(new_n736), .ZN(new_n831));
  INV_X1    g406(.A(G1971), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n736), .A2(G23), .ZN(new_n834));
  INV_X1    g409(.A(G288), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n835), .B2(new_n736), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT33), .B(G1976), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n829), .A2(new_n833), .A3(new_n838), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT34), .Z(new_n840));
  NOR2_X1   g415(.A1(new_n619), .A2(new_n736), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(new_n736), .B2(G24), .ZN(new_n842));
  INV_X1    g417(.A(G1986), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n741), .A2(G25), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT94), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n484), .A2(G131), .ZN(new_n847));
  OAI21_X1  g422(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n848));
  INV_X1    g423(.A(G107), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n848), .B1(new_n849), .B2(G2105), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(new_n489), .B2(G119), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n846), .B1(new_n852), .B2(G29), .ZN(new_n853));
  XNOR2_X1  g428(.A(KEYINPUT35), .B(G1991), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT95), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n853), .B(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(new_n842), .B2(new_n843), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n840), .A2(new_n844), .A3(new_n857), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n858), .A2(KEYINPUT36), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(KEYINPUT36), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n825), .B1(new_n859), .B2(new_n860), .ZN(G311));
  INV_X1    g436(.A(G311), .ZN(G150));
  AOI22_X1  g437(.A1(new_n542), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n863), .A2(new_n549), .ZN(new_n864));
  INV_X1    g439(.A(G93), .ZN(new_n865));
  INV_X1    g440(.A(G55), .ZN(new_n866));
  OAI22_X1  g441(.A1(new_n524), .A2(new_n865), .B1(new_n527), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(G860), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT37), .Z(new_n871));
  NAND2_X1  g446(.A1(new_n636), .A2(G559), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT38), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n868), .A2(new_n557), .A3(new_n561), .ZN(new_n874));
  OAI22_X1  g449(.A1(new_n556), .A2(new_n560), .B1(new_n864), .B2(new_n867), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n873), .B(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(G860), .B1(new_n877), .B2(new_n878), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n879), .A2(KEYINPUT105), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT105), .B1(new_n879), .B2(new_n880), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n871), .B1(new_n881), .B2(new_n882), .ZN(G145));
  NAND2_X1  g458(.A1(new_n484), .A2(G142), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n489), .A2(G130), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n461), .A2(G118), .ZN(new_n886));
  OAI21_X1  g461(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n884), .B(new_n885), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n667), .ZN(new_n889));
  INV_X1    g464(.A(new_n852), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n889), .A2(new_n890), .ZN(new_n893));
  NOR3_X1   g468(.A1(new_n892), .A2(new_n762), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n762), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n889), .A2(new_n890), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n895), .B1(new_n896), .B2(new_n891), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n798), .A2(new_n821), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n510), .A2(KEYINPUT4), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n509), .B1(new_n476), .B2(new_n506), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n513), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n501), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n798), .A2(new_n821), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n898), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n903), .B1(new_n898), .B2(new_n904), .ZN(new_n907));
  OAI22_X1  g482(.A1(new_n894), .A2(new_n897), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n907), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n762), .B1(new_n892), .B2(new_n893), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n896), .A2(new_n895), .A3(new_n891), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .A4(new_n905), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n491), .B(G160), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n913), .B(new_n663), .Z(new_n914));
  NAND3_X1  g489(.A1(new_n908), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G37), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n914), .B1(new_n908), .B2(new_n912), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT40), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT40), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n917), .A2(new_n922), .A3(new_n919), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n921), .A2(new_n923), .ZN(G395));
  NAND2_X1  g499(.A1(new_n635), .A2(G299), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n627), .A2(new_n629), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n633), .A2(new_n634), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n643), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n650), .A2(new_n876), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n650), .A2(new_n876), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n925), .B(new_n928), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n931), .ZN(new_n933));
  INV_X1    g508(.A(new_n925), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n635), .A2(G299), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT41), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT41), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n928), .A2(new_n937), .A3(new_n925), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n933), .A2(new_n939), .A3(new_n929), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT108), .B1(new_n932), .B2(new_n940), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n932), .A2(new_n940), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT108), .ZN(new_n943));
  XOR2_X1   g518(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(G305), .B1(new_n617), .B2(new_n618), .ZN(new_n946));
  INV_X1    g521(.A(new_n618), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n947), .A2(new_n604), .A3(new_n616), .ZN(new_n948));
  XNOR2_X1  g523(.A(G303), .B(G288), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n949), .B1(new_n946), .B2(new_n948), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n945), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OR2_X1    g527(.A1(new_n952), .A2(KEYINPUT107), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(KEYINPUT107), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n950), .A2(new_n951), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT42), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n953), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n941), .B1(new_n943), .B2(new_n958), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n957), .A2(new_n942), .A3(KEYINPUT108), .ZN(new_n960));
  OAI21_X1  g535(.A(G868), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n869), .A2(new_n641), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(G295));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n962), .ZN(G331));
  INV_X1    g539(.A(new_n546), .ZN(new_n965));
  NAND3_X1  g540(.A1(G171), .A2(new_n536), .A3(new_n965), .ZN(new_n966));
  OAI22_X1  g541(.A1(new_n537), .A2(new_n546), .B1(new_n550), .B2(new_n553), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n876), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n876), .A2(new_n968), .A3(KEYINPUT110), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT110), .B1(new_n876), .B2(new_n968), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n934), .A2(new_n969), .A3(new_n935), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n876), .A2(new_n968), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n939), .A2(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(G37), .B1(new_n976), .B2(new_n955), .ZN(new_n977));
  XNOR2_X1  g552(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT111), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n938), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n928), .A2(KEYINPUT111), .A3(new_n937), .A4(new_n925), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(new_n936), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n970), .A2(new_n975), .ZN(new_n983));
  OR2_X1    g558(.A1(new_n971), .A2(new_n972), .ZN(new_n984));
  AOI22_X1  g559(.A1(new_n982), .A2(new_n983), .B1(new_n974), .B2(new_n984), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n977), .B(new_n978), .C1(new_n985), .C2(new_n955), .ZN(new_n986));
  INV_X1    g561(.A(new_n978), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n939), .A2(new_n973), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n974), .A2(new_n975), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n988), .A2(new_n955), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n916), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n976), .A2(new_n955), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n987), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT44), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n986), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n982), .A2(new_n983), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n984), .A2(new_n974), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n955), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT43), .B1(new_n991), .B2(new_n998), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n977), .B(new_n978), .C1(new_n955), .C2(new_n976), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n994), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT112), .B1(new_n995), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT43), .ZN(new_n1003));
  INV_X1    g578(.A(new_n998), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1003), .B1(new_n1004), .B2(new_n977), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n991), .A2(new_n992), .A3(new_n987), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT44), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n986), .A2(new_n993), .A3(new_n994), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1002), .A2(new_n1010), .ZN(G397));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n1012));
  INV_X1    g587(.A(G1384), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n903), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT114), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1016));
  INV_X1    g591(.A(new_n479), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n471), .A2(new_n472), .ZN(new_n1018));
  OAI211_X1 g593(.A(G40), .B(new_n1017), .C1(new_n1018), .C2(new_n461), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT119), .B(G2084), .Z(new_n1020));
  NOR2_X1   g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(G1384), .B1(new_n901), .B2(new_n902), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n1023), .A3(new_n1012), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1015), .A2(new_n1016), .A3(new_n1021), .A4(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1966), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n1027));
  NOR3_X1   g602(.A1(G164), .A2(new_n1027), .A3(G1384), .ZN(new_n1028));
  INV_X1    g603(.A(G40), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n473), .A2(new_n1029), .A3(new_n479), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(new_n1022), .B2(KEYINPUT45), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1026), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT124), .B1(new_n1025), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1025), .A2(new_n1032), .A3(KEYINPUT124), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1034), .A2(G168), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT51), .ZN(new_n1037));
  INV_X1    g612(.A(G8), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1038), .B1(new_n1025), .B2(new_n1032), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(G168), .A2(new_n1038), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(KEYINPUT51), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n1036), .A2(new_n1039), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1035), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1042), .B1(new_n1045), .B2(new_n1033), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT62), .B1(new_n1044), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n1045), .A2(new_n1033), .A3(G286), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1039), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT62), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1052), .A2(new_n1053), .A3(new_n1046), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1038), .B1(new_n1030), .B2(new_n1022), .ZN(new_n1055));
  OAI21_X1  g630(.A(G1981), .B1(new_n596), .B2(new_n599), .ZN(new_n1056));
  INV_X1    g631(.A(G1981), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT117), .B1(new_n600), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n1059));
  NOR4_X1   g634(.A1(new_n596), .A2(new_n599), .A3(new_n1059), .A4(G1981), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1056), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT49), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1055), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1056), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n600), .A2(new_n1057), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n1059), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n600), .A2(KEYINPUT117), .A3(new_n1057), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1065), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1064), .B1(new_n1069), .B2(KEYINPUT49), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1061), .A2(KEYINPUT118), .A3(new_n1062), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1063), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n590), .A2(new_n592), .A3(new_n1073), .A4(G1976), .ZN(new_n1074));
  INV_X1    g649(.A(G1976), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT116), .B1(G288), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1055), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT52), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1079), .B1(new_n835), .B2(G1976), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1078), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1072), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n501), .B1(new_n511), .B2(new_n513), .ZN(new_n1083));
  NOR4_X1   g658(.A1(new_n1083), .A2(KEYINPUT114), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n899), .A2(new_n900), .ZN(new_n1085));
  INV_X1    g660(.A(new_n513), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n499), .A2(KEYINPUT69), .A3(new_n500), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT69), .B1(new_n499), .B2(new_n500), .ZN(new_n1088));
  OAI22_X1  g663(.A1(new_n1085), .A2(new_n1086), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1012), .B1(new_n1089), .B2(new_n1013), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1084), .A2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1091), .A2(new_n746), .A3(new_n1030), .A4(new_n1015), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n903), .A2(KEYINPUT45), .A3(new_n1013), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n1030), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT45), .B1(new_n1089), .B2(new_n1013), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n832), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT113), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n503), .A2(new_n504), .ZN(new_n1098));
  AOI21_X1  g673(.A(G1384), .B1(new_n1098), .B2(new_n901), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1093), .B(new_n1030), .C1(new_n1099), .C2(KEYINPUT45), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT113), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1100), .A2(new_n1101), .A3(new_n832), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1092), .A2(new_n1097), .A3(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(G166), .A2(new_n1038), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT115), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1105), .A2(KEYINPUT55), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1108), .B1(new_n1104), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1103), .A2(G8), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1110), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1089), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT50), .B1(new_n1083), .B2(G1384), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(new_n1114), .A3(new_n1030), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1115), .A2(G2090), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1116), .B1(new_n832), .B2(new_n1100), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1112), .B1(new_n1117), .B2(new_n1038), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1082), .A2(new_n1111), .A3(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1015), .A2(new_n1016), .A3(new_n1030), .A4(new_n1024), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n813), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1122));
  INV_X1    g697(.A(G2078), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1122), .A2(KEYINPUT53), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n1100), .B2(G2078), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1121), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(G171), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1119), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1048), .A2(new_n1054), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1063), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(G288), .A2(G1976), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1133), .A2(new_n1134), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1055), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1082), .ZN(new_n1137));
  OAI22_X1  g712(.A1(new_n1135), .A2(new_n1136), .B1(new_n1137), .B2(new_n1111), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT63), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT120), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1040), .A2(new_n1140), .A3(G168), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1140), .B1(new_n1040), .B2(G168), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1139), .B1(new_n1119), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1103), .A2(G8), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1139), .B1(new_n1146), .B2(new_n1112), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1025), .A2(new_n1032), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1148), .A2(G8), .A3(G168), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(KEYINPUT120), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n1141), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1147), .A2(new_n1111), .A3(new_n1082), .A4(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1138), .B1(new_n1145), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(G1956), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1115), .A2(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g730(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(G299), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n577), .A2(new_n585), .A3(new_n1156), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1027), .B1(G164), .B2(G1384), .ZN(new_n1161));
  XNOR2_X1  g736(.A(KEYINPUT56), .B(G2072), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1161), .A2(new_n1030), .A3(new_n1093), .A4(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1155), .A2(new_n1160), .A3(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1120), .A2(new_n752), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1030), .A2(new_n1022), .A3(new_n803), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n636), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1160), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1019), .B1(new_n1099), .B2(new_n1012), .ZN(new_n1171));
  AOI21_X1  g746(.A(G1956), .B1(new_n1171), .B2(new_n1114), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1162), .ZN(new_n1173));
  NOR3_X1   g748(.A1(new_n1094), .A2(new_n1095), .A3(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1170), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1165), .B1(new_n1169), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(KEYINPUT60), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1166), .A2(KEYINPUT60), .A3(new_n1167), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n636), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1166), .A2(KEYINPUT60), .A3(new_n635), .A4(new_n1167), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1177), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1164), .A2(KEYINPUT122), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT122), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1155), .A2(new_n1160), .A3(new_n1183), .A4(new_n1163), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1182), .A2(KEYINPUT61), .A3(new_n1175), .A4(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1030), .A2(new_n1022), .ZN(new_n1186));
  XOR2_X1   g761(.A(KEYINPUT58), .B(G1341), .Z(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1188), .B1(new_n1100), .B2(G1996), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(new_n563), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT59), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1189), .A2(new_n1192), .A3(new_n563), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT61), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1160), .B1(new_n1155), .B2(new_n1163), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1195), .B1(new_n1165), .B2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1185), .A2(new_n1194), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1181), .B1(new_n1198), .B2(KEYINPUT123), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT123), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1185), .A2(new_n1194), .A3(new_n1197), .A4(new_n1200), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1176), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1052), .A2(new_n1046), .ZN(new_n1203));
  XNOR2_X1  g778(.A(KEYINPUT125), .B(KEYINPUT54), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1093), .A2(KEYINPUT53), .A3(new_n1123), .ZN(new_n1205));
  OR2_X1    g780(.A1(new_n1205), .A2(new_n1031), .ZN(new_n1206));
  NAND4_X1  g781(.A1(new_n1121), .A2(G301), .A3(new_n1126), .A4(new_n1206), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1204), .B1(new_n1128), .B2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n1119), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1121), .A2(new_n1126), .A3(new_n1206), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1210), .A2(G171), .ZN(new_n1211));
  OAI211_X1 g786(.A(new_n1211), .B(KEYINPUT54), .C1(G171), .C2(new_n1127), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1203), .A2(new_n1209), .A3(new_n1212), .ZN(new_n1213));
  OAI211_X1 g788(.A(new_n1130), .B(new_n1153), .C1(new_n1202), .C2(new_n1213), .ZN(new_n1214));
  NOR3_X1   g789(.A1(new_n1019), .A2(new_n1022), .A3(KEYINPUT45), .ZN(new_n1215));
  XNOR2_X1  g790(.A(new_n798), .B(new_n803), .ZN(new_n1216));
  XNOR2_X1  g791(.A(new_n762), .B(G1996), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n890), .A2(new_n855), .ZN(new_n1218));
  OR2_X1    g793(.A1(new_n890), .A2(new_n855), .ZN(new_n1219));
  NAND4_X1  g794(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(G290), .A2(G1986), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n619), .A2(new_n843), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1215), .B1(new_n1220), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1214), .A2(new_n1224), .ZN(new_n1225));
  NOR2_X1   g800(.A1(new_n798), .A2(G2067), .ZN(new_n1226));
  INV_X1    g801(.A(new_n1226), .ZN(new_n1227));
  INV_X1    g802(.A(new_n1215), .ZN(new_n1228));
  AOI21_X1  g803(.A(new_n1228), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1229));
  OAI21_X1  g804(.A(new_n1227), .B1(new_n1229), .B2(new_n1218), .ZN(new_n1230));
  INV_X1    g805(.A(KEYINPUT126), .ZN(new_n1231));
  OR2_X1    g806(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1233));
  NAND3_X1  g808(.A1(new_n1232), .A2(new_n1215), .A3(new_n1233), .ZN(new_n1234));
  NOR2_X1   g809(.A1(new_n1228), .A2(G1996), .ZN(new_n1235));
  XNOR2_X1  g810(.A(new_n1235), .B(KEYINPUT46), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n1216), .A2(new_n762), .ZN(new_n1237));
  AOI21_X1  g812(.A(new_n1236), .B1(new_n1237), .B2(new_n1215), .ZN(new_n1238));
  XOR2_X1   g813(.A(new_n1238), .B(KEYINPUT47), .Z(new_n1239));
  NAND2_X1  g814(.A1(new_n1220), .A2(new_n1215), .ZN(new_n1240));
  OR2_X1    g815(.A1(new_n1240), .A2(KEYINPUT127), .ZN(new_n1241));
  NAND2_X1  g816(.A1(new_n1240), .A2(KEYINPUT127), .ZN(new_n1242));
  NOR2_X1   g817(.A1(new_n1222), .A2(new_n1228), .ZN(new_n1243));
  XOR2_X1   g818(.A(new_n1243), .B(KEYINPUT48), .Z(new_n1244));
  NAND3_X1  g819(.A1(new_n1241), .A2(new_n1242), .A3(new_n1244), .ZN(new_n1245));
  AND3_X1   g820(.A1(new_n1234), .A2(new_n1239), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g821(.A1(new_n1225), .A2(new_n1246), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g822(.A1(G227), .A2(new_n459), .ZN(new_n1249));
  INV_X1    g823(.A(new_n1249), .ZN(new_n1250));
  AOI21_X1  g824(.A(new_n1250), .B1(new_n687), .B2(new_n689), .ZN(new_n1251));
  OAI211_X1 g825(.A(new_n734), .B(new_n1251), .C1(new_n917), .C2(new_n919), .ZN(new_n1252));
  NAND2_X1  g826(.A1(new_n986), .A2(new_n993), .ZN(new_n1253));
  INV_X1    g827(.A(new_n1253), .ZN(new_n1254));
  NOR2_X1   g828(.A1(new_n1252), .A2(new_n1254), .ZN(G308));
  NAND2_X1  g829(.A1(new_n918), .A2(new_n920), .ZN(new_n1256));
  NAND4_X1  g830(.A1(new_n1256), .A2(new_n734), .A3(new_n1253), .A4(new_n1251), .ZN(G225));
endmodule


