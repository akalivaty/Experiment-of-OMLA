//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0 1 0 0 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1287, new_n1288, new_n1289, new_n1290, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  INV_X1    g0017(.A(G97), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n208), .B1(new_n214), .B2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT65), .Z(new_n222));
  INV_X1    g0022(.A(KEYINPUT1), .ZN(new_n223));
  OR2_X1    g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n222), .A2(new_n223), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n208), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT0), .ZN(new_n228));
  INV_X1    g0028(.A(KEYINPUT64), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(new_n206), .ZN(new_n230));
  NAND2_X1  g0030(.A1(KEYINPUT64), .A2(G20), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n202), .A2(G50), .ZN(new_n236));
  OAI22_X1  g0036(.A1(new_n227), .A2(new_n228), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  AOI21_X1  g0037(.A(new_n237), .B1(new_n228), .B2(new_n227), .ZN(new_n238));
  AND3_X1   g0038(.A1(new_n224), .A2(new_n225), .A3(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n217), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT2), .B(G226), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n243), .B(new_n247), .ZN(G358));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT66), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(G87), .B(G97), .Z(new_n253));
  XOR2_X1   g0053(.A(G107), .B(G116), .Z(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n252), .B(new_n255), .ZN(G351));
  OAI21_X1  g0056(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G150), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT64), .A2(G20), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT64), .A2(G20), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G33), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT8), .B(G58), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n257), .B(new_n259), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n233), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(new_n267), .ZN(new_n271));
  INV_X1    g0071(.A(G50), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n272), .B1(new_n205), .B2(G20), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n271), .A2(new_n273), .B1(new_n272), .B2(new_n270), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n275), .B(KEYINPUT9), .ZN(new_n276));
  OR2_X1    g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  AOI21_X1  g0078(.A(G1698), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G222), .ZN(new_n280));
  INV_X1    g0080(.A(G77), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT3), .B(G33), .ZN(new_n282));
  INV_X1    g0082(.A(G223), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(G1698), .ZN(new_n284));
  OAI221_X1 g0084(.A(new_n280), .B1(new_n281), .B2(new_n282), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n288));
  INV_X1    g0088(.A(G274), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(G1), .A3(G13), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n288), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n290), .B1(new_n294), .B2(G226), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n287), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G200), .ZN(new_n297));
  INV_X1    g0097(.A(G190), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n276), .B(new_n297), .C1(new_n298), .C2(new_n296), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT70), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT10), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n300), .A2(new_n301), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n275), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n307), .B1(new_n296), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT67), .ZN(new_n310));
  OR2_X1    g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(new_n310), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n311), .B(new_n312), .C1(G179), .C2(new_n296), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n303), .A2(new_n305), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n306), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n264), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT68), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n316), .B1(new_n317), .B2(new_n258), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n318), .B1(new_n317), .B2(new_n258), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT15), .B(G87), .ZN(new_n320));
  OAI22_X1  g0120(.A1(new_n263), .A2(new_n320), .B1(new_n281), .B2(new_n262), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n267), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n266), .A2(new_n233), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n323), .A2(KEYINPUT69), .A3(new_n269), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT69), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(new_n270), .B2(new_n267), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n205), .A2(G20), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(G77), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n270), .A2(new_n281), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n322), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G1698), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n282), .A2(G232), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G107), .ZN(new_n335));
  OAI221_X1 g0135(.A(new_n334), .B1(new_n335), .B2(new_n282), .C1(new_n284), .C2(new_n211), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n286), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n290), .B1(new_n294), .B2(G244), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(G179), .ZN(new_n340));
  AOI21_X1  g0140(.A(G169), .B1(new_n337), .B2(new_n338), .ZN(new_n341));
  NOR3_X1   g0141(.A1(new_n332), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n331), .B1(G200), .B2(new_n339), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n344), .B1(new_n298), .B2(new_n339), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n315), .A2(new_n346), .ZN(new_n347));
  AND2_X1   g0147(.A1(G58), .A2(G68), .ZN(new_n348));
  OAI21_X1  g0148(.A(G20), .B1(new_n348), .B2(new_n201), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n258), .A2(G159), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  AND2_X1   g0152(.A1(KEYINPUT3), .A2(G33), .ZN(new_n353));
  NOR2_X1   g0153(.A1(KEYINPUT3), .A2(G33), .ZN(new_n354));
  NOR3_X1   g0154(.A1(new_n353), .A2(new_n354), .A3(G20), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT7), .ZN(new_n356));
  OAI21_X1  g0156(.A(G68), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NOR3_X1   g0157(.A1(new_n232), .A2(new_n282), .A3(KEYINPUT7), .ZN(new_n358));
  OAI211_X1 g0158(.A(KEYINPUT16), .B(new_n352), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n267), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT7), .B1(new_n232), .B2(new_n282), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n355), .A2(new_n356), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(new_n362), .A3(G68), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT16), .B1(new_n363), .B2(new_n352), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT72), .B1(new_n360), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n352), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT16), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n277), .A2(new_n206), .A3(new_n278), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n210), .B1(new_n369), .B2(KEYINPUT7), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n353), .A2(new_n354), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n262), .A2(new_n371), .A3(new_n356), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n351), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n323), .B1(new_n373), .B2(KEYINPUT16), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT72), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n368), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n264), .B1(new_n205), .B2(G20), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n377), .A2(new_n271), .B1(new_n270), .B2(new_n264), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT73), .ZN(new_n379));
  XNOR2_X1  g0179(.A(new_n378), .B(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n365), .A2(new_n376), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G226), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G1698), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n282), .B(new_n383), .C1(G223), .C2(G1698), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G33), .A2(G87), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n292), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G179), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n293), .A2(new_n217), .B1(new_n289), .B2(new_n288), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  OR2_X1    g0189(.A1(new_n386), .A2(new_n388), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n389), .B1(new_n390), .B2(G169), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n381), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT18), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT18), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n381), .A2(new_n395), .A3(new_n392), .ZN(new_n396));
  INV_X1    g0196(.A(G200), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n386), .B2(new_n388), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(new_n390), .B2(G190), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n365), .A2(new_n399), .A3(new_n376), .A4(new_n380), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT17), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n376), .A2(new_n380), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n403), .A2(KEYINPUT17), .A3(new_n365), .A4(new_n399), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n394), .A2(new_n396), .A3(new_n402), .A4(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n279), .A2(G226), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n282), .A2(G232), .A3(G1698), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G97), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n286), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT13), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n290), .B1(new_n294), .B2(G238), .ZN(new_n413));
  AND3_X1   g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n412), .B1(new_n411), .B2(new_n413), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT14), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n416), .A2(new_n417), .A3(G169), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n414), .A2(new_n415), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT14), .B1(new_n419), .B2(new_n308), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT71), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n421), .B1(new_n419), .B2(G179), .ZN(new_n422));
  NOR4_X1   g0222(.A1(new_n414), .A2(new_n415), .A3(KEYINPUT71), .A4(new_n387), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n418), .B(new_n420), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n262), .A2(G33), .A3(G77), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n258), .A2(G50), .B1(G20), .B2(new_n210), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n323), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n427), .A2(KEYINPUT11), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT12), .B1(new_n269), .B2(G68), .ZN(new_n429));
  OR3_X1    g0229(.A1(new_n269), .A2(KEYINPUT12), .A3(G68), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n427), .A2(KEYINPUT11), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n327), .A2(G68), .A3(new_n328), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n428), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n424), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n416), .A2(G200), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n433), .B1(new_n419), .B2(G190), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n347), .A2(new_n406), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n205), .A2(G45), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n440), .A2(new_n289), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n213), .B1(new_n205), .B2(G45), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n292), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT76), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n442), .A2(new_n292), .A3(KEYINPUT76), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n441), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(G244), .B(G1698), .C1(new_n353), .C2(new_n354), .ZN(new_n448));
  OAI211_X1 g0248(.A(G238), .B(new_n333), .C1(new_n353), .C2(new_n354), .ZN(new_n449));
  NAND2_X1  g0249(.A1(G33), .A2(G116), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n286), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n447), .A2(new_n452), .A3(new_n387), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT77), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT77), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n447), .A2(new_n452), .A3(new_n455), .A4(new_n387), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n451), .A2(new_n286), .ZN(new_n457));
  INV_X1    g0257(.A(new_n446), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT76), .B1(new_n442), .B2(new_n292), .ZN(new_n459));
  OAI22_X1  g0259(.A1(new_n458), .A2(new_n459), .B1(new_n289), .B2(new_n440), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n308), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n230), .A2(G33), .A3(G97), .A4(new_n231), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT19), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n262), .A2(new_n282), .A3(G68), .ZN(new_n465));
  NAND3_X1  g0265(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n230), .A2(new_n231), .A3(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(G97), .A2(G107), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n212), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n464), .A2(new_n465), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n267), .ZN(new_n472));
  INV_X1    g0272(.A(new_n320), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(new_n269), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(KEYINPUT78), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n205), .A2(G33), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n269), .A2(new_n477), .A3(new_n233), .A4(new_n266), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT78), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n320), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n476), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n472), .A2(new_n475), .A3(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n454), .A2(new_n456), .A3(new_n461), .A4(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT79), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n447), .A2(new_n452), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G200), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n478), .A2(new_n212), .ZN(new_n488));
  AOI211_X1 g0288(.A(new_n474), .B(new_n488), .C1(new_n471), .C2(new_n267), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n447), .A2(new_n452), .A3(G190), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n487), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n484), .A2(new_n485), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n485), .B1(new_n484), .B2(new_n491), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n361), .A2(new_n362), .A3(G107), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT6), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n218), .A2(new_n335), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n497), .B1(new_n498), .B2(new_n468), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n335), .A2(KEYINPUT6), .A3(G97), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n232), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n258), .A2(G77), .ZN(new_n503));
  XOR2_X1   g0303(.A(new_n503), .B(KEYINPUT74), .Z(new_n504));
  NAND3_X1  g0304(.A1(new_n496), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n267), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n269), .A2(G97), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n507), .B1(new_n479), .B2(G97), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g0309(.A(KEYINPUT5), .B(G41), .ZN(new_n510));
  INV_X1    g0310(.A(G45), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(G1), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n510), .A2(new_n292), .A3(G274), .A4(new_n512), .ZN(new_n513));
  AND2_X1   g0313(.A1(KEYINPUT5), .A2(G41), .ZN(new_n514));
  NOR2_X1   g0314(.A1(KEYINPUT5), .A2(G41), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n292), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n513), .B1(new_n517), .B2(new_n219), .ZN(new_n518));
  OAI211_X1 g0318(.A(G244), .B(new_n333), .C1(new_n353), .C2(new_n354), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT4), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n282), .A2(KEYINPUT4), .A3(G244), .A4(new_n333), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G33), .A2(G283), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n282), .A2(G250), .A3(G1698), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n521), .A2(new_n522), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n518), .B1(new_n525), .B2(new_n286), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n387), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n286), .ZN(new_n528));
  INV_X1    g0328(.A(new_n518), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n308), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n509), .A2(new_n527), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n508), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n533), .B1(new_n505), .B2(new_n267), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n528), .A2(new_n298), .A3(new_n529), .ZN(new_n535));
  AOI21_X1  g0335(.A(G200), .B1(new_n528), .B2(new_n529), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT75), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT75), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n539), .B(new_n534), .C1(new_n535), .C2(new_n536), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n532), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT21), .ZN(new_n542));
  OAI211_X1 g0342(.A(G264), .B(G1698), .C1(new_n353), .C2(new_n354), .ZN(new_n543));
  OAI211_X1 g0343(.A(G257), .B(new_n333), .C1(new_n353), .C2(new_n354), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n277), .A2(G303), .A3(new_n278), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n546), .A2(KEYINPUT80), .A3(new_n286), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(KEYINPUT80), .B1(new_n546), .B2(new_n286), .ZN(new_n549));
  INV_X1    g0349(.A(G270), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n513), .B1(new_n517), .B2(new_n550), .ZN(new_n551));
  NOR3_X1   g0351(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(G116), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n553), .B1(new_n205), .B2(G33), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n324), .A2(new_n326), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n270), .A2(new_n553), .ZN(new_n556));
  INV_X1    g0356(.A(G33), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G97), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n230), .A2(new_n558), .A3(new_n231), .A4(new_n523), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n266), .A2(new_n233), .B1(G20), .B2(new_n553), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n559), .A2(KEYINPUT20), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT20), .B1(new_n559), .B2(new_n560), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n555), .B(new_n556), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G169), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n542), .B1(new_n552), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n552), .A2(G179), .A3(new_n563), .ZN(new_n566));
  INV_X1    g0366(.A(new_n549), .ZN(new_n567));
  INV_X1    g0367(.A(new_n551), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(new_n568), .A3(new_n547), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n569), .A2(KEYINPUT21), .A3(G169), .A4(new_n563), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n565), .A2(new_n566), .A3(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(G250), .B(new_n333), .C1(new_n353), .C2(new_n354), .ZN(new_n572));
  OAI211_X1 g0372(.A(G257), .B(G1698), .C1(new_n353), .C2(new_n354), .ZN(new_n573));
  NAND2_X1  g0373(.A1(G33), .A2(G294), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n286), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n286), .B1(new_n512), .B2(new_n510), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G264), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n578), .A3(new_n513), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n308), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n286), .A2(new_n575), .B1(new_n577), .B2(G264), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n581), .A2(new_n387), .A3(new_n513), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n262), .A2(new_n282), .A3(G87), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT22), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT22), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n262), .A2(new_n282), .A3(new_n586), .A4(G87), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT24), .ZN(new_n589));
  NAND2_X1  g0389(.A1(KEYINPUT23), .A2(G107), .ZN(new_n590));
  AOI21_X1  g0390(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n590), .B1(new_n591), .B2(G20), .ZN(new_n592));
  NOR2_X1   g0392(.A1(KEYINPUT23), .A2(G107), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n592), .B1(new_n232), .B2(new_n593), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n588), .A2(new_n589), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n589), .B1(new_n588), .B2(new_n594), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n267), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT25), .B1(new_n270), .B2(new_n335), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n270), .A2(KEYINPUT25), .A3(new_n335), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n599), .A2(new_n600), .B1(G107), .B2(new_n479), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n583), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n571), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n588), .A2(new_n594), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(KEYINPUT24), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n588), .A2(new_n589), .A3(new_n594), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n323), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n601), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(G200), .B1(new_n581), .B2(new_n513), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT81), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n579), .A2(new_n397), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT81), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n581), .A2(new_n298), .A3(new_n513), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n612), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n552), .A2(G190), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n563), .B1(new_n569), .B2(G200), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n609), .A2(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n495), .A2(new_n541), .A3(new_n603), .A4(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n439), .A2(new_n620), .ZN(G372));
  AND3_X1   g0421(.A1(new_n381), .A2(new_n395), .A3(new_n392), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n395), .B1(new_n381), .B2(new_n392), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n437), .A2(new_n342), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n434), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT83), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n404), .A2(new_n402), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n626), .A2(new_n627), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n624), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n306), .A2(new_n314), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n313), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n484), .A2(new_n491), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(KEYINPUT79), .ZN(new_n638));
  XOR2_X1   g0438(.A(KEYINPUT82), .B(KEYINPUT26), .Z(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n638), .A2(new_n492), .A3(new_n532), .A4(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT26), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n461), .A2(new_n483), .A3(new_n453), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n491), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n509), .A2(new_n531), .A3(new_n527), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n583), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n648), .B1(new_n607), .B2(new_n608), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n649), .A2(new_n566), .A3(new_n565), .A4(new_n570), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n644), .B1(new_n609), .B2(new_n616), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n541), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n647), .A2(new_n652), .A3(new_n643), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n636), .B1(new_n439), .B2(new_n654), .ZN(G369));
  INV_X1    g0455(.A(KEYINPUT84), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n205), .A2(G13), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n656), .B1(new_n232), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT27), .ZN(new_n659));
  INV_X1    g0459(.A(new_n657), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n262), .A2(KEYINPUT84), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n658), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G213), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n659), .B1(new_n658), .B2(new_n661), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT85), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n658), .A2(new_n661), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT85), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n667), .A2(new_n668), .A3(G213), .A4(new_n662), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G343), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT86), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT86), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n665), .A2(new_n669), .A3(new_n673), .A4(G343), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n563), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT87), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n676), .B(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n571), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n676), .B(KEYINPUT87), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n618), .A2(new_n617), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g0485(.A(KEYINPUT88), .B(G330), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n675), .A2(new_n649), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n615), .B1(new_n610), .B2(new_n611), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n613), .A2(KEYINPUT81), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n597), .B(new_n601), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n672), .A2(new_n674), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n691), .B1(new_n692), .B2(new_n609), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n688), .B1(new_n693), .B2(new_n649), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n685), .A2(new_n687), .A3(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n679), .A2(new_n675), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n688), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(G399));
  INV_X1    g0498(.A(new_n226), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(G41), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n469), .A2(G116), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G1), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n236), .B2(new_n701), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT28), .Z(new_n705));
  INV_X1    g0505(.A(KEYINPUT29), .ZN(new_n706));
  INV_X1    g0506(.A(new_n644), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n691), .B(new_n707), .C1(new_n571), .C2(new_n602), .ZN(new_n708));
  INV_X1    g0508(.A(new_n540), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n528), .A2(new_n529), .A3(new_n298), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(G200), .B2(new_n526), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n539), .B1(new_n711), .B2(new_n534), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n645), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n643), .B1(new_n708), .B2(new_n713), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n644), .A2(new_n645), .A3(new_n642), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n638), .A2(new_n492), .A3(new_n532), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n715), .B1(new_n716), .B2(new_n639), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n692), .B1(new_n714), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(KEYINPUT91), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT91), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n720), .B(new_n692), .C1(new_n714), .C2(new_n717), .ZN(new_n721));
  AOI211_X1 g0521(.A(KEYINPUT92), .B(new_n706), .C1(new_n719), .C2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT92), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n719), .A2(new_n721), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(KEYINPUT29), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n641), .A2(new_n646), .ZN(new_n726));
  OAI211_X1 g0526(.A(KEYINPUT90), .B(new_n692), .C1(new_n726), .C2(new_n714), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(KEYINPUT90), .B1(new_n653), .B2(new_n692), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n706), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n722), .B1(new_n725), .B2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT31), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n579), .A2(new_n486), .A3(new_n387), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(new_n569), .A3(new_n530), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT30), .ZN(new_n736));
  INV_X1    g0536(.A(new_n486), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(new_n526), .A3(new_n581), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n567), .A2(new_n568), .A3(G179), .A4(new_n547), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n736), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT89), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n735), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n737), .A2(new_n526), .A3(new_n581), .ZN(new_n743));
  INV_X1    g0543(.A(new_n739), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n743), .A2(new_n744), .A3(KEYINPUT30), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(KEYINPUT89), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n742), .B1(new_n740), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n733), .B1(new_n747), .B2(new_n692), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n745), .A2(new_n740), .A3(new_n735), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(KEYINPUT31), .A3(new_n675), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n748), .B(new_n750), .C1(new_n620), .C2(new_n675), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n687), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n732), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n705), .B1(new_n753), .B2(new_n205), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n754), .B(KEYINPUT93), .Z(G364));
  NOR2_X1   g0555(.A1(G179), .A2(G200), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n232), .A2(new_n298), .A3(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n758), .A2(G329), .ZN(new_n759));
  INV_X1    g0559(.A(G303), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n397), .A2(G179), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n761), .A2(G20), .A3(G190), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n262), .B1(G190), .B2(new_n756), .ZN(new_n763));
  INV_X1    g0563(.A(G294), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n371), .B1(new_n760), .B2(new_n762), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n232), .A2(new_n298), .A3(new_n761), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n759), .B(new_n765), .C1(G283), .C2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n262), .A2(new_n387), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n770), .A2(KEYINPUT97), .ZN(new_n771));
  AOI21_X1  g0571(.A(G200), .B1(new_n770), .B2(KEYINPUT97), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n771), .A2(G190), .A3(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G322), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n771), .A2(new_n298), .A3(new_n772), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G311), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n769), .A2(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n298), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n769), .A2(new_n298), .A3(G200), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  XNOR2_X1  g0582(.A(KEYINPUT33), .B(G317), .ZN(new_n783));
  AOI22_X1  g0583(.A1(G326), .A2(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n768), .A2(new_n775), .A3(new_n778), .A4(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n282), .B1(new_n762), .B2(new_n212), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n763), .A2(new_n218), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n786), .B(new_n787), .C1(G107), .C2(new_n767), .ZN(new_n788));
  INV_X1    g0588(.A(G159), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n757), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT32), .ZN(new_n791));
  AOI22_X1  g0591(.A1(G50), .A2(new_n780), .B1(new_n782), .B2(G68), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n788), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n216), .A2(new_n773), .B1(new_n776), .B2(new_n281), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n785), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT95), .ZN(new_n796));
  OAI21_X1  g0596(.A(G20), .B1(new_n796), .B2(G169), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n308), .A2(KEYINPUT95), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n234), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n799), .A2(KEYINPUT96), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(KEYINPUT96), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n795), .A2(new_n802), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n262), .A2(G13), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n205), .B1(new_n804), .B2(G45), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n700), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n252), .A2(G45), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n226), .A2(new_n371), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT94), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n809), .B(new_n811), .C1(G45), .C2(new_n236), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n699), .A2(new_n371), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n813), .A2(G355), .B1(new_n553), .B2(new_n699), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(G13), .A2(G33), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(G20), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n802), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n808), .B1(new_n815), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n818), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n803), .B(new_n820), .C1(new_n685), .C2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n685), .A2(new_n687), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n808), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n685), .A2(new_n687), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n822), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT98), .Z(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(G396));
  NOR2_X1   g0628(.A1(new_n343), .A2(new_n675), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n675), .A2(new_n331), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n342), .B1(new_n830), .B2(new_n345), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n730), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n831), .A2(new_n829), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n653), .A2(new_n833), .A3(new_n692), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n807), .B1(new_n835), .B2(new_n752), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n752), .B2(new_n835), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n802), .A2(new_n816), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n808), .B1(new_n838), .B2(new_n281), .ZN(new_n839));
  INV_X1    g0639(.A(new_n762), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n282), .B(new_n787), .C1(G107), .C2(new_n840), .ZN(new_n841));
  AOI22_X1  g0641(.A1(G87), .A2(new_n767), .B1(new_n758), .B2(G311), .ZN(new_n842));
  INV_X1    g0642(.A(new_n780), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n841), .B(new_n842), .C1(new_n760), .C2(new_n843), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n781), .B(KEYINPUT99), .ZN(new_n845));
  XNOR2_X1  g0645(.A(KEYINPUT100), .B(G283), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n777), .A2(G116), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n848), .A2(KEYINPUT101), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n844), .B(new_n849), .C1(G294), .C2(new_n774), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n848), .A2(KEYINPUT101), .ZN(new_n851));
  AOI22_X1  g0651(.A1(G137), .A2(new_n780), .B1(new_n782), .B2(G150), .ZN(new_n852));
  INV_X1    g0652(.A(G143), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n852), .B1(new_n853), .B2(new_n773), .C1(new_n789), .C2(new_n776), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT34), .ZN(new_n855));
  OR2_X1    g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(G132), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n282), .B1(new_n272), .B2(new_n762), .C1(new_n757), .C2(new_n857), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n763), .A2(new_n216), .B1(new_n766), .B2(new_n210), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n858), .B(new_n859), .C1(new_n854), .C2(new_n855), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n850), .A2(new_n851), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n802), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n839), .B1(new_n833), .B2(new_n817), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n837), .A2(new_n863), .ZN(G384));
  INV_X1    g0664(.A(new_n439), .ZN(new_n865));
  NOR3_X1   g0665(.A1(new_n728), .A2(new_n729), .A3(KEYINPUT29), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n706), .B1(new_n719), .B2(new_n721), .ZN(new_n867));
  NOR3_X1   g0667(.A1(new_n866), .A2(new_n867), .A3(new_n723), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n865), .B1(new_n868), .B2(new_n722), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n636), .ZN(new_n870));
  XOR2_X1   g0670(.A(new_n870), .B(KEYINPUT106), .Z(new_n871));
  NOR2_X1   g0671(.A1(new_n434), .A2(new_n675), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT38), .ZN(new_n874));
  INV_X1    g0674(.A(new_n378), .ZN(new_n875));
  OR2_X1    g0675(.A1(new_n373), .A2(KEYINPUT16), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n875), .B1(new_n876), .B2(new_n374), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n877), .A2(new_n670), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n629), .B2(new_n624), .ZN(new_n880));
  INV_X1    g0680(.A(new_n670), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n381), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT37), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n393), .A2(new_n882), .A3(new_n883), .A4(new_n400), .ZN(new_n884));
  INV_X1    g0684(.A(new_n400), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n877), .B1(new_n391), .B2(new_n670), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT37), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n874), .B1(new_n880), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n405), .A2(new_n878), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT103), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n891), .A2(new_n892), .A3(KEYINPUT38), .A4(new_n888), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n405), .A2(new_n878), .B1(new_n884), .B2(new_n887), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n892), .B1(new_n895), .B2(KEYINPUT38), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT39), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n891), .A2(KEYINPUT38), .A3(new_n888), .ZN(new_n898));
  XOR2_X1   g0698(.A(KEYINPUT105), .B(KEYINPUT39), .Z(new_n899));
  AOI21_X1  g0699(.A(new_n882), .B1(new_n629), .B2(new_n624), .ZN(new_n900));
  INV_X1    g0700(.A(new_n884), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n393), .A2(new_n882), .A3(new_n400), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT37), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n901), .B1(KEYINPUT104), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT104), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n902), .A2(new_n905), .A3(KEYINPUT37), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n900), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n898), .B(new_n899), .C1(new_n907), .C2(KEYINPUT38), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n873), .B1(new_n897), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n894), .A2(new_n896), .ZN(new_n910));
  INV_X1    g0710(.A(new_n829), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n834), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n675), .A2(new_n433), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n434), .A2(new_n437), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n424), .A2(new_n433), .A3(new_n675), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  OAI22_X1  g0717(.A1(new_n910), .A2(new_n917), .B1(new_n624), .B2(new_n881), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n909), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n871), .B(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT40), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n898), .B1(new_n907), .B2(KEYINPUT38), .ZN(new_n923));
  INV_X1    g0723(.A(new_n735), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT30), .B1(new_n743), .B2(new_n744), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n924), .B1(new_n925), .B2(KEYINPUT89), .ZN(new_n926));
  NOR3_X1   g0726(.A1(new_n738), .A2(new_n739), .A3(new_n736), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n740), .B1(new_n927), .B2(new_n741), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n692), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT31), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n748), .B(new_n930), .C1(new_n620), .C2(new_n675), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n931), .A2(new_n833), .A3(new_n916), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n922), .B1(new_n923), .B2(new_n932), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n931), .A2(new_n922), .A3(new_n833), .A4(new_n916), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n910), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n931), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n439), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n936), .B(new_n938), .Z(new_n939));
  NOR2_X1   g0739(.A1(new_n939), .A2(new_n686), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n921), .A2(new_n940), .B1(new_n205), .B2(new_n804), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n921), .B2(new_n940), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n501), .B(KEYINPUT102), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n943), .A2(KEYINPUT35), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n943), .A2(KEYINPUT35), .ZN(new_n945));
  NOR4_X1   g0745(.A1(new_n944), .A2(new_n945), .A3(new_n553), .A4(new_n235), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT36), .ZN(new_n947));
  OR3_X1    g0747(.A1(new_n236), .A2(new_n281), .A3(new_n348), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n272), .A2(G68), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n205), .B(G13), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  OR3_X1    g0750(.A1(new_n942), .A2(new_n947), .A3(new_n950), .ZN(G367));
  INV_X1    g0751(.A(new_n819), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n811), .A2(new_n246), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n226), .B2(new_n320), .ZN(new_n954));
  INV_X1    g0754(.A(new_n763), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n780), .A2(G143), .B1(G68), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(G150), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n956), .B1(new_n773), .B2(new_n957), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT110), .Z(new_n959));
  NAND2_X1  g0759(.A1(new_n767), .A2(G77), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n371), .B1(new_n840), .B2(G58), .ZN(new_n961));
  XNOR2_X1  g0761(.A(KEYINPUT111), .B(G137), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n960), .B(new_n961), .C1(new_n757), .C2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n777), .B2(G50), .ZN(new_n964));
  INV_X1    g0764(.A(new_n845), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n959), .B(new_n964), .C1(new_n789), .C2(new_n965), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n777), .A2(new_n847), .B1(G294), .B2(new_n845), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n774), .A2(G303), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n763), .A2(new_n335), .B1(new_n766), .B2(new_n218), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(G317), .B2(new_n758), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT46), .B1(new_n840), .B2(G116), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n840), .A2(KEYINPUT46), .A3(G116), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n371), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n971), .B(new_n973), .C1(G311), .C2(new_n780), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n967), .A2(new_n968), .A3(new_n970), .A4(new_n974), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n966), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(KEYINPUT47), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n802), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n976), .A2(KEYINPUT47), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n807), .B1(new_n952), .B2(new_n954), .C1(new_n978), .C2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n692), .A2(new_n489), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n981), .A2(new_n644), .ZN(new_n982));
  INV_X1    g0782(.A(new_n643), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n982), .B1(new_n983), .B2(new_n981), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n980), .B1(new_n818), .B2(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT112), .Z(new_n986));
  INV_X1    g0786(.A(KEYINPUT42), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n694), .A2(new_n696), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n675), .A2(new_n509), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n541), .A2(new_n989), .B1(new_n532), .B2(new_n675), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n987), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n990), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n694), .A2(new_n992), .A3(KEYINPUT42), .A4(new_n696), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n602), .B1(new_n709), .B2(new_n712), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n675), .B1(new_n995), .B2(new_n645), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT107), .ZN(new_n999));
  INV_X1    g0799(.A(new_n984), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n998), .A2(KEYINPUT43), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n996), .B1(new_n991), .B2(new_n993), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n984), .B1(new_n1003), .B2(KEYINPUT107), .ZN(new_n1004));
  AND3_X1   g0804(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT43), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1007));
  OAI21_X1  g0807(.A(KEYINPUT108), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(KEYINPUT43), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT108), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1008), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n695), .A2(new_n990), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1008), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AND2_X1   g0819(.A1(new_n732), .A2(new_n752), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT109), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT45), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n688), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n988), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1022), .B1(new_n1024), .B2(new_n990), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n697), .A2(KEYINPUT45), .A3(new_n992), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1024), .A2(KEYINPUT44), .A3(new_n990), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT44), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n697), .B2(new_n992), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  AND3_X1   g0831(.A1(new_n1027), .A2(new_n695), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n695), .B1(new_n1027), .B2(new_n1031), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1021), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1033), .A2(new_n1021), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n694), .B(new_n696), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n823), .B(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1020), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n700), .B(KEYINPUT41), .Z(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n806), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n986), .B1(new_n1019), .B2(new_n1042), .ZN(G387));
  INV_X1    g0843(.A(new_n702), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n813), .A2(new_n1044), .B1(new_n335), .B2(new_n699), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n243), .A2(new_n511), .ZN(new_n1046));
  AOI21_X1  g0846(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1047));
  AND3_X1   g0847(.A1(new_n316), .A2(KEYINPUT50), .A3(new_n272), .ZN(new_n1048));
  AOI21_X1  g0848(.A(KEYINPUT50), .B1(new_n316), .B2(new_n272), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n702), .B(new_n1047), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n811), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1045), .B1(new_n1046), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n808), .B1(new_n1052), .B2(new_n819), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n694), .B2(new_n821), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n282), .B1(new_n758), .B2(G326), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n845), .A2(G311), .B1(G322), .B2(new_n780), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n774), .A2(G317), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(new_n760), .C2(new_n776), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT114), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n1059), .A2(KEYINPUT48), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(KEYINPUT48), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n955), .A2(new_n847), .B1(new_n840), .B2(G294), .ZN(new_n1062));
  AND3_X1   g0862(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(KEYINPUT115), .B(KEYINPUT49), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1055), .B1(new_n553), .B2(new_n766), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n776), .A2(new_n210), .B1(new_n264), .B2(new_n781), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT113), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n282), .B1(new_n281), .B2(new_n762), .C1(new_n766), .C2(new_n218), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n476), .A2(new_n481), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n1071), .A2(new_n763), .B1(new_n957), .B2(new_n757), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1070), .B(new_n1072), .C1(G159), .C2(new_n780), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n272), .B2(new_n773), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1067), .B1(new_n1069), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1054), .B1(new_n1075), .B2(new_n802), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1038), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1076), .B1(new_n806), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1020), .A2(new_n1077), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n753), .A2(new_n1038), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n700), .B(KEYINPUT116), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1078), .A2(new_n1082), .ZN(G393));
  AOI22_X1  g0883(.A1(new_n811), .A2(new_n255), .B1(G97), .B2(new_n699), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n808), .B1(new_n1084), .B2(new_n819), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n774), .A2(G311), .B1(G317), .B2(new_n780), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT52), .Z(new_n1087));
  AOI22_X1  g0887(.A1(new_n955), .A2(G116), .B1(new_n758), .B2(G322), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n282), .B1(new_n840), .B2(new_n847), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1088), .B(new_n1089), .C1(new_n335), .C2(new_n766), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n776), .A2(new_n764), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1090), .B(new_n1091), .C1(G303), .C2(new_n845), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n773), .A2(new_n789), .B1(new_n957), .B2(new_n843), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT51), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n955), .A2(G77), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n767), .A2(G87), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n371), .B1(new_n840), .B2(G68), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n758), .A2(G143), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n776), .A2(new_n264), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1099), .B(new_n1100), .C1(G50), .C2(new_n845), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1087), .A2(new_n1092), .B1(new_n1094), .B2(new_n1101), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1085), .B1(new_n1102), .B2(new_n862), .C1(new_n821), .C2(new_n992), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1081), .B1(new_n1036), .B2(new_n1079), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1104), .B1(new_n1020), .B2(new_n1077), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1103), .B1(new_n805), .B2(new_n1105), .C1(new_n1106), .C2(new_n1107), .ZN(G390));
  AOI21_X1  g0908(.A(new_n831), .B1(new_n719), .B2(new_n721), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n916), .B1(new_n1109), .B2(new_n829), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n903), .A2(KEYINPUT104), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1111), .A2(new_n884), .A3(new_n906), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n406), .B2(new_n882), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n874), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n872), .B1(new_n1114), .B2(new_n898), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1110), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n917), .A2(new_n873), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1117), .A2(new_n897), .A3(new_n908), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n751), .A2(new_n687), .A3(new_n833), .A4(new_n916), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1116), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n898), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n1113), .B2(new_n874), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n898), .A2(KEYINPUT103), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1123), .A2(new_n893), .A3(new_n890), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1122), .A2(new_n899), .B1(new_n1124), .B2(KEYINPUT39), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1125), .A2(new_n1117), .B1(new_n1110), .B2(new_n1115), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n931), .A2(G330), .A3(new_n833), .A4(new_n916), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1120), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n938), .A2(G330), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n620), .A2(new_n675), .B1(new_n929), .B2(KEYINPUT31), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n750), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n687), .B(new_n833), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n916), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n1127), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n912), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n831), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n724), .A2(new_n1137), .ZN(new_n1138));
  NOR3_X1   g0938(.A1(new_n747), .A2(new_n733), .A3(new_n692), .ZN(new_n1139));
  OAI211_X1 g0939(.A(G330), .B(new_n833), .C1(new_n1130), .C2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n1133), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1138), .A2(new_n911), .A3(new_n1119), .A4(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1136), .A2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n869), .A2(new_n636), .A3(new_n1129), .A4(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1128), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n1081), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n636), .B(new_n1129), .C1(new_n732), .C2(new_n439), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1143), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1116), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1127), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT117), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1149), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(KEYINPUT117), .B1(new_n1128), .B2(new_n1144), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1146), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1125), .A2(new_n816), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n838), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n807), .B1(new_n1158), .B2(new_n316), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n763), .A2(new_n789), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n840), .A2(G150), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT53), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1160), .B(new_n1162), .C1(G125), .C2(new_n758), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n282), .B1(new_n766), .B2(new_n272), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n780), .B2(G128), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(KEYINPUT54), .B(G143), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1163), .B(new_n1165), .C1(new_n776), .C2(new_n1166), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n965), .A2(new_n962), .B1(new_n857), .B2(new_n773), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n965), .A2(new_n335), .B1(new_n553), .B2(new_n773), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1095), .B1(new_n764), .B2(new_n757), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n371), .B1(new_n212), .B2(new_n762), .C1(new_n766), .C2(new_n210), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n780), .A2(G283), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1172), .B(new_n1173), .C1(new_n218), .C2(new_n776), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n1167), .A2(new_n1168), .B1(new_n1169), .B2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1159), .B1(new_n1175), .B2(new_n802), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1157), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n1128), .B2(new_n805), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1156), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(G378));
  AOI21_X1  g0980(.A(new_n808), .B1(new_n838), .B2(new_n272), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n774), .A2(G128), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n777), .A2(G137), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n763), .A2(new_n957), .B1(new_n762), .B2(new_n1166), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n781), .A2(new_n857), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n1184), .B(new_n1185), .C1(G125), .C2(new_n780), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1182), .A2(new_n1183), .A3(new_n1186), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1187), .A2(KEYINPUT59), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(KEYINPUT59), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n767), .A2(G159), .ZN(new_n1190));
  AOI211_X1 g0990(.A(G33), .B(G41), .C1(new_n758), .C2(G124), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n780), .A2(G116), .B1(G68), .B2(new_n955), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1193), .B(KEYINPUT118), .Z(new_n1194));
  NOR2_X1   g0994(.A1(new_n781), .A2(new_n218), .ZN(new_n1195));
  AOI211_X1 g0995(.A(G41), .B(new_n282), .C1(new_n840), .C2(G77), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n758), .A2(G283), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1196), .B(new_n1197), .C1(new_n216), .C2(new_n766), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1195), .B(new_n1198), .C1(new_n774), .C2(G107), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1194), .B(new_n1199), .C1(new_n1071), .C2(new_n776), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT58), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n272), .B1(new_n353), .B2(G41), .ZN(new_n1204));
  AND4_X1   g1004(.A1(new_n1192), .A2(new_n1202), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n670), .A2(new_n307), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n315), .B(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n315), .A2(new_n1206), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n315), .A2(new_n1206), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1211), .A2(new_n1212), .A3(new_n1208), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1210), .A2(new_n1213), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1181), .B1(new_n862), .B2(new_n1205), .C1(new_n1214), .C2(new_n817), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT119), .ZN(new_n1216));
  OAI21_X1  g1016(.A(KEYINPUT121), .B1(new_n919), .B2(KEYINPUT120), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT120), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT121), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(new_n909), .C2(new_n918), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1217), .A2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(G330), .B1(new_n933), .B2(new_n935), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1214), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1214), .B(G330), .C1(new_n933), .C2(new_n935), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1221), .B(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1216), .B1(new_n1227), .B2(new_n805), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1081), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1147), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1153), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1128), .A2(new_n1144), .A3(KEYINPUT117), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1230), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  AND3_X1   g1033(.A1(new_n1224), .A2(new_n919), .A3(new_n1225), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n919), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1235));
  OAI21_X1  g1035(.A(KEYINPUT57), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1229), .B1(new_n1233), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT57), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1147), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1239), .B1(new_n1240), .B2(new_n1227), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1228), .B1(new_n1238), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(KEYINPUT122), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1216), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1221), .A2(new_n1226), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n1217), .A2(new_n1220), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1244), .B1(new_n1247), .B2(new_n806), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT57), .B1(new_n1233), .B2(new_n1247), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1081), .B1(new_n1240), .B2(new_n1236), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1248), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT122), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1243), .A2(new_n1253), .ZN(G375));
  NAND2_X1  g1054(.A1(new_n960), .A2(new_n371), .ZN(new_n1255));
  XOR2_X1   g1055(.A(new_n1255), .B(KEYINPUT124), .Z(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n335), .B2(new_n776), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(G116), .B2(new_n845), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1071), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n1259), .A2(new_n955), .B1(G97), .B2(new_n840), .ZN(new_n1260));
  OAI221_X1 g1060(.A(new_n1260), .B1(new_n760), .B2(new_n757), .C1(new_n843), .C2(new_n764), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(G283), .B2(new_n774), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n282), .B1(new_n762), .B2(new_n789), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(new_n767), .B2(G58), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n955), .A2(G50), .B1(new_n758), .B2(G128), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1264), .B(new_n1265), .C1(new_n857), .C2(new_n843), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(G150), .B2(new_n777), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n962), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1166), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n774), .A2(new_n1268), .B1(new_n845), .B2(new_n1269), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n1258), .A2(new_n1262), .B1(new_n1267), .B2(new_n1270), .ZN(new_n1271));
  OAI221_X1 g1071(.A(new_n807), .B1(G68), .B2(new_n1158), .C1(new_n1271), .C2(new_n862), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(new_n816), .B2(new_n1133), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(new_n1143), .B2(new_n806), .ZN(new_n1274));
  XOR2_X1   g1074(.A(new_n1040), .B(KEYINPUT123), .Z(new_n1275));
  NAND2_X1  g1075(.A1(new_n1144), .A2(new_n1275), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1274), .B1(new_n1276), .B2(new_n1277), .ZN(G381));
  AOI21_X1  g1078(.A(G378), .B1(new_n1243), .B2(new_n1253), .ZN(new_n1279));
  INV_X1    g1079(.A(G390), .ZN(new_n1280));
  INV_X1    g1080(.A(G384), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1078), .A2(new_n827), .A3(new_n1082), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1280), .A2(new_n1281), .A3(new_n1283), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1284), .A2(G387), .A3(G381), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1279), .A2(new_n1285), .ZN(G407));
  AND2_X1   g1086(.A1(new_n671), .A2(G213), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1279), .A2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(G407), .A2(new_n1288), .A3(G213), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT125), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1289), .B(new_n1290), .ZN(G409));
  OAI21_X1  g1091(.A(new_n806), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n1216), .ZN(new_n1293));
  NOR3_X1   g1093(.A1(new_n1156), .A2(new_n1293), .A3(new_n1178), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1233), .A2(new_n1247), .A3(new_n1275), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1287), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1296), .B1(new_n1242), .B2(new_n1179), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1277), .A2(KEYINPUT60), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1149), .A2(new_n1229), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT60), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1300), .B1(new_n1230), .B2(new_n1143), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1298), .A2(new_n1299), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1274), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1281), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1302), .A2(G384), .A3(new_n1274), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1287), .A2(G2897), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1304), .A2(new_n1305), .A3(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1306), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT61), .B1(new_n1297), .B2(new_n1309), .ZN(new_n1310));
  AND2_X1   g1110(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1296), .B(new_n1311), .C1(new_n1242), .C2(new_n1179), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT63), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1310), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1251), .A2(G378), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1316), .A2(KEYINPUT63), .A3(new_n1311), .A4(new_n1296), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(G387), .A2(new_n1280), .ZN(new_n1318));
  XNOR2_X1  g1118(.A(G393), .B(new_n827), .ZN(new_n1319));
  OAI211_X1 g1119(.A(G390), .B(new_n986), .C1(new_n1019), .C2(new_n1042), .ZN(new_n1320));
  AND3_X1   g1120(.A1(new_n1318), .A2(new_n1319), .A3(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1319), .B1(new_n1318), .B2(new_n1320), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1317), .A2(new_n1323), .ZN(new_n1324));
  OAI21_X1  g1124(.A(KEYINPUT126), .B1(new_n1315), .B2(new_n1324), .ZN(new_n1325));
  AND2_X1   g1125(.A1(new_n1317), .A2(new_n1323), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT126), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1326), .A2(new_n1327), .A3(new_n1314), .A4(new_n1310), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1325), .A2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT62), .ZN(new_n1330));
  AND2_X1   g1130(.A1(new_n1312), .A2(new_n1330), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1312), .A2(new_n1330), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1310), .B1(new_n1331), .B2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT127), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(new_n1323), .B(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1333), .A2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1329), .A2(new_n1336), .ZN(G405));
  INV_X1    g1137(.A(new_n1311), .ZN(new_n1338));
  OAI211_X1 g1138(.A(new_n1338), .B(new_n1316), .C1(G375), .C2(G378), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1316), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1311), .B1(new_n1279), .B2(new_n1340), .ZN(new_n1341));
  AND3_X1   g1141(.A1(new_n1339), .A2(new_n1341), .A3(new_n1323), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1323), .B1(new_n1339), .B2(new_n1341), .ZN(new_n1343));
  NOR2_X1   g1143(.A1(new_n1342), .A2(new_n1343), .ZN(G402));
endmodule


