//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 1 0 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1327, new_n1328;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  INV_X1    g0005(.A(G87), .ZN(new_n206));
  INV_X1    g0006(.A(G250), .ZN(new_n207));
  INV_X1    g0007(.A(G97), .ZN(new_n208));
  INV_X1    g0008(.A(G257), .ZN(new_n209));
  OAI22_X1  g0009(.A1(new_n206), .A2(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AOI21_X1  g0010(.A(new_n210), .B1(G68), .B2(G238), .ZN(new_n211));
  INV_X1    g0011(.A(G107), .ZN(new_n212));
  INV_X1    g0012(.A(G264), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n214), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G77), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AND2_X1   g0020(.A1(G58), .A2(G232), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n205), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n205), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  AOI211_X1 g0025(.A(new_n207), .B(new_n225), .C1(new_n209), .C2(new_n213), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n226), .A2(KEYINPUT0), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(KEYINPUT0), .ZN(new_n228));
  NOR2_X1   g0028(.A1(G58), .A2(G68), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT64), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  INV_X1    g0033(.A(G20), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g0036(.A1(new_n227), .A2(new_n228), .A3(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n237), .B(KEYINPUT65), .Z(new_n238));
  NOR2_X1   g0038(.A1(new_n223), .A2(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n213), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G270), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G358));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n250), .B(new_n253), .Z(G351));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n255), .B1(G41), .B2(G45), .ZN(new_n256));
  OR2_X1    g0056(.A1(new_n256), .A2(KEYINPUT66), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(KEYINPUT66), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  OAI211_X1 g0060(.A(G1), .B(G13), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n257), .A2(G274), .A3(new_n258), .A4(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n256), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(new_n217), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT3), .B(G33), .ZN(new_n266));
  INV_X1    g0066(.A(G1698), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(G222), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(G1698), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT67), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n269), .B(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G223), .ZN(new_n272));
  OAI221_X1 g0072(.A(new_n268), .B1(new_n218), .B2(new_n266), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n274));
  AOI211_X1 g0074(.A(new_n263), .B(new_n265), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G190), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT70), .B(G200), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n277), .B1(new_n278), .B2(new_n275), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT71), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n233), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n255), .A2(G20), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G50), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n255), .A2(G13), .A3(G20), .ZN(new_n288));
  OAI21_X1  g0088(.A(G20), .B1(new_n230), .B2(G50), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n234), .A2(new_n259), .A3(KEYINPUT69), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT69), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n291), .B1(G20), .B2(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G150), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n289), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n259), .A2(G20), .ZN(new_n297));
  NOR2_X1   g0097(.A1(KEYINPUT8), .A2(G58), .ZN(new_n298));
  NAND2_X1  g0098(.A1(KEYINPUT68), .A2(G58), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(KEYINPUT68), .A2(G58), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n298), .B1(new_n302), .B2(KEYINPUT8), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n296), .B1(new_n297), .B2(new_n303), .ZN(new_n304));
  OAI221_X1 g0104(.A(new_n287), .B1(G50), .B2(new_n288), .C1(new_n304), .C2(new_n283), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT9), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n275), .A2(new_n276), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n275), .A2(new_n278), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT10), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n280), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n279), .B(new_n306), .C1(KEYINPUT71), .C2(KEYINPUT10), .ZN(new_n312));
  AND2_X1   g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AND2_X1   g0113(.A1(KEYINPUT3), .A2(G33), .ZN(new_n314));
  NOR2_X1   g0114(.A1(KEYINPUT3), .A2(G33), .ZN(new_n315));
  OAI211_X1 g0115(.A(G226), .B(new_n267), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  OAI211_X1 g0116(.A(G232), .B(G1698), .C1(new_n314), .C2(new_n315), .ZN(new_n317));
  NAND2_X1  g0117(.A1(G33), .A2(G97), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n274), .ZN(new_n320));
  INV_X1    g0120(.A(new_n264), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G238), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n262), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT13), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT13), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n320), .A2(new_n325), .A3(new_n322), .A4(new_n262), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n324), .A2(KEYINPUT72), .A3(new_n326), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n320), .A2(new_n322), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT72), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n328), .A2(new_n329), .A3(new_n325), .A4(new_n262), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n327), .A2(G169), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT14), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT14), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n327), .A2(new_n333), .A3(G169), .A4(new_n330), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n324), .A2(G179), .A3(new_n326), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G68), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G20), .ZN(new_n338));
  INV_X1    g0138(.A(G13), .ZN(new_n339));
  NOR3_X1   g0139(.A1(new_n338), .A2(G1), .A3(new_n339), .ZN(new_n340));
  XOR2_X1   g0140(.A(new_n340), .B(KEYINPUT12), .Z(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(new_n337), .B2(new_n285), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT73), .B1(new_n294), .B2(new_n216), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n297), .A2(G77), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT73), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n293), .A2(new_n345), .A3(G50), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n343), .A2(new_n338), .A3(new_n344), .A4(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n282), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT11), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT11), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n347), .A2(new_n350), .A3(new_n282), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n342), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n336), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n327), .A2(G200), .A3(new_n330), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n324), .A2(G190), .A3(new_n326), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n356), .A2(new_n352), .A3(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G179), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n275), .A2(new_n360), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n361), .B(new_n305), .C1(G169), .C2(new_n275), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n314), .A2(new_n315), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(G107), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n266), .A2(G232), .A3(new_n267), .ZN(new_n365));
  INV_X1    g0165(.A(G238), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n364), .B(new_n365), .C1(new_n271), .C2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n274), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n264), .A2(new_n219), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n262), .A3(new_n370), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n371), .A2(new_n278), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n288), .A2(G77), .ZN(new_n373));
  XOR2_X1   g0173(.A(KEYINPUT15), .B(G87), .Z(new_n374));
  AOI22_X1  g0174(.A1(new_n374), .A2(new_n297), .B1(G20), .B2(G77), .ZN(new_n375));
  XOR2_X1   g0175(.A(KEYINPUT8), .B(G58), .Z(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n293), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n283), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  AOI211_X1 g0178(.A(new_n373), .B(new_n378), .C1(G77), .C2(new_n286), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(new_n371), .B2(new_n276), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n372), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n313), .A2(new_n359), .A3(new_n362), .A4(new_n382), .ZN(new_n383));
  NOR3_X1   g0183(.A1(new_n300), .A2(new_n301), .A3(new_n337), .ZN(new_n384));
  OAI21_X1  g0184(.A(G20), .B1(new_n384), .B2(new_n229), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT75), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT74), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n293), .B2(G159), .ZN(new_n388));
  INV_X1    g0188(.A(G159), .ZN(new_n389));
  AOI211_X1 g0189(.A(KEYINPUT74), .B(new_n389), .C1(new_n290), .C2(new_n292), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n385), .B(new_n386), .C1(new_n388), .C2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT16), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n385), .B1(new_n388), .B2(new_n390), .ZN(new_n393));
  OR2_X1    g0193(.A1(KEYINPUT3), .A2(G33), .ZN(new_n394));
  NAND2_X1  g0194(.A1(KEYINPUT3), .A2(G33), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(new_n234), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n394), .A2(KEYINPUT7), .A3(new_n234), .A4(new_n395), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n337), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n391), .B(new_n392), .C1(new_n393), .C2(new_n400), .ZN(new_n401));
  OR2_X1    g0201(.A1(KEYINPUT68), .A2(G58), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n402), .A2(G68), .A3(new_n299), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n234), .B1(new_n403), .B2(new_n230), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n291), .A2(G20), .A3(G33), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT69), .B1(new_n234), .B2(new_n259), .ZN(new_n406));
  OAI21_X1  g0206(.A(G159), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT74), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n293), .A2(new_n387), .A3(G159), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n404), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n400), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n410), .B(new_n411), .C1(new_n386), .C2(KEYINPUT16), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n401), .A2(new_n412), .A3(new_n282), .ZN(new_n413));
  INV_X1    g0213(.A(G200), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n272), .A2(new_n267), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n217), .A2(G1698), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n415), .B(new_n416), .C1(new_n314), .C2(new_n315), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G33), .A2(G87), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n417), .A2(KEYINPUT76), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT76), .B1(new_n417), .B2(new_n418), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n419), .A2(new_n420), .A3(new_n261), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n321), .A2(G232), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n262), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n414), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n422), .A2(new_n262), .ZN(new_n425));
  INV_X1    g0225(.A(new_n420), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n417), .A2(KEYINPUT76), .A3(new_n418), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n426), .A2(new_n274), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n425), .A2(new_n428), .A3(new_n276), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n424), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT77), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n303), .A2(new_n288), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n286), .B2(new_n303), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n413), .A2(new_n430), .A3(new_n431), .A4(new_n433), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n434), .B(KEYINPUT17), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n413), .A2(new_n433), .ZN(new_n436));
  OAI21_X1  g0236(.A(G169), .B1(new_n421), .B2(new_n423), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n425), .A2(new_n428), .A3(G179), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT18), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n436), .A2(KEYINPUT18), .A3(new_n439), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n368), .A2(new_n360), .A3(new_n262), .A4(new_n370), .ZN(new_n445));
  INV_X1    g0245(.A(new_n379), .ZN(new_n446));
  AOI211_X1 g0246(.A(new_n263), .B(new_n369), .C1(new_n367), .C2(new_n274), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n445), .B(new_n446), .C1(new_n447), .C2(G169), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n435), .A2(new_n444), .A3(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n383), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n266), .A2(KEYINPUT4), .A3(G244), .A4(new_n267), .ZN(new_n451));
  OAI21_X1  g0251(.A(G244), .B1(new_n314), .B2(new_n315), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT4), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G283), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n451), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n266), .A2(G250), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n267), .B1(new_n457), .B2(KEYINPUT4), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n274), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n255), .A2(G45), .ZN(new_n460));
  OR2_X1    g0260(.A1(KEYINPUT5), .A2(G41), .ZN(new_n461));
  NAND2_X1  g0261(.A1(KEYINPUT5), .A2(G41), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT79), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(new_n464), .A3(G274), .ZN(new_n465));
  INV_X1    g0265(.A(G45), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(G1), .ZN(new_n467));
  NOR2_X1   g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  AND2_X1   g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n467), .B(G274), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT79), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n467), .B1(new_n469), .B2(new_n468), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n261), .ZN(new_n474));
  OAI21_X1  g0274(.A(KEYINPUT80), .B1(new_n474), .B2(new_n209), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT80), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n473), .A2(new_n476), .A3(G257), .A4(new_n261), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n459), .A2(new_n472), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(G169), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n288), .A2(G97), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n259), .A2(G1), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n283), .B1(KEYINPUT78), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(KEYINPUT78), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n288), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G97), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n212), .B1(new_n398), .B2(new_n399), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n294), .A2(new_n218), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT6), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n208), .A2(new_n212), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n492), .B1(new_n493), .B2(new_n202), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n212), .A2(KEYINPUT6), .A3(G97), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n234), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n490), .A2(new_n491), .A3(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n483), .B(new_n489), .C1(new_n497), .C2(new_n283), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n207), .B1(new_n394), .B2(new_n395), .ZN(new_n499));
  OAI21_X1  g0299(.A(G1698), .B1(new_n499), .B2(new_n453), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n452), .A2(new_n453), .B1(G33), .B2(G283), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n500), .A2(new_n501), .A3(new_n451), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n502), .A2(new_n274), .B1(new_n465), .B2(new_n471), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n503), .A2(new_n360), .A3(new_n478), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n481), .A2(new_n498), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT81), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n481), .A2(new_n498), .A3(new_n504), .A4(KEYINPUT81), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OR3_X1    g0309(.A1(new_n466), .A2(G1), .A3(G274), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n460), .A2(new_n207), .ZN(new_n511));
  AND3_X1   g0311(.A1(new_n510), .A2(new_n261), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G116), .ZN(new_n513));
  OAI22_X1  g0313(.A1(new_n314), .A2(new_n315), .B1(G244), .B2(new_n267), .ZN(new_n514));
  NOR2_X1   g0314(.A1(G238), .A2(G1698), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n512), .B1(new_n274), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n278), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(G190), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n266), .A2(new_n234), .A3(G68), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n318), .A2(new_n234), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n522), .B(KEYINPUT19), .C1(new_n203), .C2(G87), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n318), .A2(G20), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n521), .B(new_n523), .C1(KEYINPUT19), .C2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n288), .ZN(new_n526));
  INV_X1    g0326(.A(new_n374), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n525), .A2(new_n282), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n488), .A2(G87), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n519), .A2(new_n520), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n488), .A2(new_n374), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n518), .A2(new_n480), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n517), .A2(new_n360), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n479), .A2(new_n276), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n414), .B1(new_n503), .B2(new_n478), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n498), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n509), .A2(new_n536), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(KEYINPUT23), .B1(new_n234), .B2(G107), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT23), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n544), .A2(new_n212), .A3(G20), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT85), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n513), .B2(G20), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n234), .A2(KEYINPUT85), .A3(G33), .A4(G116), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n546), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n234), .B(G87), .C1(new_n314), .C2(new_n315), .ZN(new_n551));
  XOR2_X1   g0351(.A(KEYINPUT84), .B(KEYINPUT22), .Z(new_n552));
  AND2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n551), .A2(new_n552), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n550), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT86), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(KEYINPUT86), .B(new_n550), .C1(new_n553), .C2(new_n554), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n558), .A3(KEYINPUT24), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT24), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n555), .A2(new_n556), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n282), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n488), .A2(G107), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n526), .B(new_n212), .C1(KEYINPUT87), .C2(KEYINPUT25), .ZN(new_n564));
  NAND2_X1  g0364(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n565));
  XNOR2_X1  g0365(.A(new_n564), .B(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n562), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  OAI22_X1  g0367(.A1(new_n314), .A2(new_n315), .B1(G250), .B2(G1698), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n267), .A2(G257), .ZN(new_n569));
  INV_X1    g0369(.A(G294), .ZN(new_n570));
  OAI22_X1  g0370(.A1(new_n568), .A2(new_n569), .B1(new_n259), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n463), .A2(new_n274), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n274), .A2(new_n571), .B1(new_n572), .B2(G264), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n573), .A2(new_n472), .ZN(new_n574));
  OAI21_X1  g0374(.A(KEYINPUT88), .B1(new_n574), .B2(new_n480), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(G179), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n573), .A2(new_n472), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT88), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n577), .A2(new_n578), .A3(G169), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n575), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n567), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n577), .A2(new_n276), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n577), .A2(G200), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n562), .A2(new_n563), .A3(new_n566), .A4(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n581), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n267), .A2(G257), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n266), .B(new_n586), .C1(new_n213), .C2(new_n267), .ZN(new_n587));
  INV_X1    g0387(.A(G303), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n363), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n274), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n473), .A2(G270), .A3(new_n261), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n472), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT82), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n472), .A2(KEYINPUT82), .A3(new_n592), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n591), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G190), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n455), .B(new_n234), .C1(G33), .C2(new_n208), .ZN(new_n599));
  INV_X1    g0399(.A(G116), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(G20), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n282), .A3(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT20), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n603), .A2(KEYINPUT83), .ZN(new_n604));
  OR2_X1    g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n602), .A2(new_n604), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n605), .A2(new_n606), .B1(KEYINPUT83), .B2(new_n603), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(G116), .B1(new_n485), .B2(new_n487), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n288), .A2(new_n600), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n598), .B(new_n613), .C1(new_n414), .C2(new_n597), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n597), .A2(new_n612), .A3(G179), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n595), .A2(new_n596), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n590), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n480), .B1(new_n608), .B2(new_n611), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n617), .A2(new_n618), .A3(KEYINPUT21), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT21), .ZN(new_n620));
  INV_X1    g0420(.A(new_n611), .ZN(new_n621));
  OAI21_X1  g0421(.A(G169), .B1(new_n621), .B2(new_n607), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n620), .B1(new_n622), .B2(new_n597), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n614), .A2(new_n615), .A3(new_n619), .A4(new_n623), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n542), .A2(new_n585), .A3(new_n624), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n450), .A2(new_n625), .ZN(G372));
  INV_X1    g0426(.A(new_n362), .ZN(new_n627));
  INV_X1    g0427(.A(new_n358), .ZN(new_n628));
  INV_X1    g0428(.A(new_n448), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n355), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT17), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n434), .B(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n444), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n627), .B1(new_n633), .B2(new_n313), .ZN(new_n634));
  INV_X1    g0434(.A(new_n450), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n507), .A2(new_n536), .A3(new_n508), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT26), .ZN(new_n637));
  INV_X1    g0437(.A(new_n505), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(new_n536), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n637), .A2(new_n535), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT90), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n535), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n644), .B1(new_n636), .B2(KEYINPUT26), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n645), .A2(KEYINPUT90), .A3(new_n640), .ZN(new_n646));
  INV_X1    g0446(.A(new_n581), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n619), .A2(new_n623), .A3(new_n615), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n647), .A2(KEYINPUT89), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT89), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n619), .A2(new_n623), .A3(new_n615), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n650), .B1(new_n651), .B2(new_n581), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n582), .ZN(new_n654));
  INV_X1    g0454(.A(new_n584), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n542), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n643), .A2(new_n646), .B1(new_n653), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n634), .B1(new_n635), .B2(new_n657), .ZN(G369));
  NAND3_X1  g0458(.A1(new_n255), .A2(new_n234), .A3(G13), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(G213), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT91), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(G343), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n567), .A2(new_n665), .ZN(new_n666));
  OAI22_X1  g0466(.A1(new_n585), .A2(new_n666), .B1(new_n581), .B2(new_n664), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n613), .A2(new_n664), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n648), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n624), .B2(new_n668), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n670), .A2(KEYINPUT92), .A3(G330), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT92), .B1(new_n670), .B2(G330), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n667), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT93), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n673), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n671), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n678), .A2(KEYINPUT93), .A3(new_n667), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n651), .A2(new_n665), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n655), .A2(new_n654), .B1(new_n567), .B2(new_n580), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n647), .A2(new_n664), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n680), .A2(new_n685), .ZN(G399));
  INV_X1    g0486(.A(KEYINPUT94), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n225), .B2(G41), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n224), .A2(KEYINPUT94), .A3(new_n260), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n202), .A2(new_n206), .A3(new_n600), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n691), .A2(new_n255), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n693), .B1(new_n232), .B2(new_n691), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n694), .B(KEYINPUT28), .Z(new_n695));
  INV_X1    g0495(.A(KEYINPUT96), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n643), .A2(new_n646), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n651), .A2(new_n581), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(KEYINPUT89), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n655), .A2(new_n654), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n530), .A2(new_n535), .ZN(new_n701));
  AOI221_X4 g0501(.A(new_n701), .B1(new_n539), .B2(new_n540), .C1(new_n507), .C2(new_n508), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n651), .A2(new_n650), .A3(new_n581), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n699), .A2(new_n700), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n665), .B1(new_n697), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n696), .B1(new_n705), .B2(KEYINPUT29), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n702), .A2(new_n700), .A3(new_n698), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n636), .A2(new_n639), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n638), .A2(new_n536), .A3(KEYINPUT26), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT98), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n638), .A2(new_n536), .A3(KEYINPUT98), .A4(KEYINPUT26), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n708), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  XOR2_X1   g0513(.A(new_n535), .B(KEYINPUT97), .Z(new_n714));
  NAND3_X1  g0514(.A1(new_n707), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n715), .A2(KEYINPUT29), .A3(new_n664), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT29), .ZN(new_n717));
  OAI211_X1 g0517(.A(KEYINPUT96), .B(new_n717), .C1(new_n657), .C2(new_n665), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n706), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n614), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n648), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n702), .A2(new_n682), .A3(new_n721), .A4(new_n664), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n573), .A2(KEYINPUT95), .A3(new_n517), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n616), .A2(G179), .A3(new_n590), .A4(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(KEYINPUT95), .B1(new_n573), .B2(new_n517), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n479), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n723), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(G179), .B1(new_n616), .B2(new_n590), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n729), .A2(new_n577), .A3(new_n518), .A4(new_n479), .ZN(new_n730));
  AOI211_X1 g0530(.A(new_n360), .B(new_n591), .C1(new_n595), .C2(new_n596), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n479), .A2(new_n726), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n731), .A2(KEYINPUT30), .A3(new_n732), .A4(new_n724), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n728), .A2(new_n730), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n665), .ZN(new_n735));
  AOI21_X1  g0535(.A(KEYINPUT31), .B1(new_n734), .B2(new_n665), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n722), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G330), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n719), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n695), .B1(new_n740), .B2(G1), .ZN(G364));
  NOR2_X1   g0541(.A1(new_n339), .A2(G20), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n255), .B1(new_n742), .B2(G45), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n691), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n670), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G13), .A2(G33), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n746), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n233), .B1(G20), .B2(new_n480), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n234), .A2(G179), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n278), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n276), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n206), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT100), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n234), .A2(new_n360), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n758), .B1(new_n760), .B2(new_n414), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n759), .A2(KEYINPUT100), .A3(G200), .ZN(new_n762));
  AND3_X1   g0562(.A1(new_n761), .A2(G190), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n757), .B1(G50), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n761), .A2(new_n276), .A3(new_n762), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n754), .A2(G190), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n764), .B1(new_n337), .B2(new_n765), .C1(new_n212), .C2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G190), .A2(G200), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n759), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n363), .B1(new_n770), .B2(G77), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n276), .A2(G179), .A3(G200), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n234), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n760), .A2(new_n276), .A3(G200), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n302), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n771), .B1(new_n208), .B2(new_n773), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n753), .A2(new_n769), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G159), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT32), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n768), .A2(new_n777), .A3(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n765), .ZN(new_n783));
  XNOR2_X1  g0583(.A(KEYINPUT33), .B(G317), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n783), .A2(new_n784), .B1(new_n766), .B2(G283), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(new_n588), .B2(new_n756), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n763), .A2(G326), .B1(G329), .B2(new_n779), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n266), .B1(new_n774), .B2(G322), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n773), .A2(new_n570), .ZN(new_n790));
  INV_X1    g0590(.A(new_n770), .ZN(new_n791));
  INV_X1    g0591(.A(G311), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR4_X1   g0593(.A1(new_n786), .A2(new_n789), .A3(new_n790), .A4(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n752), .B1(new_n782), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n750), .A2(new_n752), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n225), .A2(new_n266), .ZN(new_n798));
  INV_X1    g0598(.A(new_n232), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n799), .B2(G45), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n250), .A2(new_n466), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n800), .A2(new_n801), .B1(G116), .B2(new_n224), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n225), .A2(new_n363), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n802), .B1(G355), .B2(new_n803), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n751), .B(new_n795), .C1(new_n797), .C2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G330), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n747), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n745), .B1(new_n808), .B2(KEYINPUT99), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n677), .B(new_n671), .C1(new_n808), .C2(KEYINPUT99), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n805), .B1(new_n810), .B2(new_n811), .ZN(G396));
  AOI22_X1  g0612(.A1(new_n763), .A2(G303), .B1(G116), .B2(new_n770), .ZN(new_n813));
  INV_X1    g0613(.A(G283), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n814), .B2(new_n765), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT101), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n775), .A2(new_n570), .B1(new_n208), .B2(new_n773), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT102), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n206), .A2(new_n767), .B1(new_n756), .B2(new_n212), .ZN(new_n819));
  NOR3_X1   g0619(.A1(new_n818), .A2(new_n266), .A3(new_n819), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n816), .B(new_n820), .C1(new_n792), .C2(new_n778), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n783), .A2(G150), .B1(G143), .B2(new_n774), .ZN(new_n822));
  INV_X1    g0622(.A(G137), .ZN(new_n823));
  INV_X1    g0623(.A(new_n763), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n822), .B1(new_n823), .B2(new_n824), .C1(new_n389), .C2(new_n791), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT34), .Z(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(G50), .B2(new_n755), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n363), .B1(new_n779), .B2(G132), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n766), .A2(G68), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n776), .A2(new_n773), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n821), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT103), .Z(new_n833));
  AOI21_X1  g0633(.A(new_n746), .B1(new_n833), .B2(new_n752), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n752), .A2(new_n748), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n448), .A2(new_n665), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n372), .A2(new_n380), .B1(new_n379), .B2(new_n664), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n837), .B1(new_n838), .B2(new_n448), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n834), .B1(G77), .B2(new_n836), .C1(new_n749), .C2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n839), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n705), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(new_n739), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n746), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n840), .A2(new_n844), .ZN(G384));
  INV_X1    g0645(.A(KEYINPUT38), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n437), .A2(new_n438), .ZN(new_n847));
  INV_X1    g0647(.A(new_n663), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n847), .A2(new_n848), .B1(new_n413), .B2(new_n433), .ZN(new_n849));
  AND3_X1   g0649(.A1(new_n413), .A2(new_n430), .A3(new_n433), .ZN(new_n850));
  OAI21_X1  g0650(.A(KEYINPUT37), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AND3_X1   g0651(.A1(new_n401), .A2(new_n412), .A3(new_n282), .ZN(new_n852));
  INV_X1    g0652(.A(new_n433), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n852), .A2(new_n853), .B1(new_n439), .B2(new_n663), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT37), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n413), .A2(new_n430), .A3(new_n433), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n851), .A2(new_n857), .A3(KEYINPUT106), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT106), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n854), .A2(new_n859), .A3(new_n855), .A4(new_n856), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n436), .A2(new_n663), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n435), .B2(new_n444), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n846), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n392), .B1(new_n393), .B2(new_n400), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT16), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n865), .A2(new_n866), .A3(new_n282), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT105), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n867), .A2(new_n868), .A3(new_n433), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n868), .B1(new_n867), .B2(new_n433), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI221_X4 g0671(.A(new_n441), .B1(new_n437), .B2(new_n438), .C1(new_n413), .C2(new_n433), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT18), .B1(new_n436), .B2(new_n439), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n663), .B(new_n871), .C1(new_n632), .C2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n439), .A2(new_n663), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n869), .A2(new_n876), .A3(new_n870), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT37), .B1(new_n877), .B2(new_n850), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n857), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n875), .A2(new_n879), .A3(KEYINPUT38), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n864), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT39), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n875), .A2(new_n879), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n846), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n885), .A2(KEYINPUT39), .A3(new_n880), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n354), .A2(new_n665), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n352), .A2(new_n664), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n891), .B(new_n358), .C1(new_n336), .C2(new_n353), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n354), .A2(new_n664), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n641), .A2(new_n642), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT90), .B1(new_n645), .B2(new_n640), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n704), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(new_n664), .A3(new_n839), .ZN(new_n898));
  INV_X1    g0698(.A(new_n837), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n894), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n885), .A2(new_n880), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n874), .A2(new_n848), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n890), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n706), .A2(new_n450), .A3(new_n718), .A4(new_n716), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n634), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n904), .B(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n839), .B1(new_n892), .B2(new_n893), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n735), .A2(KEYINPUT107), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT107), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n734), .A2(new_n911), .A3(KEYINPUT31), .A4(new_n665), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n722), .A2(new_n910), .A3(new_n737), .A4(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n881), .A2(new_n909), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT40), .B1(new_n885), .B2(new_n880), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n736), .B1(new_n625), .B2(new_n664), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n910), .A2(new_n912), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n908), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI22_X1  g0718(.A1(KEYINPUT40), .A2(new_n914), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(new_n916), .B2(new_n917), .ZN(new_n920));
  INV_X1    g0720(.A(new_n919), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(G330), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n450), .A2(G330), .A3(new_n913), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n920), .A2(new_n450), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n907), .B(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n255), .B2(new_n742), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n494), .A2(new_n495), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n927), .B(KEYINPUT104), .Z(new_n928));
  AOI21_X1  g0728(.A(new_n600), .B1(new_n928), .B2(KEYINPUT35), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n929), .B(new_n235), .C1(KEYINPUT35), .C2(new_n928), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT36), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n232), .A2(G77), .A3(new_n403), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(G50), .B2(new_n337), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n933), .A2(G1), .A3(new_n339), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n926), .A2(new_n931), .A3(new_n934), .ZN(G367));
  INV_X1    g0735(.A(G317), .ZN(new_n936));
  OAI221_X1 g0736(.A(new_n363), .B1(new_n778), .B2(new_n936), .C1(new_n791), .C2(new_n814), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n766), .A2(G97), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n938), .B1(new_n570), .B2(new_n765), .C1(new_n824), .C2(new_n792), .ZN(new_n939));
  OAI21_X1  g0739(.A(KEYINPUT46), .B1(new_n756), .B2(new_n600), .ZN(new_n940));
  OR3_X1    g0740(.A1(new_n756), .A2(KEYINPUT46), .A3(new_n600), .ZN(new_n941));
  AOI211_X1 g0741(.A(new_n937), .B(new_n939), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  OAI221_X1 g0742(.A(new_n942), .B1(new_n212), .B2(new_n773), .C1(new_n588), .C2(new_n775), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT109), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n778), .A2(new_n823), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n767), .A2(new_n218), .ZN(new_n946));
  INV_X1    g0746(.A(new_n773), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n783), .A2(G159), .B1(G68), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n216), .B2(new_n791), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n946), .B(new_n949), .C1(new_n302), .C2(new_n755), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n363), .B1(new_n763), .B2(G143), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n950), .B(new_n951), .C1(new_n295), .C2(new_n775), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n944), .B1(new_n945), .B2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT47), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n752), .ZN(new_n955));
  INV_X1    g0755(.A(new_n798), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n796), .B1(new_n224), .B2(new_n527), .C1(new_n246), .C2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n528), .A2(new_n529), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n665), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n536), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n644), .A2(new_n958), .A3(new_n665), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n960), .A2(new_n750), .A3(new_n961), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n955), .A2(new_n745), .A3(new_n957), .A4(new_n962), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n509), .A2(new_n541), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n665), .A2(new_n498), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n638), .A2(new_n665), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(KEYINPUT44), .B1(new_n685), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n683), .A2(new_n684), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n964), .A2(new_n965), .B1(new_n638), .B2(new_n665), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT44), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(KEYINPUT45), .B1(new_n685), .B2(new_n968), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT45), .ZN(new_n975));
  NOR3_X1   g0775(.A1(new_n970), .A2(new_n971), .A3(new_n975), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n969), .B(new_n973), .C1(new_n974), .C2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n680), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n977), .A2(new_n676), .A3(new_n679), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n667), .A2(new_n681), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n683), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT108), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n672), .B2(new_n673), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n677), .A2(KEYINPUT108), .A3(new_n671), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n984), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n678), .A2(new_n983), .A3(new_n985), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n740), .B1(new_n981), .B2(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n690), .B(KEYINPUT41), .Z(new_n993));
  AOI21_X1  g0793(.A(new_n744), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n964), .A2(new_n681), .A3(new_n682), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT42), .Z(new_n996));
  OAI21_X1  g0796(.A(new_n509), .B1(new_n971), .B2(new_n581), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n664), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n960), .A2(new_n961), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n996), .A2(new_n998), .B1(KEYINPUT43), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n680), .B2(new_n971), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n680), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1003), .A2(new_n1007), .A3(new_n968), .A4(new_n1004), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n963), .B1(new_n994), .B2(new_n1009), .ZN(G387));
  NAND3_X1  g0810(.A1(new_n719), .A2(new_n739), .A3(new_n990), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n691), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT115), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1011), .A2(KEYINPUT115), .A3(new_n691), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1014), .A2(new_n740), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n363), .B1(new_n774), .B2(G50), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n303), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n824), .A2(KEYINPUT112), .A3(new_n389), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT112), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n763), .B2(G159), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1017), .B1(new_n1018), .B2(new_n765), .C1(new_n1019), .C2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n374), .B2(new_n947), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n770), .A2(G68), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n755), .A2(G77), .B1(G150), .B2(new_n779), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1023), .A2(new_n938), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(KEYINPUT113), .B(G322), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n763), .A2(new_n1027), .B1(G303), .B2(new_n770), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n792), .B2(new_n765), .C1(new_n936), .C2(new_n775), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT48), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n814), .B2(new_n773), .C1(new_n570), .C2(new_n756), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT49), .Z(new_n1032));
  AOI21_X1  g0832(.A(new_n266), .B1(new_n779), .B2(G326), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n767), .B2(new_n600), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1026), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT114), .Z(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n752), .ZN(new_n1037));
  OR3_X1    g0837(.A1(new_n667), .A2(G20), .A3(new_n749), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n956), .B1(new_n243), .B2(G45), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(new_n692), .B2(new_n803), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n376), .A2(new_n216), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1041), .B(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n337), .A2(new_n218), .ZN(new_n1044));
  NOR4_X1   g0844(.A1(new_n1043), .A2(G45), .A3(new_n1044), .A4(new_n692), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n1040), .A2(new_n1045), .B1(G107), .B2(new_n224), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n746), .B1(new_n1046), .B2(new_n796), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT111), .Z(new_n1048));
  NAND3_X1  g0848(.A1(new_n1037), .A2(new_n1038), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n744), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1016), .B(new_n1049), .C1(new_n1050), .C2(new_n991), .ZN(G393));
  AOI21_X1  g0851(.A(new_n690), .B1(new_n981), .B2(new_n1011), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n981), .B2(new_n1011), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n981), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n752), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n763), .A2(G317), .B1(G311), .B2(new_n774), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT52), .Z(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n212), .B2(new_n767), .C1(new_n588), .C2(new_n765), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G283), .B2(new_n755), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n947), .A2(G116), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n779), .A2(new_n1027), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n266), .B1(new_n770), .B2(G294), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n266), .B1(new_n765), .B2(new_n216), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n763), .A2(G150), .B1(G159), .B2(new_n774), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT51), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1064), .B(new_n1066), .C1(G87), .C2(new_n766), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n947), .A2(G77), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n779), .A2(G143), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n755), .A2(G68), .B1(new_n376), .B2(new_n770), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1055), .B1(new_n1063), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n253), .A2(new_n798), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n797), .B1(G97), .B2(new_n225), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n746), .B(new_n1072), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n971), .A2(new_n750), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT116), .Z(new_n1077));
  AOI22_X1  g0877(.A1(new_n1054), .A2(new_n744), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1053), .A2(new_n1078), .ZN(G390));
  NOR2_X1   g0879(.A1(new_n888), .A2(new_n749), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n755), .A2(G150), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT53), .Z(new_n1082));
  AOI21_X1  g0882(.A(new_n363), .B1(new_n783), .B2(G137), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1082), .B(new_n1083), .C1(new_n389), .C2(new_n773), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G128), .B2(new_n763), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n774), .A2(G132), .ZN(new_n1086));
  XOR2_X1   g0886(.A(KEYINPUT54), .B(G143), .Z(new_n1087));
  AOI22_X1  g0887(.A1(new_n770), .A2(new_n1087), .B1(new_n779), .B2(G125), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1085), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(G50), .B2(new_n766), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n829), .B1(new_n570), .B2(new_n778), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n363), .B1(new_n1091), .B2(KEYINPUT119), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n757), .B(new_n1092), .C1(KEYINPUT119), .C2(new_n1091), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n763), .A2(G283), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n774), .A2(G116), .B1(G97), .B2(new_n770), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1093), .A2(new_n1068), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(G107), .B2(new_n783), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n752), .B1(new_n1090), .B2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1098), .B(new_n745), .C1(new_n303), .C2(new_n836), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1080), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n887), .B1(new_n900), .B2(new_n889), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n889), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n881), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n838), .A2(new_n448), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n715), .A2(new_n664), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n899), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n894), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1103), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n738), .A2(G330), .A3(new_n839), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1110), .A2(new_n894), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n1101), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n909), .A2(G330), .A3(new_n913), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n1101), .B2(new_n1109), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1100), .B1(new_n1116), .B2(new_n744), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1101), .A2(new_n1109), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1114), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n898), .A2(new_n899), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n889), .B1(new_n1121), .B2(new_n1107), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1109), .B(new_n1112), .C1(new_n1122), .C2(new_n888), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n913), .A2(KEYINPUT118), .A3(G330), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n839), .ZN(new_n1125));
  AOI21_X1  g0925(.A(KEYINPUT118), .B1(new_n913), .B2(G330), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n894), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1106), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1127), .A2(new_n1128), .A3(new_n1112), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1110), .A2(new_n894), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n1114), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1131), .A2(new_n1121), .A3(KEYINPUT117), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(KEYINPUT117), .B1(new_n1131), .B2(new_n1121), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1129), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n905), .A2(new_n923), .A3(new_n634), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1120), .A2(new_n1123), .A3(new_n1135), .A4(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n691), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n837), .B1(new_n705), .B2(new_n839), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1102), .B1(new_n1141), .B2(new_n894), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1108), .B1(new_n1142), .B2(new_n887), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1123), .B1(new_n1143), .B2(new_n1114), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1140), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1117), .B1(new_n1139), .B2(new_n1146), .ZN(G378));
  OAI21_X1  g0947(.A(new_n745), .B1(G50), .B2(new_n836), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n824), .A2(new_n600), .B1(new_n337), .B2(new_n773), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n266), .B(new_n1149), .C1(G107), .C2(new_n774), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n756), .A2(new_n218), .B1(new_n765), .B2(new_n208), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n767), .A2(new_n776), .B1(new_n814), .B2(new_n778), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1151), .A2(new_n1152), .A3(G41), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1150), .B(new_n1153), .C1(new_n527), .C2(new_n791), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT58), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(G124), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n259), .B1(new_n778), .B2(new_n1157), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n783), .A2(G132), .B1(G137), .B2(new_n770), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n763), .A2(G125), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n755), .A2(new_n1087), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(G128), .A2(new_n774), .B1(new_n947), .B2(G150), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  AOI211_X1 g0963(.A(G41), .B(new_n1158), .C1(new_n1163), .C2(KEYINPUT59), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1164), .B1(KEYINPUT59), .B2(new_n1163), .C1(new_n389), .C2(new_n767), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1166));
  AOI21_X1  g0966(.A(G50), .B1(new_n395), .B2(new_n260), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT120), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1156), .A2(new_n1165), .A3(new_n1166), .A4(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1148), .B1(new_n1169), .B2(new_n752), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n311), .A2(new_n312), .A3(new_n362), .ZN(new_n1171));
  XOR2_X1   g0971(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1172));
  OR2_X1    g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n305), .A2(new_n663), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1173), .A2(new_n305), .A3(new_n663), .A4(new_n1174), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1170), .B1(new_n1180), .B2(new_n749), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1181), .A2(KEYINPUT121), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1181), .A2(KEYINPUT121), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT122), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n919), .B2(new_n806), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n915), .A2(new_n918), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT40), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n918), .B2(new_n881), .ZN(new_n1189));
  OAI211_X1 g0989(.A(KEYINPUT122), .B(G330), .C1(new_n1187), .C2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1186), .A2(new_n1190), .A3(new_n1180), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n921), .A2(new_n1179), .A3(KEYINPUT122), .A4(G330), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1191), .A2(KEYINPUT123), .A3(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n904), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1191), .A2(KEYINPUT123), .A3(new_n904), .A4(new_n1192), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1184), .B1(new_n1197), .B2(new_n744), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n913), .A2(G330), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT118), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1201), .A2(new_n839), .A3(new_n1124), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1111), .B1(new_n1202), .B2(new_n894), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT117), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n918), .A2(G330), .B1(new_n1110), .B2(new_n894), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1204), .B1(new_n1205), .B2(new_n1141), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1128), .A2(new_n1203), .B1(new_n1206), .B2(new_n1132), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1137), .B1(new_n1144), .B2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT57), .B1(new_n1197), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n904), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1191), .A2(new_n1194), .A3(new_n1192), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1208), .A2(new_n1211), .A3(KEYINPUT57), .A4(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n691), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1198), .B1(new_n1209), .B2(new_n1214), .ZN(G375));
  AOI21_X1  g1015(.A(KEYINPUT124), .B1(new_n1207), .B2(new_n1136), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1206), .A2(new_n1132), .ZN(new_n1217));
  AND4_X1   g1017(.A1(KEYINPUT124), .A2(new_n1136), .A3(new_n1217), .A4(new_n1129), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n993), .B(new_n1140), .C1(new_n1216), .C2(new_n1218), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n766), .A2(new_n302), .B1(G50), .B2(new_n947), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n295), .B2(new_n791), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n783), .B2(new_n1087), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n779), .A2(G128), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n363), .B1(new_n755), .B2(G159), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G132), .B2(new_n763), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n823), .B2(new_n775), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n946), .B1(G107), .B2(new_n770), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n570), .B2(new_n824), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n775), .A2(new_n814), .B1(new_n527), .B2(new_n773), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n363), .B1(new_n756), .B2(new_n208), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1232), .B1(new_n600), .B2(new_n765), .C1(new_n588), .C2(new_n778), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1227), .A2(new_n1233), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n745), .B1(G68), .B2(new_n836), .C1(new_n1234), .C2(new_n1055), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n894), .B2(new_n748), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n1135), .B2(new_n744), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1219), .A2(new_n1237), .ZN(G381));
  AOI22_X1  g1038(.A1(new_n1195), .A2(new_n1196), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n691), .B(new_n1213), .C1(new_n1239), .C2(KEYINPUT57), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n1144), .A2(new_n743), .B1(new_n1080), .B2(new_n1099), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1207), .A2(new_n1136), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n690), .B1(new_n1116), .B2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1241), .B1(new_n1243), .B2(new_n1145), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1240), .A2(new_n1244), .A3(new_n1198), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(G387), .A2(G384), .A3(G390), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(G381), .A2(G393), .A3(G396), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .ZN(G407));
  OAI211_X1 g1049(.A(G407), .B(G213), .C1(G343), .C2(new_n1245), .ZN(G409));
  INV_X1    g1050(.A(G213), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1251), .A2(G343), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(G2897), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT60), .B1(new_n1207), .B2(new_n1136), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(KEYINPUT60), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1256), .A2(new_n691), .A3(new_n1258), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1259), .A2(G384), .A3(new_n1237), .ZN(new_n1260));
  AOI21_X1  g1060(.A(G384), .B1(new_n1259), .B2(new_n1237), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1254), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1259), .A2(new_n1237), .ZN(new_n1263));
  INV_X1    g1063(.A(G384), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1259), .A2(G384), .A3(new_n1237), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1265), .A2(new_n1266), .A3(new_n1253), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1244), .B1(new_n1240), .B2(new_n1198), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1197), .A2(new_n993), .A3(new_n1208), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1184), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1211), .A2(new_n744), .A3(new_n1212), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1269), .A2(new_n1244), .A3(new_n1270), .A4(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1252), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1262), .B(new_n1267), .C1(new_n1268), .C2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT61), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(KEYINPUT127), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT62), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1268), .A2(new_n1274), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1279), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(G375), .A2(G378), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1271), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(G378), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1184), .B1(new_n1239), .B2(new_n993), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1252), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  AND4_X1   g1087(.A1(new_n1279), .A2(new_n1283), .A3(new_n1281), .A4(new_n1287), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1282), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT127), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1275), .A2(new_n1290), .A3(new_n1276), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1278), .A2(new_n1289), .A3(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT125), .ZN(new_n1293));
  INV_X1    g1093(.A(G390), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1293), .B1(new_n1294), .B2(G387), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(G393), .A2(G396), .ZN(new_n1296));
  INV_X1    g1096(.A(G396), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1049), .ZN(new_n1298));
  AND3_X1   g1098(.A1(new_n1011), .A2(KEYINPUT115), .A3(new_n691), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT115), .B1(new_n1011), .B2(new_n691), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n743), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1298), .B1(new_n1301), .B2(new_n990), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1297), .B1(new_n1302), .B2(new_n1016), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1295), .B1(new_n1296), .B2(new_n1303), .ZN(new_n1304));
  XNOR2_X1  g1104(.A(G387), .B(G390), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1305), .B(new_n1295), .C1(new_n1296), .C2(new_n1303), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1292), .A2(new_n1310), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1283), .A2(new_n1281), .A3(KEYINPUT63), .A4(new_n1287), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1312), .A2(new_n1309), .A3(new_n1276), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT126), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT63), .ZN(new_n1315));
  AND2_X1   g1115(.A1(new_n1262), .A2(new_n1267), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1283), .A2(new_n1287), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1315), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1281), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1317), .A2(new_n1319), .ZN(new_n1320));
  OAI211_X1 g1120(.A(new_n1313), .B(new_n1314), .C1(new_n1318), .C2(new_n1320), .ZN(new_n1321));
  AOI22_X1  g1121(.A1(new_n1275), .A2(KEYINPUT63), .B1(new_n1281), .B2(new_n1280), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1312), .A2(new_n1309), .A3(new_n1276), .ZN(new_n1323));
  OAI21_X1  g1123(.A(KEYINPUT126), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1321), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1311), .A2(new_n1325), .ZN(G405));
  NAND2_X1  g1126(.A1(new_n1283), .A2(new_n1245), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(new_n1327), .B(new_n1319), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(new_n1328), .B(new_n1310), .ZN(G402));
endmodule


