

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749;

  NOR2_X1 U369 ( .A1(n646), .A2(n658), .ZN(n647) );
  NOR2_X1 U370 ( .A1(n659), .A2(n658), .ZN(n660) );
  AND2_X1 U371 ( .A1(n378), .A2(n377), .ZN(n374) );
  OR2_X1 U372 ( .A1(n687), .A2(n686), .ZN(n541) );
  NAND2_X1 U373 ( .A1(n471), .A2(n359), .ZN(n473) );
  BUF_X1 U374 ( .A(G104), .Z(n346) );
  XNOR2_X1 U375 ( .A(KEYINPUT66), .B(G101), .ZN(n478) );
  XNOR2_X1 U376 ( .A(KEYINPUT95), .B(G110), .ZN(n379) );
  XNOR2_X2 U377 ( .A(n382), .B(KEYINPUT0), .ZN(n532) );
  BUF_X2 U378 ( .A(n564), .Z(n608) );
  NAND2_X1 U379 ( .A1(n347), .A2(n397), .ZN(n396) );
  NAND2_X1 U380 ( .A1(n617), .A2(n361), .ZN(n347) );
  NOR2_X1 U381 ( .A1(G953), .A2(G237), .ZN(n443) );
  XNOR2_X1 U382 ( .A(G119), .B(G110), .ZN(n503) );
  NOR2_X2 U383 ( .A1(n671), .A2(n579), .ZN(n580) );
  NOR2_X2 U384 ( .A1(n672), .A2(n576), .ZN(n578) );
  OR2_X2 U385 ( .A1(n491), .A2(n357), .ZN(n492) );
  XNOR2_X2 U386 ( .A(n738), .B(n353), .ZN(n491) );
  NAND2_X1 U387 ( .A1(n677), .A2(n674), .ZN(n704) );
  XNOR2_X2 U388 ( .A(G119), .B(G116), .ZN(n410) );
  AND2_X1 U389 ( .A1(n394), .A2(n363), .ZN(n397) );
  NOR2_X1 U390 ( .A1(n381), .A2(KEYINPUT89), .ZN(n617) );
  AND2_X1 U391 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U392 ( .A(n538), .B(KEYINPUT35), .ZN(n641) );
  NAND2_X1 U393 ( .A1(n374), .A2(n373), .ZN(n630) );
  NOR2_X1 U394 ( .A1(n573), .A2(n582), .ZN(n366) );
  OR2_X1 U395 ( .A1(n649), .A2(G902), .ZN(n484) );
  XNOR2_X1 U396 ( .A(n467), .B(KEYINPUT20), .ZN(n511) );
  XNOR2_X1 U397 ( .A(KEYINPUT94), .B(KEYINPUT15), .ZN(n424) );
  XNOR2_X1 U398 ( .A(KEYINPUT16), .B(G122), .ZN(n409) );
  XNOR2_X1 U399 ( .A(G107), .B(G104), .ZN(n380) );
  XNOR2_X1 U400 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n458) );
  NAND2_X1 U401 ( .A1(n523), .A2(n687), .ZN(n348) );
  NAND2_X1 U402 ( .A1(n523), .A2(n687), .ZN(n552) );
  BUF_X1 U403 ( .A(n481), .Z(n349) );
  XNOR2_X1 U404 ( .A(n380), .B(n379), .ZN(n481) );
  BUF_X1 U405 ( .A(n736), .Z(n350) );
  XNOR2_X2 U406 ( .A(n473), .B(n472), .ZN(n523) );
  XNOR2_X1 U407 ( .A(KEYINPUT30), .B(n351), .ZN(n592) );
  NOR2_X1 U408 ( .A1(n573), .A2(n429), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n366), .B(n365), .ZN(n601) );
  XNOR2_X2 U410 ( .A(n463), .B(G134), .ZN(n477) );
  XNOR2_X1 U411 ( .A(KEYINPUT10), .B(KEYINPUT70), .ZN(n436) );
  XNOR2_X1 U412 ( .A(KEYINPUT4), .B(G137), .ZN(n474) );
  INV_X1 U413 ( .A(KEYINPUT73), .ZN(n372) );
  INV_X1 U414 ( .A(KEYINPUT48), .ZN(n368) );
  NAND2_X1 U415 ( .A1(n541), .A2(n531), .ZN(n393) );
  AND2_X1 U416 ( .A1(n390), .A2(n391), .ZN(n389) );
  OR2_X1 U417 ( .A1(n530), .A2(n392), .ZN(n391) );
  NAND2_X1 U418 ( .A1(n386), .A2(n385), .ZN(n390) );
  INV_X1 U419 ( .A(KEYINPUT102), .ZN(n439) );
  NAND2_X1 U420 ( .A1(n404), .A2(KEYINPUT36), .ZN(n403) );
  INV_X1 U421 ( .A(n407), .ZN(n404) );
  XNOR2_X1 U422 ( .A(n384), .B(n383), .ZN(n574) );
  INV_X1 U423 ( .A(KEYINPUT19), .ZN(n383) );
  INV_X1 U424 ( .A(KEYINPUT28), .ZN(n365) );
  OR2_X1 U425 ( .A1(n352), .A2(KEYINPUT109), .ZN(n377) );
  AND2_X1 U426 ( .A1(n530), .A2(n392), .ZN(n385) );
  INV_X1 U427 ( .A(G237), .ZN(n425) );
  INV_X1 U428 ( .A(KEYINPUT71), .ZN(n438) );
  NAND2_X1 U429 ( .A1(G237), .A2(G234), .ZN(n431) );
  XNOR2_X1 U430 ( .A(G113), .B(KEYINPUT76), .ZN(n411) );
  XOR2_X1 U431 ( .A(KEYINPUT85), .B(KEYINPUT23), .Z(n506) );
  XNOR2_X1 U432 ( .A(G116), .B(G107), .ZN(n454) );
  XOR2_X1 U433 ( .A(KEYINPUT105), .B(G122), .Z(n455) );
  XNOR2_X1 U434 ( .A(KEYINPUT72), .B(G140), .ZN(n499) );
  XNOR2_X1 U435 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n419) );
  INV_X1 U436 ( .A(G128), .ZN(n414) );
  XNOR2_X1 U437 ( .A(KEYINPUT86), .B(KEYINPUT4), .ZN(n416) );
  XNOR2_X1 U438 ( .A(n369), .B(n368), .ZN(n367) );
  AND2_X1 U439 ( .A1(n388), .A2(n393), .ZN(n387) );
  XOR2_X1 U440 ( .A(G143), .B(G122), .Z(n446) );
  NOR2_X1 U441 ( .A1(n457), .A2(G952), .ZN(n658) );
  OR2_X1 U442 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U443 ( .A1(n610), .A2(n674), .ZN(n595) );
  AND2_X1 U444 ( .A1(n401), .A2(n400), .ZN(n679) );
  NAND2_X1 U445 ( .A1(n520), .A2(n403), .ZN(n402) );
  OR2_X2 U446 ( .A1(n601), .A2(n575), .ZN(n672) );
  AND2_X1 U447 ( .A1(n352), .A2(KEYINPUT109), .ZN(n375) );
  AND2_X1 U448 ( .A1(n573), .A2(n517), .ZN(n352) );
  XOR2_X1 U449 ( .A(n478), .B(G146), .Z(n353) );
  AND2_X1 U450 ( .A1(n389), .A2(n393), .ZN(n354) );
  OR2_X1 U451 ( .A1(n381), .A2(n621), .ZN(n355) );
  INV_X1 U452 ( .A(n684), .ZN(n395) );
  XOR2_X1 U453 ( .A(n349), .B(n480), .Z(n356) );
  XOR2_X1 U454 ( .A(n490), .B(n489), .Z(n357) );
  NAND2_X1 U455 ( .A1(n520), .A2(n395), .ZN(n358) );
  NOR2_X1 U456 ( .A1(n702), .A2(n470), .ZN(n359) );
  AND2_X2 U457 ( .A1(n396), .A2(n355), .ZN(n653) );
  NOR2_X1 U458 ( .A1(n549), .A2(n563), .ZN(n360) );
  INV_X1 U459 ( .A(KEYINPUT36), .ZN(n408) );
  NAND2_X1 U460 ( .A1(n619), .A2(n618), .ZN(n361) );
  XOR2_X1 U461 ( .A(n604), .B(KEYINPUT91), .Z(n362) );
  AND2_X1 U462 ( .A1(n398), .A2(n620), .ZN(n363) );
  XNOR2_X1 U463 ( .A(n364), .B(n362), .ZN(n370) );
  NOR2_X1 U464 ( .A1(n748), .A2(n749), .ZN(n364) );
  NAND2_X1 U465 ( .A1(n389), .A2(n387), .ZN(n534) );
  XNOR2_X1 U466 ( .A(n491), .B(n356), .ZN(n649) );
  AND2_X2 U467 ( .A1(n367), .A2(n612), .ZN(n736) );
  NAND2_X1 U468 ( .A1(n371), .A2(n370), .ZN(n369) );
  XNOR2_X1 U469 ( .A(n586), .B(n372), .ZN(n371) );
  NAND2_X1 U470 ( .A1(n628), .A2(n630), .ZN(n527) );
  NAND2_X1 U471 ( .A1(n376), .A2(n375), .ZN(n373) );
  INV_X1 U472 ( .A(n348), .ZN(n376) );
  NAND2_X1 U473 ( .A1(n552), .A2(n518), .ZN(n378) );
  NAND2_X1 U474 ( .A1(n381), .A2(KEYINPUT89), .ZN(n394) );
  XNOR2_X1 U475 ( .A(n381), .B(KEYINPUT2), .ZN(n722) );
  NAND2_X2 U476 ( .A1(n728), .A2(n736), .ZN(n381) );
  NAND2_X1 U477 ( .A1(n574), .A2(n433), .ZN(n382) );
  NOR2_X2 U478 ( .A1(n564), .A2(n429), .ZN(n384) );
  INV_X1 U479 ( .A(n541), .ZN(n386) );
  INV_X1 U480 ( .A(n547), .ZN(n388) );
  INV_X1 U481 ( .A(n531), .ZN(n392) );
  OR2_X1 U482 ( .A1(n530), .A2(n395), .ZN(n551) );
  NAND2_X1 U483 ( .A1(n530), .A2(n360), .ZN(n581) );
  NOR2_X1 U484 ( .A1(n358), .A2(n530), .ZN(n522) );
  XNOR2_X2 U485 ( .A(n692), .B(KEYINPUT6), .ZN(n530) );
  NAND2_X1 U486 ( .A1(n361), .A2(n616), .ZN(n398) );
  OR2_X1 U487 ( .A1(n583), .A2(n408), .ZN(n400) );
  NOR2_X1 U488 ( .A1(n405), .A2(n402), .ZN(n401) );
  AND2_X1 U489 ( .A1(n583), .A2(n406), .ZN(n405) );
  AND2_X1 U490 ( .A1(n407), .A2(n408), .ZN(n406) );
  NAND2_X1 U491 ( .A1(n583), .A2(n699), .ZN(n605) );
  NOR2_X1 U492 ( .A1(n608), .A2(n429), .ZN(n407) );
  INV_X1 U493 ( .A(KEYINPUT47), .ZN(n577) );
  XNOR2_X1 U494 ( .A(n475), .B(n439), .ZN(n440) );
  INV_X1 U495 ( .A(n499), .ZN(n500) );
  XNOR2_X1 U496 ( .A(n501), .B(n500), .ZN(n737) );
  XNOR2_X1 U497 ( .A(n498), .B(G137), .ZN(n502) );
  XNOR2_X1 U498 ( .A(n502), .B(n737), .ZN(n510) );
  INV_X4 U499 ( .A(G953), .ZN(n457) );
  BUF_X1 U500 ( .A(n532), .Z(n547) );
  INV_X1 U501 ( .A(KEYINPUT123), .ZN(n625) );
  XNOR2_X1 U502 ( .A(n595), .B(KEYINPUT40), .ZN(n749) );
  XNOR2_X1 U503 ( .A(n481), .B(n409), .ZN(n413) );
  XNOR2_X1 U504 ( .A(n410), .B(KEYINPUT3), .ZN(n412) );
  XNOR2_X1 U505 ( .A(n412), .B(n411), .ZN(n489) );
  XNOR2_X1 U506 ( .A(n489), .B(n413), .ZN(n725) );
  XNOR2_X2 U507 ( .A(G143), .B(KEYINPUT88), .ZN(n415) );
  XNOR2_X2 U508 ( .A(n415), .B(n414), .ZN(n463) );
  XNOR2_X1 U509 ( .A(n478), .B(n416), .ZN(n417) );
  XNOR2_X1 U510 ( .A(n463), .B(n417), .ZN(n422) );
  XNOR2_X2 U511 ( .A(G146), .B(G125), .ZN(n437) );
  NAND2_X1 U512 ( .A1(n457), .A2(G224), .ZN(n418) );
  XNOR2_X1 U513 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U514 ( .A(n437), .B(n420), .ZN(n421) );
  XNOR2_X1 U515 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U516 ( .A(n725), .B(n423), .ZN(n655) );
  XNOR2_X1 U517 ( .A(n424), .B(G902), .ZN(n619) );
  INV_X1 U518 ( .A(n619), .ZN(n615) );
  OR2_X2 U519 ( .A1(n655), .A2(n615), .ZN(n427) );
  INV_X1 U520 ( .A(G902), .ZN(n494) );
  NAND2_X1 U521 ( .A1(n494), .A2(n425), .ZN(n428) );
  NAND2_X1 U522 ( .A1(n428), .A2(G210), .ZN(n426) );
  XNOR2_X2 U523 ( .A(n427), .B(n426), .ZN(n564) );
  NAND2_X1 U524 ( .A1(n428), .A2(G214), .ZN(n699) );
  INV_X1 U525 ( .A(n699), .ZN(n429) );
  NOR2_X1 U526 ( .A1(G898), .A2(n457), .ZN(n726) );
  NAND2_X1 U527 ( .A1(n726), .A2(G902), .ZN(n430) );
  NAND2_X1 U528 ( .A1(n457), .A2(G952), .ZN(n560) );
  NAND2_X1 U529 ( .A1(n430), .A2(n560), .ZN(n432) );
  XNOR2_X1 U530 ( .A(n431), .B(KEYINPUT14), .ZN(n682) );
  AND2_X1 U531 ( .A1(n432), .A2(n682), .ZN(n433) );
  INV_X1 U532 ( .A(n532), .ZN(n471) );
  XOR2_X1 U533 ( .A(KEYINPUT101), .B(KEYINPUT11), .Z(n435) );
  XNOR2_X1 U534 ( .A(G140), .B(KEYINPUT12), .ZN(n434) );
  XNOR2_X1 U535 ( .A(n435), .B(n434), .ZN(n442) );
  XNOR2_X1 U536 ( .A(n437), .B(n436), .ZN(n501) );
  XNOR2_X1 U537 ( .A(n438), .B(G131), .ZN(n475) );
  XNOR2_X1 U538 ( .A(n501), .B(n440), .ZN(n441) );
  XOR2_X1 U539 ( .A(n442), .B(n441), .Z(n449) );
  XOR2_X1 U540 ( .A(KEYINPUT83), .B(n443), .Z(n485) );
  NAND2_X1 U541 ( .A1(n485), .A2(G214), .ZN(n445) );
  XOR2_X1 U542 ( .A(n346), .B(G113), .Z(n444) );
  XNOR2_X1 U543 ( .A(n445), .B(n444), .ZN(n447) );
  XNOR2_X1 U544 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U545 ( .A(n449), .B(n448), .ZN(n643) );
  NAND2_X1 U546 ( .A1(n643), .A2(n494), .ZN(n453) );
  XOR2_X1 U547 ( .A(KEYINPUT13), .B(KEYINPUT104), .Z(n451) );
  XNOR2_X1 U548 ( .A(KEYINPUT103), .B(G475), .ZN(n450) );
  XNOR2_X1 U549 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X2 U550 ( .A(n453), .B(n452), .ZN(n549) );
  XNOR2_X1 U551 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U552 ( .A(n456), .B(KEYINPUT9), .Z(n462) );
  NAND2_X1 U553 ( .A1(n457), .A2(G234), .ZN(n459) );
  XNOR2_X1 U554 ( .A(n459), .B(n458), .ZN(n497) );
  NAND2_X1 U555 ( .A1(n497), .A2(G217), .ZN(n460) );
  XNOR2_X1 U556 ( .A(n460), .B(KEYINPUT7), .ZN(n461) );
  XNOR2_X1 U557 ( .A(n462), .B(n461), .ZN(n465) );
  INV_X1 U558 ( .A(n477), .ZN(n464) );
  XNOR2_X1 U559 ( .A(n465), .B(n464), .ZN(n632) );
  NAND2_X1 U560 ( .A1(n632), .A2(n494), .ZN(n466) );
  XNOR2_X1 U561 ( .A(n466), .B(G478), .ZN(n563) );
  INV_X1 U562 ( .A(n563), .ZN(n535) );
  NAND2_X1 U563 ( .A1(n549), .A2(n535), .ZN(n702) );
  NAND2_X1 U564 ( .A1(n619), .A2(G234), .ZN(n467) );
  NAND2_X1 U565 ( .A1(n511), .A2(G221), .ZN(n469) );
  INV_X1 U566 ( .A(KEYINPUT21), .ZN(n468) );
  XNOR2_X1 U567 ( .A(n469), .B(n468), .ZN(n683) );
  INV_X1 U568 ( .A(n683), .ZN(n470) );
  XNOR2_X1 U569 ( .A(KEYINPUT81), .B(KEYINPUT22), .ZN(n472) );
  XNOR2_X1 U570 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X2 U571 ( .A(n477), .B(n476), .ZN(n738) );
  AND2_X1 U572 ( .A1(n457), .A2(G227), .ZN(n479) );
  XNOR2_X1 U573 ( .A(n499), .B(n479), .ZN(n480) );
  XNOR2_X1 U574 ( .A(KEYINPUT75), .B(G469), .ZN(n482) );
  XNOR2_X1 U575 ( .A(n482), .B(KEYINPUT74), .ZN(n483) );
  XNOR2_X2 U576 ( .A(n484), .B(n483), .ZN(n568) );
  XNOR2_X2 U577 ( .A(n568), .B(KEYINPUT1), .ZN(n687) );
  NAND2_X1 U578 ( .A1(n485), .A2(G210), .ZN(n488) );
  XOR2_X1 U579 ( .A(KEYINPUT5), .B(KEYINPUT99), .Z(n486) );
  XNOR2_X1 U580 ( .A(n486), .B(KEYINPUT98), .ZN(n487) );
  XNOR2_X1 U581 ( .A(n488), .B(n487), .ZN(n490) );
  NAND2_X1 U582 ( .A1(n491), .A2(n357), .ZN(n493) );
  NAND2_X1 U583 ( .A1(n492), .A2(n493), .ZN(n635) );
  NAND2_X1 U584 ( .A1(n635), .A2(n494), .ZN(n496) );
  XOR2_X1 U585 ( .A(KEYINPUT80), .B(G472), .Z(n495) );
  XNOR2_X2 U586 ( .A(n496), .B(n495), .ZN(n521) );
  XNOR2_X2 U587 ( .A(n521), .B(KEYINPUT108), .ZN(n573) );
  NAND2_X1 U588 ( .A1(n497), .A2(G221), .ZN(n498) );
  XOR2_X1 U589 ( .A(KEYINPUT77), .B(KEYINPUT24), .Z(n504) );
  XNOR2_X1 U590 ( .A(n504), .B(n503), .ZN(n508) );
  XNOR2_X1 U591 ( .A(G128), .B(KEYINPUT96), .ZN(n505) );
  XNOR2_X1 U592 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U593 ( .A(n508), .B(n507), .Z(n509) );
  XNOR2_X1 U594 ( .A(n510), .B(n509), .ZN(n622) );
  NOR2_X1 U595 ( .A1(n622), .A2(G902), .ZN(n516) );
  XOR2_X1 U596 ( .A(KEYINPUT97), .B(KEYINPUT84), .Z(n513) );
  NAND2_X1 U597 ( .A1(n511), .A2(G217), .ZN(n512) );
  XNOR2_X1 U598 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U599 ( .A(n514), .B(KEYINPUT25), .ZN(n515) );
  XNOR2_X2 U600 ( .A(n516), .B(n515), .ZN(n571) );
  INV_X1 U601 ( .A(n571), .ZN(n517) );
  INV_X1 U602 ( .A(KEYINPUT109), .ZN(n518) );
  INV_X1 U603 ( .A(n687), .ZN(n520) );
  INV_X1 U604 ( .A(KEYINPUT107), .ZN(n519) );
  XNOR2_X1 U605 ( .A(n571), .B(n519), .ZN(n684) );
  BUF_X2 U606 ( .A(n521), .Z(n692) );
  NAND2_X1 U607 ( .A1(n523), .A2(n522), .ZN(n526) );
  INV_X1 U608 ( .A(KEYINPUT87), .ZN(n524) );
  XNOR2_X1 U609 ( .A(n524), .B(KEYINPUT32), .ZN(n525) );
  XNOR2_X1 U610 ( .A(n526), .B(n525), .ZN(n628) );
  XNOR2_X1 U611 ( .A(n527), .B(KEYINPUT92), .ZN(n539) );
  NAND2_X1 U612 ( .A1(n571), .A2(n683), .ZN(n529) );
  INV_X1 U613 ( .A(KEYINPUT67), .ZN(n528) );
  XNOR2_X2 U614 ( .A(n529), .B(n528), .ZN(n686) );
  XNOR2_X1 U615 ( .A(KEYINPUT93), .B(KEYINPUT33), .ZN(n531) );
  XNOR2_X1 U616 ( .A(KEYINPUT79), .B(KEYINPUT34), .ZN(n533) );
  XNOR2_X1 U617 ( .A(n534), .B(n533), .ZN(n537) );
  NOR2_X1 U618 ( .A1(n549), .A2(n535), .ZN(n536) );
  NAND2_X1 U619 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X2 U620 ( .A1(n539), .A2(n641), .ZN(n540) );
  XNOR2_X1 U621 ( .A(n540), .B(KEYINPUT44), .ZN(n555) );
  OR2_X1 U622 ( .A1(n541), .A2(n692), .ZN(n542) );
  XNOR2_X1 U623 ( .A(n542), .B(KEYINPUT100), .ZN(n694) );
  OR2_X1 U624 ( .A1(n694), .A2(n547), .ZN(n544) );
  INV_X1 U625 ( .A(KEYINPUT31), .ZN(n543) );
  XNOR2_X1 U626 ( .A(n544), .B(n543), .ZN(n676) );
  NOR2_X1 U627 ( .A1(n686), .A2(n568), .ZN(n545) );
  NAND2_X1 U628 ( .A1(n545), .A2(n692), .ZN(n546) );
  OR2_X1 U629 ( .A1(n547), .A2(n546), .ZN(n662) );
  NAND2_X1 U630 ( .A1(n676), .A2(n662), .ZN(n550) );
  NAND2_X1 U631 ( .A1(n563), .A2(n549), .ZN(n548) );
  XNOR2_X2 U632 ( .A(KEYINPUT106), .B(n548), .ZN(n677) );
  INV_X1 U633 ( .A(n360), .ZN(n674) );
  NAND2_X1 U634 ( .A1(n550), .A2(n704), .ZN(n553) );
  OR2_X1 U635 ( .A1(n348), .A2(n551), .ZN(n627) );
  AND2_X1 U636 ( .A1(n553), .A2(n627), .ZN(n554) );
  NAND2_X1 U637 ( .A1(n555), .A2(n554), .ZN(n557) );
  XNOR2_X1 U638 ( .A(KEYINPUT90), .B(KEYINPUT45), .ZN(n556) );
  XNOR2_X2 U639 ( .A(n557), .B(n556), .ZN(n728) );
  NOR2_X1 U640 ( .A1(G900), .A2(n457), .ZN(n558) );
  NAND2_X1 U641 ( .A1(G902), .A2(n558), .ZN(n559) );
  NAND2_X1 U642 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U643 ( .A1(n682), .A2(n561), .ZN(n587) );
  INV_X1 U644 ( .A(n587), .ZN(n562) );
  NAND2_X1 U645 ( .A1(n563), .A2(n562), .ZN(n565) );
  OR2_X1 U646 ( .A1(n565), .A2(n608), .ZN(n566) );
  OR2_X1 U647 ( .A1(n549), .A2(n566), .ZN(n567) );
  NOR2_X1 U648 ( .A1(n686), .A2(n567), .ZN(n569) );
  INV_X1 U649 ( .A(n568), .ZN(n599) );
  AND2_X1 U650 ( .A1(n569), .A2(n599), .ZN(n570) );
  AND2_X1 U651 ( .A1(n592), .A2(n570), .ZN(n671) );
  NOR2_X1 U652 ( .A1(n571), .A2(n587), .ZN(n572) );
  NAND2_X1 U653 ( .A1(n572), .A2(n683), .ZN(n582) );
  NAND2_X1 U654 ( .A1(n599), .A2(n574), .ZN(n575) );
  NAND2_X1 U655 ( .A1(n704), .A2(KEYINPUT68), .ZN(n576) );
  XNOR2_X1 U656 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U657 ( .A(n580), .B(KEYINPUT82), .ZN(n585) );
  NOR2_X1 U658 ( .A1(n582), .A2(n581), .ZN(n583) );
  INV_X1 U659 ( .A(n679), .ZN(n584) );
  OR2_X2 U660 ( .A1(n686), .A2(n587), .ZN(n589) );
  INV_X1 U661 ( .A(KEYINPUT38), .ZN(n588) );
  XNOR2_X1 U662 ( .A(n608), .B(n588), .ZN(n596) );
  NOR2_X1 U663 ( .A1(n589), .A2(n596), .ZN(n590) );
  AND2_X1 U664 ( .A1(n590), .A2(n599), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n594) );
  XOR2_X1 U666 ( .A(KEYINPUT78), .B(KEYINPUT39), .Z(n593) );
  XNOR2_X1 U667 ( .A(n594), .B(n593), .ZN(n610) );
  XOR2_X1 U668 ( .A(KEYINPUT112), .B(KEYINPUT42), .Z(n603) );
  INV_X1 U669 ( .A(n596), .ZN(n700) );
  NAND2_X1 U670 ( .A1(n700), .A2(n699), .ZN(n705) );
  NOR2_X1 U671 ( .A1(n702), .A2(n705), .ZN(n598) );
  XNOR2_X1 U672 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n597) );
  XNOR2_X1 U673 ( .A(n598), .B(n597), .ZN(n718) );
  NAND2_X1 U674 ( .A1(n718), .A2(n599), .ZN(n600) );
  XNOR2_X1 U675 ( .A(n603), .B(n602), .ZN(n748) );
  XNOR2_X1 U676 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n604) );
  XOR2_X1 U677 ( .A(n605), .B(KEYINPUT110), .Z(n606) );
  NAND2_X1 U678 ( .A1(n606), .A2(n687), .ZN(n607) );
  XNOR2_X1 U679 ( .A(n607), .B(KEYINPUT43), .ZN(n609) );
  NAND2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n629) );
  NOR2_X1 U681 ( .A1(n610), .A2(n677), .ZN(n681) );
  INV_X1 U682 ( .A(n681), .ZN(n611) );
  AND2_X1 U683 ( .A1(n629), .A2(n611), .ZN(n612) );
  INV_X1 U684 ( .A(KEYINPUT65), .ZN(n613) );
  NAND2_X1 U685 ( .A1(n613), .A2(KEYINPUT2), .ZN(n614) );
  NAND2_X1 U686 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U687 ( .A1(KEYINPUT89), .A2(KEYINPUT65), .ZN(n618) );
  INV_X1 U688 ( .A(KEYINPUT2), .ZN(n621) );
  NAND2_X1 U689 ( .A1(n621), .A2(KEYINPUT65), .ZN(n620) );
  NAND2_X1 U690 ( .A1(n653), .A2(G217), .ZN(n623) );
  XNOR2_X1 U691 ( .A(n623), .B(n622), .ZN(n624) );
  NOR2_X2 U692 ( .A1(n624), .A2(n658), .ZN(n626) );
  XNOR2_X1 U693 ( .A(n626), .B(n625), .ZN(G66) );
  XNOR2_X1 U694 ( .A(n627), .B(G101), .ZN(G3) );
  XNOR2_X1 U695 ( .A(n628), .B(G119), .ZN(G21) );
  XNOR2_X1 U696 ( .A(n629), .B(G140), .ZN(G42) );
  XNOR2_X1 U697 ( .A(n630), .B(G110), .ZN(G12) );
  AND2_X2 U698 ( .A1(n653), .A2(G478), .ZN(n631) );
  XNOR2_X1 U699 ( .A(n631), .B(n632), .ZN(n633) );
  NOR2_X1 U700 ( .A1(n633), .A2(n658), .ZN(n634) );
  XNOR2_X1 U701 ( .A(n634), .B(KEYINPUT122), .ZN(G63) );
  INV_X1 U702 ( .A(KEYINPUT63), .ZN(n640) );
  NAND2_X1 U703 ( .A1(n653), .A2(G472), .ZN(n637) );
  XOR2_X1 U704 ( .A(KEYINPUT62), .B(n635), .Z(n636) );
  XNOR2_X1 U705 ( .A(n637), .B(n636), .ZN(n638) );
  NOR2_X2 U706 ( .A1(n638), .A2(n658), .ZN(n639) );
  XNOR2_X1 U707 ( .A(n640), .B(n639), .ZN(G57) );
  XOR2_X1 U708 ( .A(n641), .B(G122), .Z(G24) );
  NAND2_X1 U709 ( .A1(n653), .A2(G475), .ZN(n645) );
  XOR2_X1 U710 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n642) );
  XNOR2_X1 U711 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U712 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U713 ( .A(n647), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U714 ( .A1(n653), .A2(G469), .ZN(n651) );
  XOR2_X1 U715 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n648) );
  XNOR2_X1 U716 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U717 ( .A(n651), .B(n650), .ZN(n652) );
  NOR2_X1 U718 ( .A1(n652), .A2(n658), .ZN(G54) );
  NAND2_X1 U719 ( .A1(n653), .A2(G210), .ZN(n657) );
  XOR2_X1 U720 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n654) );
  XNOR2_X1 U721 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U722 ( .A(n657), .B(n656), .ZN(n659) );
  XNOR2_X1 U723 ( .A(n660), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X1 U724 ( .A1(n674), .A2(n662), .ZN(n661) );
  XOR2_X1 U725 ( .A(n346), .B(n661), .Z(G6) );
  NOR2_X1 U726 ( .A1(n677), .A2(n662), .ZN(n667) );
  XOR2_X1 U727 ( .A(KEYINPUT27), .B(KEYINPUT114), .Z(n664) );
  XNOR2_X1 U728 ( .A(G107), .B(KEYINPUT113), .ZN(n663) );
  XNOR2_X1 U729 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U730 ( .A(KEYINPUT26), .B(n665), .ZN(n666) );
  XNOR2_X1 U731 ( .A(n667), .B(n666), .ZN(G9) );
  NOR2_X1 U732 ( .A1(n672), .A2(n677), .ZN(n669) );
  XNOR2_X1 U733 ( .A(KEYINPUT29), .B(KEYINPUT115), .ZN(n668) );
  XNOR2_X1 U734 ( .A(n669), .B(n668), .ZN(n670) );
  XOR2_X1 U735 ( .A(G128), .B(n670), .Z(G30) );
  XOR2_X1 U736 ( .A(G143), .B(n671), .Z(G45) );
  NOR2_X1 U737 ( .A1(n672), .A2(n674), .ZN(n673) );
  XOR2_X1 U738 ( .A(G146), .B(n673), .Z(G48) );
  NOR2_X1 U739 ( .A1(n674), .A2(n676), .ZN(n675) );
  XOR2_X1 U740 ( .A(G113), .B(n675), .Z(G15) );
  NOR2_X1 U741 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U742 ( .A(G116), .B(n678), .Z(G18) );
  XNOR2_X1 U743 ( .A(n679), .B(G125), .ZN(n680) );
  XNOR2_X1 U744 ( .A(n680), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U745 ( .A(G134), .B(n681), .Z(G36) );
  INV_X1 U746 ( .A(n682), .ZN(n716) );
  NOR2_X1 U747 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U748 ( .A(KEYINPUT49), .B(n685), .Z(n690) );
  NAND2_X1 U749 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U750 ( .A(KEYINPUT50), .B(n688), .Z(n689) );
  NOR2_X1 U751 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U752 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U753 ( .A(KEYINPUT116), .B(n693), .ZN(n695) );
  NAND2_X1 U754 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U755 ( .A(n696), .B(KEYINPUT117), .ZN(n697) );
  XNOR2_X1 U756 ( .A(n697), .B(KEYINPUT51), .ZN(n698) );
  NAND2_X1 U757 ( .A1(n698), .A2(n718), .ZN(n712) );
  NOR2_X1 U758 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U759 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U760 ( .A(KEYINPUT118), .B(n703), .Z(n709) );
  INV_X1 U761 ( .A(n704), .ZN(n706) );
  NOR2_X1 U762 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U763 ( .A(KEYINPUT119), .B(n707), .ZN(n708) );
  NAND2_X1 U764 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U765 ( .A1(n710), .A2(n354), .ZN(n711) );
  NAND2_X1 U766 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U767 ( .A(n713), .B(KEYINPUT120), .ZN(n714) );
  XOR2_X1 U768 ( .A(KEYINPUT52), .B(n714), .Z(n715) );
  NOR2_X1 U769 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U770 ( .A1(n717), .A2(G952), .ZN(n720) );
  NAND2_X1 U771 ( .A1(n718), .A2(n354), .ZN(n719) );
  NAND2_X1 U772 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U773 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U774 ( .A1(n457), .A2(n723), .ZN(n724) );
  XOR2_X1 U775 ( .A(KEYINPUT53), .B(n724), .Z(G75) );
  XOR2_X1 U776 ( .A(n725), .B(G101), .Z(n727) );
  NOR2_X1 U777 ( .A1(n727), .A2(n726), .ZN(n735) );
  NAND2_X1 U778 ( .A1(n728), .A2(n457), .ZN(n733) );
  NAND2_X1 U779 ( .A1(G224), .A2(G953), .ZN(n729) );
  XNOR2_X1 U780 ( .A(n729), .B(KEYINPUT124), .ZN(n730) );
  XNOR2_X1 U781 ( .A(KEYINPUT61), .B(n730), .ZN(n731) );
  NAND2_X1 U782 ( .A1(G898), .A2(n731), .ZN(n732) );
  NAND2_X1 U783 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U784 ( .A(n735), .B(n734), .ZN(G69) );
  XOR2_X1 U785 ( .A(n738), .B(n737), .Z(n742) );
  XNOR2_X1 U786 ( .A(n742), .B(KEYINPUT125), .ZN(n739) );
  XNOR2_X1 U787 ( .A(n350), .B(n739), .ZN(n740) );
  NAND2_X1 U788 ( .A1(n740), .A2(n457), .ZN(n747) );
  XNOR2_X1 U789 ( .A(G227), .B(KEYINPUT126), .ZN(n741) );
  XNOR2_X1 U790 ( .A(n742), .B(n741), .ZN(n743) );
  NAND2_X1 U791 ( .A1(n743), .A2(G900), .ZN(n744) );
  NAND2_X1 U792 ( .A1(n744), .A2(G953), .ZN(n745) );
  XOR2_X1 U793 ( .A(KEYINPUT127), .B(n745), .Z(n746) );
  NAND2_X1 U794 ( .A1(n747), .A2(n746), .ZN(G72) );
  XOR2_X1 U795 ( .A(G137), .B(n748), .Z(G39) );
  XOR2_X1 U796 ( .A(n749), .B(G131), .Z(G33) );
endmodule

