//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 0 1 0 1 0 1 1 1 1 0 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1324, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1400, new_n1401,
    new_n1402, new_n1403, new_n1404, new_n1405, new_n1406;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G107), .ZN(new_n219));
  INV_X1    g0019(.A(G264), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n209), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT65), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT1), .ZN(new_n224));
  AND2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n223), .A2(new_n224), .ZN(new_n226));
  INV_X1    g0026(.A(KEYINPUT64), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(G1), .B2(G13), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(KEYINPUT64), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(G50), .B1(G58), .B2(G68), .ZN(new_n232));
  NOR3_X1   g0032(.A1(new_n231), .A2(new_n207), .A3(new_n232), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n209), .A2(G13), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n234), .B(G250), .C1(G257), .C2(G264), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(KEYINPUT0), .Z(new_n236));
  NOR4_X1   g0036(.A1(new_n225), .A2(new_n226), .A3(new_n233), .A4(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  INV_X1    g0038(.A(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(KEYINPUT2), .B(G226), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G264), .B(G270), .Z(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT66), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G50), .B(G68), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G58), .B(G77), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n251), .B(new_n252), .Z(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n250), .B(new_n254), .ZN(G351));
  INV_X1    g0055(.A(KEYINPUT83), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n229), .A2(KEYINPUT64), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n227), .A2(G1), .A3(G13), .ZN(new_n258));
  AOI22_X1  g0058(.A1(new_n257), .A2(new_n258), .B1(G33), .B2(G41), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT3), .B(G33), .ZN(new_n263));
  AND3_X1   g0063(.A1(new_n262), .A2(new_n263), .A3(G223), .ZN(new_n264));
  AND2_X1   g0064(.A1(G226), .A2(G1698), .ZN(new_n265));
  AND2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n268), .B1(new_n269), .B2(new_n213), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n259), .B1(new_n264), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  INV_X1    g0072(.A(G45), .ZN(new_n273));
  AOI21_X1  g0073(.A(G1), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G1), .A3(G13), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(new_n276), .A3(G274), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n276), .A2(G232), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(G200), .B1(new_n271), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n275), .B1(new_n228), .B2(new_n230), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n269), .A2(new_n213), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n284), .B1(new_n263), .B2(new_n265), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n262), .A2(new_n263), .A3(G223), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n283), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NOR3_X1   g0087(.A1(new_n287), .A2(G190), .A3(new_n280), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n256), .B1(new_n282), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT3), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n269), .ZN(new_n291));
  NAND2_X1  g0091(.A1(KEYINPUT3), .A2(G33), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n291), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT80), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n266), .A2(new_n267), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n296), .A2(KEYINPUT80), .A3(KEYINPUT7), .A4(new_n207), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n291), .A2(new_n207), .A3(new_n292), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT7), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n295), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G68), .ZN(new_n302));
  INV_X1    g0102(.A(G58), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(new_n211), .ZN(new_n304));
  OAI21_X1  g0104(.A(G20), .B1(new_n304), .B2(new_n201), .ZN(new_n305));
  NOR2_X1   g0105(.A1(G20), .A2(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G159), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n305), .A2(KEYINPUT16), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n302), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n257), .A2(new_n258), .A3(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n211), .B1(new_n300), .B2(new_n293), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n305), .A2(new_n307), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n310), .A2(new_n312), .A3(new_n316), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT8), .B(G58), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n318), .B1(new_n206), .B2(G20), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n312), .A2(KEYINPUT69), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT69), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n257), .A2(new_n258), .A3(new_n321), .A4(new_n311), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n319), .A2(new_n320), .A3(new_n322), .A4(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n323), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n318), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G190), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n271), .A2(new_n329), .A3(new_n281), .ZN(new_n330));
  INV_X1    g0130(.A(G200), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n287), .B2(new_n280), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n330), .A2(new_n332), .A3(KEYINPUT83), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n289), .A2(new_n317), .A3(new_n328), .A4(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT17), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n257), .A2(new_n258), .A3(new_n311), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT7), .B1(new_n296), .B2(new_n207), .ZN(new_n338));
  INV_X1    g0138(.A(new_n293), .ZN(new_n339));
  OAI21_X1  g0139(.A(G68), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n340), .A2(new_n305), .A3(new_n307), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n337), .B1(new_n341), .B2(new_n313), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n327), .B1(new_n342), .B2(new_n310), .ZN(new_n343));
  NOR4_X1   g0143(.A1(new_n287), .A2(KEYINPUT82), .A3(G179), .A4(new_n280), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT82), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n285), .A2(new_n286), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n280), .B1(new_n346), .B2(new_n259), .ZN(new_n347));
  INV_X1    g0147(.A(G179), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n345), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G169), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n287), .B2(new_n280), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n344), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT18), .B1(new_n343), .B2(new_n352), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n343), .A2(KEYINPUT17), .A3(new_n289), .A4(new_n333), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n271), .A2(new_n348), .A3(new_n281), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n355), .A2(new_n351), .A3(KEYINPUT82), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n347), .A2(new_n345), .A3(new_n348), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n316), .A2(new_n312), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n308), .B1(new_n301), .B2(G68), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n328), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT18), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n358), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n336), .A2(new_n353), .A3(new_n354), .A4(new_n363), .ZN(new_n364));
  XOR2_X1   g0164(.A(KEYINPUT8), .B(G58), .Z(new_n365));
  AOI22_X1  g0165(.A1(new_n365), .A2(new_n306), .B1(G20), .B2(G77), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT71), .ZN(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT15), .B(G87), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n207), .A2(G33), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  XOR2_X1   g0170(.A(KEYINPUT15), .B(G87), .Z(new_n371));
  NOR2_X1   g0171(.A1(new_n269), .A2(G20), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(KEYINPUT71), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n366), .A2(new_n370), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT72), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n323), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n206), .A2(KEYINPUT72), .A3(G13), .A4(G20), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n374), .A2(new_n312), .B1(new_n217), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n312), .B1(new_n376), .B2(new_n377), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n217), .B1(new_n206), .B2(G20), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(KEYINPUT73), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n378), .A2(new_n337), .A3(new_n382), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT73), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n380), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n263), .A2(G238), .A3(G1698), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n296), .A2(G107), .ZN(new_n390));
  OR2_X1    g0190(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n391));
  NAND2_X1  g0191(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n391), .B(new_n392), .C1(new_n266), .C2(new_n267), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n389), .B(new_n390), .C1(new_n239), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n259), .ZN(new_n395));
  INV_X1    g0195(.A(new_n277), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n276), .A2(new_n278), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n396), .B1(G244), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n350), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n395), .A2(new_n348), .A3(new_n399), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n388), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n395), .A2(G190), .A3(new_n399), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n405), .A2(new_n380), .A3(new_n387), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n400), .A2(G200), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NOR3_X1   g0208(.A1(new_n364), .A2(new_n404), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n262), .A2(G222), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G223), .A2(G1698), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(new_n263), .A3(new_n411), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n412), .B(new_n259), .C1(G77), .C2(new_n263), .ZN(new_n413));
  XOR2_X1   g0213(.A(KEYINPUT67), .B(G226), .Z(new_n414));
  AOI21_X1  g0214(.A(new_n396), .B1(new_n398), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n350), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n306), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n372), .A2(KEYINPUT70), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT70), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n369), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n418), .B1(new_n422), .B2(new_n318), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n320), .A2(new_n322), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n423), .A2(new_n424), .B1(new_n202), .B2(new_n325), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n202), .B1(new_n206), .B2(G20), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n320), .A2(new_n322), .A3(new_n323), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n413), .A2(new_n348), .A3(new_n415), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n417), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT75), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n425), .A2(KEYINPUT9), .A3(new_n427), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n413), .A2(G190), .A3(new_n415), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT9), .B1(new_n425), .B2(new_n427), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n432), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n416), .A2(G200), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NOR3_X1   g0239(.A1(new_n435), .A2(new_n432), .A3(new_n436), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT10), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n438), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT74), .ZN(new_n443));
  AOI21_X1  g0243(.A(KEYINPUT10), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n435), .A2(new_n436), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n444), .B(new_n445), .C1(new_n443), .C2(new_n442), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n431), .B1(new_n441), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n277), .B1(new_n212), .B2(new_n397), .ZN(new_n448));
  INV_X1    g0248(.A(G1698), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n239), .A2(new_n449), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n263), .A2(new_n450), .B1(G33), .B2(G97), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n262), .A2(new_n263), .A3(G226), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n448), .B1(new_n453), .B2(new_n259), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT13), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT78), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n283), .B1(new_n451), .B2(new_n452), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT78), .ZN(new_n458));
  NOR4_X1   g0258(.A1(new_n457), .A2(new_n448), .A3(new_n458), .A4(KEYINPUT13), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT13), .B1(new_n457), .B2(new_n448), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT77), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI211_X1 g0263(.A(KEYINPUT77), .B(KEYINPUT13), .C1(new_n457), .C2(new_n448), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n460), .A2(new_n465), .A3(G190), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n306), .A2(G50), .B1(G20), .B2(new_n211), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n422), .B2(new_n217), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n424), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT11), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(KEYINPUT12), .B1(new_n378), .B2(G68), .ZN(new_n472));
  INV_X1    g0272(.A(G13), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n473), .A2(KEYINPUT12), .A3(G1), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(G20), .A3(new_n211), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n211), .B1(new_n206), .B2(G20), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n472), .A2(new_n475), .B1(new_n381), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n468), .A2(new_n424), .A3(KEYINPUT11), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n471), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT79), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT79), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n471), .A2(new_n477), .A3(new_n481), .A4(new_n478), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n453), .A2(new_n259), .ZN(new_n484));
  INV_X1    g0284(.A(new_n448), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n484), .A2(new_n455), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT76), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n486), .A2(new_n461), .A3(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(KEYINPUT76), .B(KEYINPUT13), .C1(new_n457), .C2(new_n448), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(G200), .A3(new_n489), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n466), .A2(new_n483), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n483), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n488), .A2(G169), .A3(new_n489), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT14), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n460), .A2(new_n465), .A3(G179), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT14), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n488), .A2(new_n496), .A3(G169), .A4(new_n489), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n491), .B1(new_n492), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n409), .A2(new_n447), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(G97), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n207), .B1(new_n502), .B2(G33), .ZN(new_n503));
  INV_X1    g0303(.A(G283), .ZN(new_n504));
  OAI21_X1  g0304(.A(KEYINPUT85), .B1(new_n269), .B2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT85), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n506), .A2(G33), .A3(G283), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n503), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(G116), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G20), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n509), .A2(KEYINPUT20), .A3(new_n312), .A4(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT20), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n312), .A2(new_n511), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n513), .B1(new_n514), .B2(new_n508), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n510), .B1(new_n206), .B2(G33), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n378), .A2(new_n337), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n376), .A2(new_n510), .A3(new_n377), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(G303), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n296), .A2(new_n523), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n391), .A2(G257), .A3(new_n392), .ZN(new_n525));
  OAI22_X1  g0325(.A1(new_n266), .A2(new_n267), .B1(new_n220), .B2(new_n449), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n524), .B(new_n259), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT86), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n528), .A2(new_n272), .A3(KEYINPUT5), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT5), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(KEYINPUT86), .B2(G41), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n273), .A2(G1), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n533), .A2(G270), .A3(new_n276), .ZN(new_n534));
  INV_X1    g0334(.A(G274), .ZN(new_n535));
  INV_X1    g0335(.A(new_n229), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n535), .B1(new_n536), .B2(new_n275), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n537), .A2(new_n529), .A3(new_n531), .A4(new_n532), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n527), .A2(new_n534), .A3(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n522), .A2(KEYINPUT21), .A3(G169), .A4(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT21), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n520), .B1(new_n515), .B2(new_n512), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n539), .A2(G169), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n527), .A2(G179), .A3(new_n534), .A4(new_n538), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n522), .A2(new_n546), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n538), .A2(new_n534), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n548), .A2(G190), .A3(new_n527), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n539), .A2(G200), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n542), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n540), .A2(new_n544), .A3(new_n547), .A4(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n393), .A2(new_n212), .ZN(new_n553));
  OAI211_X1 g0353(.A(G244), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n269), .B2(new_n510), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n259), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n532), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n557), .A2(G250), .A3(new_n276), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n276), .A2(G274), .ZN(new_n559));
  OAI21_X1  g0359(.A(KEYINPUT88), .B1(new_n559), .B2(new_n557), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT88), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n537), .A2(new_n561), .A3(new_n532), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n558), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n556), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n350), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n263), .A2(new_n207), .A3(G68), .ZN(new_n566));
  NAND3_X1  g0366(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n207), .ZN(new_n568));
  NOR2_X1   g0368(.A1(G97), .A2(G107), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n213), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT19), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(new_n369), .B2(new_n502), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n566), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n574), .A2(new_n312), .B1(new_n379), .B2(new_n368), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n206), .A2(G33), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n320), .A2(new_n322), .A3(new_n323), .A4(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n575), .B1(new_n368), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n556), .A2(new_n563), .A3(new_n348), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n565), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n556), .A2(new_n563), .A3(G190), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n556), .A2(new_n563), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n581), .B1(new_n582), .B2(new_n331), .ZN(new_n583));
  INV_X1    g0383(.A(new_n577), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(G87), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n575), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n580), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n552), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n533), .A2(G257), .A3(new_n276), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT87), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n538), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n590), .B1(new_n538), .B2(new_n589), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n262), .A2(new_n263), .A3(KEYINPUT4), .A4(G244), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n505), .A2(new_n507), .ZN(new_n596));
  OAI211_X1 g0396(.A(G250), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT4), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n393), .B2(new_n218), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n283), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(G200), .B1(new_n594), .B2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n219), .A2(KEYINPUT84), .A3(KEYINPUT6), .A4(G97), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT84), .ZN(new_n604));
  NAND2_X1  g0404(.A1(KEYINPUT6), .A2(G97), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n604), .B1(new_n605), .B2(G107), .ZN(new_n606));
  AND2_X1   g0406(.A1(G97), .A2(G107), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(new_n569), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n603), .B(new_n606), .C1(new_n608), .C2(KEYINPUT6), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n609), .A2(G20), .B1(G77), .B2(new_n306), .ZN(new_n610));
  OAI21_X1  g0410(.A(G107), .B1(new_n338), .B2(new_n339), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n337), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n577), .A2(new_n502), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n323), .A2(G97), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n538), .A2(new_n589), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n600), .A2(new_n596), .A3(new_n595), .A4(new_n597), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n616), .B1(new_n617), .B2(new_n259), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(G190), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n602), .A2(new_n615), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n617), .A2(new_n259), .ZN(new_n621));
  INV_X1    g0421(.A(new_n616), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n350), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n609), .A2(G20), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n306), .A2(G77), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n219), .B1(new_n300), .B2(new_n293), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n312), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n613), .ZN(new_n630));
  INV_X1    g0430(.A(new_n614), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n616), .A2(KEYINPUT87), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n591), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(new_n348), .A3(new_n621), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n624), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n620), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n391), .A2(G250), .A3(new_n392), .ZN(new_n638));
  NAND2_X1  g0438(.A1(G257), .A2(G1698), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n296), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(G33), .A2(G294), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n259), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(KEYINPUT89), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT89), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n645), .B(new_n259), .C1(new_n640), .C2(new_n642), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n533), .A2(G264), .A3(new_n276), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n538), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n644), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(G169), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n643), .A2(new_n538), .A3(new_n647), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(G179), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n207), .B(G87), .C1(new_n266), .C2(new_n267), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(KEYINPUT22), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT22), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n263), .A2(new_n656), .A3(new_n207), .A4(G87), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT24), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n269), .A2(new_n510), .A3(G20), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT23), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n207), .B2(G107), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n219), .A2(KEYINPUT23), .A3(G20), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n660), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n658), .A2(new_n659), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n659), .B1(new_n658), .B2(new_n664), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n312), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n325), .A2(new_n219), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT25), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n669), .B1(new_n584), .B2(G107), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n650), .A2(new_n653), .B1(new_n667), .B2(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n667), .A2(new_n670), .ZN(new_n672));
  OAI22_X1  g0472(.A1(new_n649), .A2(G190), .B1(new_n652), .B2(G200), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  AND4_X1   g0474(.A1(new_n501), .A2(new_n588), .A3(new_n637), .A4(new_n674), .ZN(G372));
  INV_X1    g0475(.A(KEYINPUT92), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n358), .A2(new_n361), .A3(new_n362), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n362), .B1(new_n358), .B2(new_n361), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n353), .A2(KEYINPUT92), .A3(new_n363), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n466), .A2(new_n483), .A3(new_n490), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n498), .A2(new_n492), .B1(new_n682), .B2(new_n404), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n336), .A2(new_n354), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n681), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n441), .A2(new_n446), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n431), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n672), .A2(new_n673), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n564), .A2(G200), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n689), .A2(new_n581), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT90), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n585), .A2(new_n691), .A3(new_n575), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n574), .A2(new_n312), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n379), .A2(new_n368), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n577), .A2(new_n213), .ZN(new_n696));
  OAI21_X1  g0496(.A(KEYINPUT90), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n692), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n690), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n688), .A2(new_n699), .A3(new_n636), .A4(new_n620), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n540), .A2(new_n544), .A3(new_n547), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n671), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n580), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n587), .A2(new_n636), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT26), .ZN(new_n706));
  AOI21_X1  g0506(.A(G169), .B1(new_n556), .B2(new_n563), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n348), .B2(new_n582), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n690), .A2(new_n698), .B1(new_n708), .B2(new_n578), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n624), .A2(new_n632), .A3(new_n635), .ZN(new_n710));
  AOI21_X1  g0510(.A(KEYINPUT26), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT91), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n706), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI211_X1 g0513(.A(KEYINPUT91), .B(KEYINPUT26), .C1(new_n709), .C2(new_n710), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n704), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n687), .B1(new_n716), .B2(new_n500), .ZN(G369));
  NAND2_X1  g0517(.A1(new_n650), .A2(new_n653), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n667), .A2(new_n670), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n473), .A2(G1), .A3(G20), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(G213), .B1(new_n722), .B2(KEYINPUT27), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT93), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT27), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n724), .B1(new_n721), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n722), .A2(KEYINPUT93), .A3(KEYINPUT27), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n723), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G343), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n720), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n719), .A2(new_n730), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT94), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n719), .A2(KEYINPUT94), .A3(new_n730), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n734), .A2(new_n720), .A3(new_n688), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n671), .A2(new_n730), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(KEYINPUT95), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT95), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n736), .A2(new_n737), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n701), .A2(new_n729), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n731), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n542), .A2(new_n729), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n701), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(new_n552), .B2(new_n746), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G330), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n742), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n745), .A2(new_n751), .ZN(G399));
  NAND2_X1  g0552(.A1(new_n234), .A2(new_n272), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n570), .A2(G116), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n753), .A2(G1), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(new_n232), .B2(new_n753), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT28), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT29), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n715), .A2(new_n758), .A3(new_n729), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n674), .A2(new_n588), .A3(new_n637), .A4(new_n729), .ZN(new_n760));
  AND4_X1   g0560(.A1(new_n556), .A2(new_n563), .A3(new_n643), .A4(new_n647), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT96), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n545), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n548), .A2(KEYINPUT96), .A3(G179), .A4(new_n527), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n761), .A2(new_n618), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT30), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n761), .A2(new_n763), .A3(new_n764), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n618), .A2(KEYINPUT30), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n634), .A2(new_n621), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n564), .A2(new_n651), .A3(new_n348), .A4(new_n539), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n768), .A2(new_n769), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n730), .B1(new_n767), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT31), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI211_X1 g0576(.A(KEYINPUT31), .B(new_n730), .C1(new_n767), .C2(new_n773), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n760), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G330), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n699), .A2(new_n580), .ZN(new_n780));
  OAI21_X1  g0580(.A(KEYINPUT26), .B1(new_n780), .B2(new_n636), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT26), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n705), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n703), .ZN(new_n785));
  OAI21_X1  g0585(.A(KEYINPUT29), .B1(new_n785), .B2(new_n730), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n759), .A2(new_n779), .A3(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n757), .B1(new_n788), .B2(G1), .ZN(G364));
  INV_X1    g0589(.A(new_n753), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n473), .A2(G20), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n206), .B1(new_n791), .B2(G45), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n750), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(G330), .B2(new_n748), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n234), .A2(new_n263), .ZN(new_n797));
  INV_X1    g0597(.A(G355), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n797), .A2(new_n798), .B1(G116), .B2(new_n234), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n254), .A2(G45), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n234), .A2(new_n296), .ZN(new_n801));
  INV_X1    g0601(.A(new_n232), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n801), .B1(new_n273), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n799), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n231), .B1(G20), .B2(new_n350), .ZN(new_n805));
  NOR2_X1   g0605(.A1(G13), .A2(G33), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(G20), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n794), .B1(new_n804), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(G20), .A2(G179), .ZN(new_n812));
  NOR3_X1   g0612(.A1(new_n812), .A2(G190), .A3(G200), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n263), .B1(new_n814), .B2(new_n217), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n329), .A2(G179), .A3(G200), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n207), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(G97), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n207), .A2(G190), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n820), .A2(new_n348), .A3(new_n331), .ZN(new_n821));
  INV_X1    g0621(.A(G159), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  XOR2_X1   g0624(.A(KEYINPUT99), .B(KEYINPUT32), .Z(new_n825));
  OAI21_X1  g0625(.A(new_n819), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n815), .B(new_n826), .C1(new_n824), .C2(new_n825), .ZN(new_n827));
  OR3_X1    g0627(.A1(new_n812), .A2(new_n331), .A3(KEYINPUT98), .ZN(new_n828));
  OAI21_X1  g0628(.A(KEYINPUT98), .B1(new_n812), .B2(new_n331), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(new_n329), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n828), .A2(new_n329), .A3(new_n829), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n827), .B1(new_n202), .B2(new_n832), .C1(new_n211), .C2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT100), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n331), .B2(G179), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n207), .A2(new_n329), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n348), .A2(KEYINPUT100), .A3(G200), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(G87), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n836), .A2(new_n838), .A3(new_n820), .ZN(new_n842));
  NOR3_X1   g0642(.A1(new_n812), .A2(new_n329), .A3(G200), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT97), .Z(new_n844));
  OAI221_X1 g0644(.A(new_n841), .B1(new_n219), .B2(new_n842), .C1(new_n844), .C2(new_n303), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n831), .B(KEYINPUT101), .Z(new_n846));
  INV_X1    g0646(.A(G326), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(G311), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n814), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n843), .ZN(new_n851));
  INV_X1    g0651(.A(G322), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n296), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n821), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n850), .B(new_n853), .C1(G329), .C2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n833), .ZN(new_n856));
  XNOR2_X1  g0656(.A(KEYINPUT33), .B(G317), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n818), .A2(G294), .ZN(new_n859));
  INV_X1    g0659(.A(new_n842), .ZN(new_n860));
  AOI22_X1  g0660(.A1(G303), .A2(new_n840), .B1(new_n860), .B2(G283), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n855), .A2(new_n858), .A3(new_n859), .A4(new_n861), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n834), .A2(new_n845), .B1(new_n848), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n811), .B1(new_n863), .B2(new_n805), .ZN(new_n864));
  INV_X1    g0664(.A(new_n808), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n864), .B1(new_n748), .B2(new_n865), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n796), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(G396));
  NAND2_X1  g0668(.A1(new_n403), .A2(KEYINPUT102), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT102), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n388), .A2(new_n401), .A3(new_n870), .A4(new_n402), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT103), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n729), .B1(new_n380), .B2(new_n387), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(new_n406), .B2(new_n407), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n875), .A2(new_n869), .A3(new_n871), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT103), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n730), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n715), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n716), .A2(new_n730), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n404), .A2(new_n730), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n876), .A2(new_n878), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n880), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n794), .B1(new_n884), .B2(new_n779), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n779), .B2(new_n884), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n805), .A2(new_n806), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n790), .B(new_n793), .C1(new_n887), .C2(new_n217), .ZN(new_n888));
  OAI22_X1  g0688(.A1(new_n832), .A2(new_n523), .B1(new_n504), .B2(new_n833), .ZN(new_n889));
  AOI22_X1  g0689(.A1(G107), .A2(new_n840), .B1(new_n860), .B2(G87), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n263), .B1(G294), .B2(new_n843), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n854), .A2(G311), .B1(new_n813), .B2(G116), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n890), .A2(new_n819), .A3(new_n891), .A4(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n844), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n895), .A2(G143), .B1(G159), .B2(new_n813), .ZN(new_n896));
  INV_X1    g0696(.A(G137), .ZN(new_n897));
  INV_X1    g0697(.A(G150), .ZN(new_n898));
  OAI221_X1 g0698(.A(new_n896), .B1(new_n897), .B2(new_n832), .C1(new_n898), .C2(new_n833), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT34), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n842), .A2(new_n211), .ZN(new_n901));
  INV_X1    g0701(.A(G132), .ZN(new_n902));
  OAI221_X1 g0702(.A(new_n263), .B1(new_n821), .B2(new_n902), .C1(new_n817), .C2(new_n303), .ZN(new_n903));
  AOI211_X1 g0703(.A(new_n901), .B(new_n903), .C1(G50), .C2(new_n840), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n894), .B1(new_n900), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n805), .ZN(new_n906));
  OAI221_X1 g0706(.A(new_n888), .B1(new_n883), .B2(new_n807), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n886), .A2(new_n907), .ZN(G384));
  NOR2_X1   g0708(.A1(new_n791), .A2(new_n206), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT108), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n760), .A2(new_n777), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n643), .A2(new_n647), .ZN(new_n912));
  AND4_X1   g0712(.A1(new_n582), .A2(new_n763), .A3(new_n764), .A4(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n769), .ZN(new_n914));
  INV_X1    g0714(.A(new_n772), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n913), .A2(new_n914), .B1(new_n915), .B2(new_n770), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n765), .A2(new_n766), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n729), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT107), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT31), .B1(new_n774), .B2(KEYINPUT107), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n911), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n498), .A2(new_n492), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n492), .A2(new_n730), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n923), .A2(new_n682), .A3(new_n924), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n492), .B(new_n730), .C1(new_n491), .C2(new_n498), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n883), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n910), .B1(new_n922), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n313), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n315), .B1(new_n301), .B2(G68), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n310), .B(new_n424), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n328), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n358), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n728), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n934), .A2(new_n935), .A3(new_n334), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT37), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n358), .A2(new_n361), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n361), .A2(new_n728), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT37), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n938), .A2(new_n334), .A3(new_n939), .A4(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n728), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n932), .B2(new_n328), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n937), .A2(new_n941), .B1(new_n364), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(KEYINPUT38), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n938), .A2(new_n334), .A3(new_n939), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(KEYINPUT37), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n941), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT105), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n684), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n336), .A2(new_n354), .A3(KEYINPUT105), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n681), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n939), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n949), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n945), .B1(new_n955), .B2(KEYINPUT38), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n877), .B(new_n873), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n957), .A2(new_n882), .B1(new_n925), .B2(new_n926), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n775), .B1(new_n918), .B2(new_n919), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n774), .A2(KEYINPUT107), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n777), .B(new_n760), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n958), .A2(new_n961), .A3(KEYINPUT108), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n929), .A2(new_n956), .A3(KEYINPUT40), .A4(new_n962), .ZN(new_n963));
  AND3_X1   g0763(.A1(new_n330), .A2(new_n332), .A3(KEYINPUT83), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT83), .B1(new_n330), .B2(new_n332), .ZN(new_n965));
  NOR3_X1   g0765(.A1(new_n361), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n932), .A2(new_n328), .B1(new_n356), .B2(new_n357), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n966), .A2(new_n967), .A3(new_n943), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n941), .B1(new_n968), .B2(new_n940), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n364), .A2(new_n943), .ZN(new_n970));
  AND3_X1   g0770(.A1(new_n969), .A2(KEYINPUT38), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(KEYINPUT38), .B1(new_n969), .B2(new_n970), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n958), .B(new_n961), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT40), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n963), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n501), .A2(new_n961), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(new_n977), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n978), .A2(G330), .A3(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT109), .Z(new_n981));
  NOR2_X1   g0781(.A1(new_n923), .A2(new_n730), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(KEYINPUT39), .B1(new_n971), .B2(new_n972), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n951), .A2(new_n952), .ZN(new_n985));
  NOR3_X1   g0785(.A1(new_n677), .A2(new_n678), .A3(new_n676), .ZN(new_n986));
  AOI21_X1  g0786(.A(KEYINPUT92), .B1(new_n353), .B2(new_n363), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n954), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(KEYINPUT38), .B1(new_n989), .B2(new_n948), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT39), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n945), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n984), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT106), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(KEYINPUT39), .B1(new_n944), .B2(KEYINPUT38), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n955), .B2(KEYINPUT38), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n997), .A2(KEYINPUT106), .A3(new_n984), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n983), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n872), .A2(new_n730), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(new_n715), .B2(new_n879), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n927), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n971), .A2(new_n972), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n1003), .A2(new_n1004), .B1(new_n988), .B2(new_n942), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n999), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n500), .B1(new_n759), .B2(new_n786), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n687), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1007), .B(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n909), .B1(new_n981), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n981), .B2(new_n1011), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n609), .A2(KEYINPUT35), .ZN(new_n1014));
  NOR3_X1   g0814(.A1(new_n231), .A2(new_n207), .A3(new_n510), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(KEYINPUT35), .B2(new_n609), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT104), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1014), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n1017), .B2(new_n1016), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT36), .Z(new_n1020));
  NOR3_X1   g0820(.A1(new_n304), .A2(new_n232), .A3(new_n217), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n211), .A2(G50), .ZN(new_n1022));
  OAI211_X1 g0822(.A(G1), .B(new_n473), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1013), .A2(new_n1020), .A3(new_n1023), .ZN(G367));
  OAI21_X1  g0824(.A(new_n809), .B1(new_n234), .B2(new_n368), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n245), .A2(new_n801), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n794), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n839), .A2(new_n303), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n854), .A2(G137), .B1(new_n813), .B2(G50), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n211), .B2(new_n817), .C1(new_n898), .C2(new_n851), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n1028), .B(new_n1030), .C1(G159), .C2(new_n856), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n263), .B1(new_n842), .B2(new_n217), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT115), .Z(new_n1033));
  INV_X1    g0833(.A(G143), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1031), .B(new_n1033), .C1(new_n1034), .C2(new_n846), .ZN(new_n1035));
  AOI21_X1  g0835(.A(KEYINPUT46), .B1(new_n840), .B2(G116), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT114), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n895), .A2(G303), .B1(G97), .B2(new_n860), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n856), .A2(G294), .ZN(new_n1039));
  INV_X1    g0839(.A(G317), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n296), .B1(new_n821), .B2(new_n1040), .C1(new_n814), .C2(new_n504), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G107), .B2(new_n818), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .A4(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n840), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT113), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n846), .B2(new_n849), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1035), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT47), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1027), .B1(new_n1048), .B2(new_n805), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n698), .A2(new_n729), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n709), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n1052), .A2(KEYINPUT110), .B1(new_n580), .B2(new_n1051), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(KEYINPUT110), .B2(new_n1052), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n808), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1049), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT44), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n637), .B1(new_n615), .B2(new_n729), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n710), .A2(new_n730), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1058), .B1(new_n745), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1061), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n743), .B1(new_n739), .B2(new_n741), .ZN(new_n1064));
  OAI211_X1 g0864(.A(KEYINPUT44), .B(new_n1063), .C1(new_n1064), .C2(new_n731), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n745), .A2(KEYINPUT45), .A3(new_n1061), .ZN(new_n1067));
  AND3_X1   g0867(.A1(new_n736), .A2(new_n737), .A3(new_n740), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n740), .B1(new_n736), .B2(new_n737), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n744), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n731), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1070), .A2(new_n1071), .A3(new_n1061), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT45), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1067), .A2(new_n1074), .ZN(new_n1075));
  AND3_X1   g0875(.A1(new_n1066), .A2(new_n751), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n751), .B1(new_n1066), .B2(new_n1075), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n742), .A2(new_n744), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n749), .B1(new_n1079), .B2(new_n1064), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n743), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1082), .A2(new_n750), .A3(new_n1070), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(KEYINPUT111), .B1(new_n1084), .B2(new_n787), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT111), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n788), .A2(new_n1086), .A3(new_n1083), .A4(new_n1080), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n787), .B1(new_n1078), .B2(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n753), .B(KEYINPUT41), .ZN(new_n1090));
  OAI21_X1  g0890(.A(KEYINPUT112), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1066), .A2(new_n1075), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n751), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1066), .A2(new_n751), .A3(new_n1075), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1094), .A2(new_n1087), .A3(new_n1085), .A4(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n788), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT112), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1090), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n793), .B1(new_n1091), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT43), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1054), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1064), .A2(new_n1061), .ZN(new_n1104));
  OR2_X1    g0904(.A1(new_n1104), .A2(KEYINPUT42), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n620), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n636), .B1(new_n1106), .B2(new_n720), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1104), .A2(KEYINPUT42), .B1(new_n729), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1103), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1054), .A2(new_n1102), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1109), .B(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1093), .A2(new_n1061), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1111), .B(new_n1112), .Z(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1057), .B1(new_n1101), .B2(new_n1114), .ZN(G387));
  OAI22_X1  g0915(.A1(new_n797), .A2(new_n754), .B1(G107), .B2(new_n234), .ZN(new_n1116));
  OR2_X1    g0916(.A1(new_n242), .A2(new_n273), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n754), .ZN(new_n1118));
  AOI211_X1 g0918(.A(G45), .B(new_n1118), .C1(G68), .C2(G77), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n318), .A2(G50), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT50), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n801), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1116), .B1(new_n1117), .B2(new_n1122), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n832), .A2(new_n822), .B1(new_n318), .B2(new_n833), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n817), .A2(new_n368), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n296), .B1(G50), .B2(new_n843), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1126), .B1(new_n211), .B2(new_n814), .C1(new_n898), .C2(new_n821), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n840), .A2(G77), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n502), .B2(new_n842), .ZN(new_n1129));
  NOR4_X1   g0929(.A1(new_n1124), .A2(new_n1125), .A3(new_n1127), .A4(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n296), .B1(new_n821), .B2(new_n847), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n895), .A2(G317), .B1(G303), .B2(new_n813), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n1132), .B1(new_n849), .B2(new_n833), .C1(new_n846), .C2(new_n852), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT48), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(G283), .A2(new_n818), .B1(new_n840), .B2(G294), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT49), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1131), .B(new_n1140), .C1(G116), .C2(new_n860), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1130), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n794), .B1(new_n810), .B2(new_n1123), .C1(new_n1143), .C2(new_n906), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(new_n1081), .B2(new_n808), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1084), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1145), .B1(new_n1146), .B2(new_n793), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1148), .B(new_n790), .C1(new_n788), .C2(new_n1146), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1147), .A2(new_n1149), .ZN(G393));
  OAI21_X1  g0950(.A(new_n809), .B1(new_n502), .B2(new_n234), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n249), .A2(new_n801), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n794), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n831), .A2(G317), .B1(G311), .B2(new_n843), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT52), .Z(new_n1155));
  AOI21_X1  g0955(.A(new_n263), .B1(G294), .B2(new_n813), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n852), .B2(new_n821), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(G107), .B2(new_n860), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1155), .B(new_n1158), .C1(new_n504), .C2(new_n839), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n833), .A2(new_n523), .B1(new_n510), .B2(new_n817), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1160), .B(KEYINPUT116), .Z(new_n1161));
  AOI22_X1  g0961(.A1(new_n831), .A2(G150), .B1(G159), .B2(new_n843), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT51), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n263), .B1(new_n821), .B2(new_n1034), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n817), .A2(new_n217), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1164), .B(new_n1165), .C1(new_n365), .C2(new_n813), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(G68), .A2(new_n840), .B1(new_n860), .B2(G87), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1166), .B(new_n1167), .C1(new_n202), .C2(new_n833), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n1159), .A2(new_n1161), .B1(new_n1163), .B2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1153), .B1(new_n1169), .B2(new_n805), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT117), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n865), .B2(new_n1061), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1172), .B1(new_n1173), .B2(new_n792), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT118), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n1078), .B2(new_n1088), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1173), .A2(KEYINPUT118), .A3(new_n1148), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n753), .B1(new_n1078), .B2(new_n1088), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1174), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(G390));
  INV_X1    g0981(.A(G330), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n760), .A2(new_n777), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n921), .A2(new_n920), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1182), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n778), .A2(G330), .A3(new_n883), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1185), .A2(new_n958), .B1(new_n1186), .B2(new_n1002), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n927), .B1(new_n1185), .B2(new_n883), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n879), .B1(new_n703), .B2(new_n784), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1000), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(new_n928), .C2(new_n779), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n1187), .A2(new_n1001), .B1(new_n1188), .B2(new_n1191), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n922), .A2(new_n500), .A3(new_n1182), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1008), .A2(new_n1193), .A3(new_n1009), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n983), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n995), .A2(new_n998), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n927), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1199), .A2(new_n956), .A3(new_n983), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n928), .A2(new_n779), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1197), .A2(new_n1200), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1185), .A2(new_n958), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n1197), .B2(new_n1200), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1195), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1204), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1195), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1197), .A2(new_n1200), .A3(new_n1202), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1206), .A2(new_n1212), .A3(new_n790), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n887), .ZN(new_n1214));
  INV_X1    g1014(.A(G128), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n832), .A2(new_n1215), .B1(new_n897), .B2(new_n833), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n817), .A2(new_n822), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(KEYINPUT54), .B(G143), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT119), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n1219), .A2(new_n814), .B1(new_n202), .B2(new_n842), .ZN(new_n1220));
  INV_X1    g1020(.A(G125), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n263), .B1(new_n821), .B2(new_n1221), .C1(new_n851), .C2(new_n902), .ZN(new_n1222));
  NOR4_X1   g1022(.A1(new_n1216), .A2(new_n1217), .A3(new_n1220), .A4(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n839), .A2(new_n898), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT53), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n832), .A2(new_n504), .B1(new_n219), .B2(new_n833), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n854), .A2(G294), .B1(new_n843), .B2(G116), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n502), .B2(new_n814), .ZN(new_n1228));
  NOR4_X1   g1028(.A1(new_n1226), .A2(new_n1228), .A3(new_n901), .A4(new_n1165), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n841), .A2(new_n296), .ZN(new_n1230));
  XOR2_X1   g1030(.A(new_n1230), .B(KEYINPUT120), .Z(new_n1231));
  AOI22_X1  g1031(.A1(new_n1223), .A2(new_n1225), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n794), .B1(new_n365), .B2(new_n1214), .C1(new_n1232), .C2(new_n906), .ZN(new_n1233));
  AND3_X1   g1033(.A1(new_n997), .A2(KEYINPUT106), .A3(new_n984), .ZN(new_n1234));
  AOI21_X1  g1034(.A(KEYINPUT106), .B1(new_n997), .B2(new_n984), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1233), .B1(new_n1236), .B2(new_n806), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1237), .B1(new_n1238), .B2(new_n793), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1213), .A2(new_n1239), .ZN(G378));
  AOI21_X1  g1040(.A(new_n1182), .B1(new_n973), .B2(new_n974), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n428), .A2(new_n728), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n447), .A2(new_n1242), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n447), .A2(new_n1242), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  OR3_X1    g1046(.A1(new_n1243), .A2(new_n1244), .A3(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1246), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n963), .A2(new_n1241), .A3(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1249), .B1(new_n963), .B2(new_n1241), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n1251), .A2(new_n1252), .B1(new_n999), .B2(new_n1006), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n963), .A2(new_n1241), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1249), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n982), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1256), .A2(new_n1005), .A3(new_n1257), .A4(new_n1250), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1253), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n793), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1255), .A2(new_n806), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n263), .A2(G41), .ZN(new_n1262));
  AOI211_X1 g1062(.A(G50), .B(new_n1262), .C1(new_n269), .C2(new_n272), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n371), .A2(new_n813), .B1(new_n843), .B2(G107), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n1264), .B1(new_n211), .B2(new_n817), .C1(new_n833), .C2(new_n502), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n860), .A2(G58), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n854), .A2(G283), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1128), .A2(new_n1266), .A3(new_n1262), .A4(new_n1267), .ZN(new_n1268));
  XOR2_X1   g1068(.A(new_n1268), .B(KEYINPUT121), .Z(new_n1269));
  AOI211_X1 g1069(.A(new_n1265), .B(new_n1269), .C1(G116), .C2(new_n831), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1263), .B1(new_n1270), .B2(KEYINPUT58), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(G128), .A2(new_n843), .B1(new_n813), .B2(G137), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1219), .B2(new_n839), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n831), .A2(G125), .B1(G150), .B2(new_n818), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1274), .B(KEYINPUT122), .ZN(new_n1275));
  AOI211_X1 g1075(.A(new_n1273), .B(new_n1275), .C1(G132), .C2(new_n856), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(KEYINPUT59), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n860), .A2(G159), .ZN(new_n1279));
  AOI211_X1 g1079(.A(G33), .B(G41), .C1(new_n854), .C2(G124), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1278), .A2(new_n1279), .A3(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1277), .A2(KEYINPUT59), .ZN(new_n1282));
  OAI221_X1 g1082(.A(new_n1271), .B1(KEYINPUT58), .B2(new_n1270), .C1(new_n1281), .C2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n805), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n887), .A2(new_n202), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1261), .A2(new_n794), .A3(new_n1284), .A4(new_n1285), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1260), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT57), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(new_n1253), .B2(new_n1258), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(new_n1203), .A2(new_n1205), .A3(new_n1195), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1185), .A2(new_n501), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n759), .A2(new_n786), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n687), .B(new_n1291), .C1(new_n1292), .C2(new_n500), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1289), .B1(new_n1290), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n790), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1212), .A2(new_n1194), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT57), .B1(new_n1296), .B2(new_n1259), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1287), .B1(new_n1295), .B2(new_n1297), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(new_n1298), .B(KEYINPUT123), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(G375));
  NAND2_X1  g1100(.A1(new_n1002), .A2(new_n806), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n794), .B1(new_n1214), .B2(G68), .ZN(new_n1302));
  OAI22_X1  g1102(.A1(new_n851), .A2(new_n504), .B1(new_n821), .B2(new_n523), .ZN(new_n1303));
  AOI211_X1 g1103(.A(new_n263), .B(new_n1303), .C1(G107), .C2(new_n813), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1125), .ZN(new_n1305));
  AOI22_X1  g1105(.A1(G294), .A2(new_n831), .B1(new_n856), .B2(G116), .ZN(new_n1306));
  AOI22_X1  g1106(.A1(G97), .A2(new_n840), .B1(new_n860), .B2(G77), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1304), .A2(new_n1305), .A3(new_n1306), .A4(new_n1307), .ZN(new_n1308));
  OAI221_X1 g1108(.A(new_n263), .B1(new_n821), .B2(new_n1215), .C1(new_n814), .C2(new_n898), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1309), .B1(G50), .B2(new_n818), .ZN(new_n1310));
  OAI221_X1 g1110(.A(new_n1310), .B1(new_n902), .B2(new_n832), .C1(new_n833), .C2(new_n1219), .ZN(new_n1311));
  OAI221_X1 g1111(.A(new_n1266), .B1(new_n822), .B2(new_n839), .C1(new_n844), .C2(new_n897), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1308), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1302), .B1(new_n1313), .B2(new_n805), .ZN(new_n1314));
  AOI22_X1  g1114(.A1(new_n1192), .A2(new_n793), .B1(new_n1301), .B2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1195), .A2(new_n1099), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1315), .B1(new_n1316), .B2(new_n1317), .ZN(G381));
  INV_X1    g1118(.A(G378), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(G393), .A2(G396), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(G381), .A2(G384), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1319), .A2(new_n1320), .A3(new_n1180), .A4(new_n1321), .ZN(new_n1322));
  OR3_X1    g1122(.A1(G375), .A2(G387), .A3(new_n1322), .ZN(G407));
  NAND2_X1  g1123(.A1(new_n1299), .A2(new_n1319), .ZN(new_n1324));
  OAI211_X1 g1124(.A(G407), .B(G213), .C1(G343), .C2(new_n1324), .ZN(G409));
  NAND2_X1  g1125(.A1(G387), .A2(new_n1180), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1098), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1327));
  AOI211_X1 g1127(.A(KEYINPUT112), .B(new_n1090), .C1(new_n1096), .C2(new_n788), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n792), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(new_n1113), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1330), .A2(new_n1057), .A3(G390), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1326), .A2(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n867), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1320), .A2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1332), .A2(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1326), .A2(new_n1331), .A3(new_n1334), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  OAI211_X1 g1138(.A(G378), .B(new_n1287), .C1(new_n1295), .C2(new_n1297), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1259), .A2(KEYINPUT124), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT124), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1253), .A2(new_n1258), .A3(new_n1341), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1340), .A2(new_n793), .A3(new_n1342), .ZN(new_n1343));
  OAI211_X1 g1143(.A(new_n1099), .B(new_n1259), .C1(new_n1290), .C2(new_n1293), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1343), .A2(new_n1344), .A3(new_n1286), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1345), .A2(new_n1319), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1339), .A2(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(G213), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(new_n1348), .A2(G343), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT60), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1351), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1352));
  NOR2_X1   g1152(.A1(new_n1352), .A2(new_n1317), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1001), .ZN(new_n1354));
  AND2_X1   g1154(.A1(new_n1186), .A2(new_n1002), .ZN(new_n1355));
  OAI21_X1  g1155(.A(new_n1354), .B1(new_n1208), .B2(new_n1355), .ZN(new_n1356));
  INV_X1    g1156(.A(new_n1191), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1185), .A2(new_n883), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1358), .A2(new_n1002), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1357), .A2(new_n1359), .ZN(new_n1360));
  NAND4_X1  g1160(.A1(new_n1293), .A2(new_n1356), .A3(KEYINPUT60), .A4(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1361), .A2(new_n790), .ZN(new_n1362));
  OAI21_X1  g1162(.A(new_n1315), .B1(new_n1353), .B2(new_n1362), .ZN(new_n1363));
  INV_X1    g1163(.A(G384), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1363), .A2(new_n1364), .ZN(new_n1365));
  OAI211_X1 g1165(.A(G384), .B(new_n1315), .C1(new_n1353), .C2(new_n1362), .ZN(new_n1366));
  AND2_X1   g1166(.A1(new_n1365), .A2(new_n1366), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1347), .A2(new_n1350), .A3(new_n1367), .ZN(new_n1368));
  OR2_X1    g1168(.A1(new_n1350), .A2(KEYINPUT126), .ZN(new_n1369));
  NAND3_X1  g1169(.A1(new_n1365), .A2(new_n1366), .A3(new_n1369), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1349), .A2(G2897), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1370), .A2(new_n1371), .ZN(new_n1372));
  INV_X1    g1172(.A(new_n1371), .ZN(new_n1373));
  NAND4_X1  g1173(.A1(new_n1365), .A2(new_n1366), .A3(new_n1373), .A4(new_n1369), .ZN(new_n1374));
  AND2_X1   g1174(.A1(new_n1372), .A2(new_n1374), .ZN(new_n1375));
  AOI21_X1  g1175(.A(new_n1375), .B1(new_n1347), .B2(new_n1350), .ZN(new_n1376));
  OAI21_X1  g1176(.A(new_n1368), .B1(new_n1376), .B2(KEYINPUT62), .ZN(new_n1377));
  INV_X1    g1177(.A(KEYINPUT61), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1377), .A2(new_n1378), .ZN(new_n1379));
  INV_X1    g1179(.A(KEYINPUT125), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1368), .A2(new_n1380), .ZN(new_n1381));
  AOI21_X1  g1181(.A(new_n1349), .B1(new_n1339), .B2(new_n1346), .ZN(new_n1382));
  NAND3_X1  g1182(.A1(new_n1382), .A2(KEYINPUT125), .A3(new_n1367), .ZN(new_n1383));
  AOI21_X1  g1183(.A(KEYINPUT62), .B1(new_n1381), .B2(new_n1383), .ZN(new_n1384));
  OAI21_X1  g1184(.A(new_n1338), .B1(new_n1379), .B2(new_n1384), .ZN(new_n1385));
  NAND2_X1  g1185(.A1(new_n1347), .A2(new_n1350), .ZN(new_n1386));
  INV_X1    g1186(.A(new_n1375), .ZN(new_n1387));
  AOI21_X1  g1187(.A(KEYINPUT127), .B1(new_n1386), .B2(new_n1387), .ZN(new_n1388));
  INV_X1    g1188(.A(KEYINPUT127), .ZN(new_n1389));
  NOR3_X1   g1189(.A1(new_n1382), .A2(new_n1389), .A3(new_n1375), .ZN(new_n1390));
  NOR2_X1   g1190(.A1(new_n1388), .A2(new_n1390), .ZN(new_n1391));
  INV_X1    g1191(.A(new_n1337), .ZN(new_n1392));
  AOI21_X1  g1192(.A(new_n1334), .B1(new_n1326), .B2(new_n1331), .ZN(new_n1393));
  NOR3_X1   g1193(.A1(new_n1392), .A2(new_n1393), .A3(KEYINPUT61), .ZN(new_n1394));
  INV_X1    g1194(.A(KEYINPUT63), .ZN(new_n1395));
  NAND3_X1  g1195(.A1(new_n1381), .A2(new_n1395), .A3(new_n1383), .ZN(new_n1396));
  NAND3_X1  g1196(.A1(new_n1382), .A2(KEYINPUT63), .A3(new_n1367), .ZN(new_n1397));
  NAND4_X1  g1197(.A1(new_n1391), .A2(new_n1394), .A3(new_n1396), .A4(new_n1397), .ZN(new_n1398));
  NAND2_X1  g1198(.A1(new_n1385), .A2(new_n1398), .ZN(G405));
  INV_X1    g1199(.A(new_n1367), .ZN(new_n1400));
  OAI21_X1  g1200(.A(new_n1400), .B1(new_n1392), .B2(new_n1393), .ZN(new_n1401));
  NAND2_X1  g1201(.A1(new_n1298), .A2(G378), .ZN(new_n1402));
  NAND2_X1  g1202(.A1(new_n1324), .A2(new_n1402), .ZN(new_n1403));
  NAND3_X1  g1203(.A1(new_n1336), .A2(new_n1337), .A3(new_n1367), .ZN(new_n1404));
  AND3_X1   g1204(.A1(new_n1401), .A2(new_n1403), .A3(new_n1404), .ZN(new_n1405));
  AOI21_X1  g1205(.A(new_n1403), .B1(new_n1401), .B2(new_n1404), .ZN(new_n1406));
  NOR2_X1   g1206(.A1(new_n1405), .A2(new_n1406), .ZN(G402));
endmodule


