//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n557, new_n559,
    new_n560, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1100,
    new_n1101;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  XOR2_X1   g028(.A(KEYINPUT64), .B(KEYINPUT65), .Z(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n452), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n452), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n467), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n469), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n468), .A2(new_n470), .A3(new_n471), .A4(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n463), .B(new_n466), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n469), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(new_n472), .ZN(new_n478));
  INV_X1    g053(.A(G125), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n475), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n466), .B1(new_n473), .B2(new_n474), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(KEYINPUT67), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n482), .A2(new_n484), .ZN(G160));
  INV_X1    g060(.A(new_n473), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n468), .A2(new_n470), .A3(G2105), .A4(new_n472), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT68), .B1(G100), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NOR3_X1   g067(.A1(KEYINPUT68), .A2(G100), .A3(G2105), .ZN(new_n493));
  OAI221_X1 g068(.A(G2104), .B1(G112), .B2(new_n471), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n487), .A2(new_n490), .A3(new_n494), .ZN(new_n495));
  XNOR2_X1  g070(.A(new_n495), .B(KEYINPUT69), .ZN(G162));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  OR3_X1    g072(.A1(new_n497), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(new_n478), .ZN(new_n499));
  AOI21_X1  g074(.A(KEYINPUT66), .B1(new_n469), .B2(G2104), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n469), .A2(G2104), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n502), .A2(G138), .A3(new_n471), .A4(new_n470), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n499), .B1(new_n503), .B2(KEYINPUT4), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n471), .A2(G102), .ZN(new_n506));
  NAND2_X1  g081(.A1(G114), .A2(G2105), .ZN(new_n507));
  AOI211_X1 g082(.A(new_n505), .B(new_n464), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G102), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n507), .B1(new_n509), .B2(G2105), .ZN(new_n510));
  AOI21_X1  g085(.A(KEYINPUT70), .B1(new_n510), .B2(G2104), .ZN(new_n511));
  INV_X1    g086(.A(G126), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n508), .A2(new_n511), .B1(new_n488), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n504), .A2(new_n513), .ZN(G164));
  NAND2_X1  g089(.A1(KEYINPUT71), .A2(G651), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n515), .B(new_n516), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n517), .A2(G543), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT5), .B(G543), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(G50), .A2(new_n518), .B1(new_n520), .B2(G88), .ZN(new_n521));
  XOR2_X1   g096(.A(new_n521), .B(KEYINPUT72), .Z(new_n522));
  AOI22_X1  g097(.A1(new_n519), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n522), .A2(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n517), .A2(G543), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n517), .A2(new_n519), .ZN(new_n530));
  INV_X1    g105(.A(G89), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n528), .A2(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT73), .ZN(new_n533));
  INV_X1    g108(.A(new_n519), .ZN(new_n534));
  NAND2_X1  g109(.A1(G63), .A2(G651), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n519), .A2(KEYINPUT73), .A3(G63), .A4(G651), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n532), .A2(new_n540), .ZN(G286));
  INV_X1    g116(.A(G286), .ZN(G168));
  AOI22_X1  g117(.A1(G52), .A2(new_n518), .B1(new_n520), .B2(G90), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n524), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT74), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI211_X1 g122(.A(new_n543), .B(KEYINPUT74), .C1(new_n524), .C2(new_n544), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(G171));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  INV_X1    g125(.A(G81), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n550), .A2(new_n529), .B1(new_n530), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n519), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n524), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G188));
  AND2_X1   g136(.A1(KEYINPUT75), .A2(G53), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n518), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n518), .A2(KEYINPUT9), .A3(new_n562), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n520), .A2(G91), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT76), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n519), .B(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n570), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n571), .A2(new_n524), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G299));
  INV_X1    g149(.A(G171), .ZN(G301));
  NAND2_X1  g150(.A1(new_n520), .A2(G87), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n518), .A2(G49), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(G288));
  INV_X1    g154(.A(G48), .ZN(new_n580));
  OR3_X1    g155(.A1(new_n529), .A2(KEYINPUT78), .A3(new_n580), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT78), .B1(new_n529), .B2(new_n580), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n581), .A2(new_n582), .B1(G86), .B2(new_n520), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n519), .A2(G61), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT77), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n585), .A2(new_n586), .B1(G73), .B2(G543), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n584), .A2(KEYINPUT77), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n524), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n583), .A2(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(G47), .A2(new_n518), .B1(new_n520), .B2(G85), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n524), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT79), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  XOR2_X1   g171(.A(KEYINPUT80), .B(G66), .Z(new_n597));
  AND2_X1   g172(.A1(new_n570), .A2(new_n597), .ZN(new_n598));
  AND2_X1   g173(.A1(G79), .A2(G543), .ZN(new_n599));
  OAI21_X1  g174(.A(G651), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n520), .A2(KEYINPUT10), .A3(G92), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n530), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n601), .A2(new_n604), .B1(G54), .B2(new_n518), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT81), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n596), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n596), .B1(new_n607), .B2(G868), .ZN(G321));
  MUX2_X1   g184(.A(G299), .B(G286), .S(G868), .Z(G280));
  XNOR2_X1  g185(.A(G280), .B(KEYINPUT82), .ZN(G297));
  XOR2_X1   g186(.A(KEYINPUT83), .B(G559), .Z(new_n612));
  OAI21_X1  g187(.A(new_n607), .B1(G860), .B2(new_n612), .ZN(G148));
  INV_X1    g188(.A(new_n555), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n607), .A2(new_n612), .ZN(new_n615));
  MUX2_X1   g190(.A(new_n614), .B(new_n615), .S(G868), .Z(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g192(.A1(new_n471), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2100), .ZN(new_n621));
  INV_X1    g196(.A(G123), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT84), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(new_n471), .B2(G111), .ZN(new_n624));
  OR2_X1    g199(.A1(G99), .A2(G2105), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n624), .A2(G2104), .A3(new_n625), .ZN(new_n626));
  NOR3_X1   g201(.A1(new_n623), .A2(new_n471), .A3(G111), .ZN(new_n627));
  OAI22_X1  g202(.A1(new_n488), .A2(new_n622), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(new_n486), .B2(G135), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n630), .A2(G2096), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(G2096), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n621), .A2(new_n631), .A3(new_n632), .ZN(G156));
  INV_X1    g208(.A(KEYINPUT14), .ZN(new_n634));
  XOR2_X1   g209(.A(KEYINPUT15), .B(G2435), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2427), .ZN(new_n637));
  INV_X1    g212(.A(G2430), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n634), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(new_n638), .B2(new_n637), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT85), .B(KEYINPUT16), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G1341), .B(G1348), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n640), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n640), .A2(new_n647), .ZN(new_n649));
  AND3_X1   g224(.A1(new_n648), .A2(G14), .A3(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NOR3_X1   g230(.A1(new_n652), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT18), .ZN(new_n657));
  INV_X1    g232(.A(new_n653), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT17), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n654), .B1(new_n660), .B2(new_n651), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n661), .B1(new_n652), .B2(new_n659), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n652), .A2(new_n655), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n658), .B1(new_n663), .B2(KEYINPUT17), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n657), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT86), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2096), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n667), .A2(G2100), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(G2100), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(G227));
  XOR2_X1   g245(.A(G1971), .B(G1976), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1956), .B(G2474), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1961), .B(G1966), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n673), .A2(new_n674), .ZN(new_n676));
  NOR3_X1   g251(.A1(new_n672), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n672), .A2(new_n675), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT20), .Z(new_n679));
  AOI211_X1 g254(.A(new_n677), .B(new_n679), .C1(new_n672), .C2(new_n676), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n681));
  XOR2_X1   g256(.A(new_n680), .B(new_n681), .Z(new_n682));
  XNOR2_X1  g257(.A(G1991), .B(G1996), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n682), .B(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(G229));
  NOR2_X1   g262(.A1(G16), .A2(G23), .ZN(new_n688));
  INV_X1    g263(.A(G288), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n688), .B1(new_n689), .B2(G16), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT33), .B(G1976), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT87), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n690), .B(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(G166), .A2(G16), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G16), .B2(G22), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT88), .B(G1971), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n693), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  MUX2_X1   g272(.A(G6), .B(G305), .S(G16), .Z(new_n698));
  XOR2_X1   g273(.A(KEYINPUT32), .B(G1981), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n697), .B(new_n700), .C1(new_n695), .C2(new_n696), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n701), .A2(KEYINPUT34), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(KEYINPUT34), .ZN(new_n703));
  MUX2_X1   g278(.A(G24), .B(G290), .S(G16), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(G1986), .ZN(new_n705));
  NOR2_X1   g280(.A1(G25), .A2(G29), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n486), .A2(G131), .ZN(new_n707));
  INV_X1    g282(.A(G119), .ZN(new_n708));
  AND2_X1   g283(.A1(G107), .A2(G2105), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G95), .B2(new_n471), .ZN(new_n710));
  OAI22_X1  g285(.A1(new_n488), .A2(new_n708), .B1(new_n710), .B2(new_n464), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n706), .B1(new_n712), .B2(G29), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT35), .B(G1991), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n705), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n702), .A2(new_n703), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT36), .ZN(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G21), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G168), .B2(new_n719), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT93), .B(G1966), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT94), .Z(new_n725));
  NOR2_X1   g300(.A1(G16), .A2(G19), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n555), .B2(G16), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(G1341), .Z(new_n728));
  XOR2_X1   g303(.A(KEYINPUT31), .B(G11), .Z(new_n729));
  INV_X1    g304(.A(G29), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT30), .B(G28), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n630), .B2(new_n730), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n721), .B2(new_n723), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n725), .A2(new_n728), .A3(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(G5), .A2(G16), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G171), .B2(G16), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(G1961), .ZN(new_n738));
  NAND3_X1  g313(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT26), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n739), .A2(new_n740), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n741), .A2(new_n742), .B1(G105), .B2(new_n465), .ZN(new_n743));
  INV_X1    g318(.A(G129), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n488), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n486), .B2(G141), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n746), .A2(new_n730), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n730), .B2(G32), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT27), .B(G1996), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n730), .A2(G26), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT28), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n486), .A2(G140), .ZN(new_n753));
  INV_X1    g328(.A(G128), .ZN(new_n754));
  AND2_X1   g329(.A1(G116), .A2(G2105), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G104), .B2(new_n471), .ZN(new_n756));
  OAI22_X1  g331(.A1(new_n488), .A2(new_n754), .B1(new_n756), .B2(new_n464), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n752), .B1(new_n758), .B2(new_n730), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT89), .B(G2067), .Z(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n750), .A2(new_n761), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n748), .A2(new_n749), .B1(new_n759), .B2(new_n760), .ZN(new_n763));
  INV_X1    g338(.A(G2084), .ZN(new_n764));
  NAND2_X1  g339(.A1(G160), .A2(G29), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT24), .B(G34), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(new_n730), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT92), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n762), .B(new_n763), .C1(new_n764), .C2(new_n769), .ZN(new_n770));
  NOR3_X1   g345(.A1(new_n735), .A2(new_n738), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n730), .A2(G33), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n465), .A2(G103), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT90), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT25), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n486), .A2(G139), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n477), .A2(new_n472), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n777), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n775), .B(new_n776), .C1(new_n471), .C2(new_n778), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT91), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n772), .B1(new_n780), .B2(new_n730), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(G2072), .Z(new_n782));
  NAND2_X1  g357(.A1(new_n737), .A2(G1961), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT95), .Z(new_n784));
  NAND3_X1  g359(.A1(new_n771), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n719), .A2(G20), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT23), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n573), .B2(new_n719), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(G1956), .Z(new_n789));
  NOR2_X1   g364(.A1(G27), .A2(G29), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G164), .B2(G29), .ZN(new_n791));
  INV_X1    g366(.A(G2078), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n769), .A2(new_n764), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n789), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(G29), .A2(G35), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G162), .B2(G29), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT29), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n795), .B1(G2090), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(G4), .A2(G16), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n607), .B2(G16), .ZN(new_n801));
  INV_X1    g376(.A(G1348), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n799), .B(new_n803), .C1(G2090), .C2(new_n798), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n785), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n718), .A2(new_n805), .ZN(G150));
  INV_X1    g381(.A(G150), .ZN(G311));
  NAND2_X1  g382(.A1(new_n520), .A2(G93), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT97), .B(G55), .Z(new_n810));
  OAI221_X1 g385(.A(new_n808), .B1(new_n524), .B2(new_n809), .C1(new_n529), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(G860), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT99), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT37), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n607), .A2(G559), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n811), .B(new_n555), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT39), .ZN(new_n820));
  AOI21_X1  g395(.A(G860), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n820), .B2(new_n819), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n822), .A2(KEYINPUT98), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n822), .A2(KEYINPUT98), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n814), .B1(new_n823), .B2(new_n824), .ZN(G145));
  INV_X1    g400(.A(KEYINPUT100), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n513), .A2(new_n826), .ZN(new_n827));
  OAI221_X1 g402(.A(KEYINPUT100), .B1(new_n488), .B2(new_n512), .C1(new_n508), .C2(new_n511), .ZN(new_n828));
  OAI21_X1  g403(.A(KEYINPUT4), .B1(new_n473), .B2(new_n497), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n478), .B2(new_n498), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n827), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(new_n758), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(new_n746), .ZN(new_n833));
  MUX2_X1   g408(.A(new_n780), .B(new_n779), .S(new_n833), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n712), .B(new_n619), .ZN(new_n835));
  MUX2_X1   g410(.A(G106), .B(G118), .S(G2105), .Z(new_n836));
  AOI22_X1  g411(.A1(new_n489), .A2(G130), .B1(G2104), .B2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT101), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n486), .A2(new_n838), .A3(G142), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n838), .B1(new_n486), .B2(G142), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n837), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n835), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n834), .B(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(G162), .B(G160), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n629), .ZN(new_n845));
  AOI21_X1  g420(.A(G37), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(new_n845), .B2(new_n843), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g423(.A1(new_n811), .A2(G868), .ZN(new_n849));
  OR3_X1    g424(.A1(new_n573), .A2(new_n606), .A3(KEYINPUT102), .ZN(new_n850));
  OAI21_X1  g425(.A(KEYINPUT102), .B1(new_n573), .B2(new_n606), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n573), .A2(new_n606), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(KEYINPUT41), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT41), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n852), .A2(new_n856), .A3(new_n853), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n615), .B(new_n816), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(new_n854), .B2(new_n859), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT42), .ZN(new_n862));
  XNOR2_X1  g437(.A(G303), .B(G305), .ZN(new_n863));
  XNOR2_X1  g438(.A(G288), .B(KEYINPUT103), .ZN(new_n864));
  XNOR2_X1  g439(.A(G290), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n863), .B(new_n865), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n866), .A2(KEYINPUT104), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n862), .B(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n849), .B1(new_n868), .B2(G868), .ZN(G295));
  AOI21_X1  g444(.A(new_n849), .B1(new_n868), .B2(G868), .ZN(G331));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n871));
  INV_X1    g446(.A(new_n816), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT105), .ZN(new_n873));
  NAND2_X1  g448(.A1(G171), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n547), .A2(KEYINPUT105), .A3(new_n548), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n874), .A2(G286), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(G286), .B1(new_n874), .B2(new_n875), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n872), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n874), .A2(new_n875), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(G168), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n874), .A2(G286), .A3(new_n875), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n880), .A2(new_n881), .A3(new_n816), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n878), .A2(new_n882), .A3(new_n854), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT106), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR3_X1   g460(.A1(new_n876), .A2(new_n877), .A3(new_n872), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n816), .B1(new_n880), .B2(new_n881), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n855), .B(new_n857), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n878), .A2(new_n882), .A3(KEYINPUT106), .A4(new_n854), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n885), .A2(new_n888), .A3(new_n866), .A4(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(G37), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT43), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n885), .A2(new_n888), .A3(new_n889), .ZN(new_n894));
  INV_X1    g469(.A(new_n866), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n892), .A2(new_n893), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n888), .A2(new_n883), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n895), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n899), .A2(new_n890), .A3(new_n891), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(KEYINPUT43), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n871), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT107), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n892), .A2(new_n903), .A3(new_n893), .A4(new_n899), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n899), .A2(new_n890), .A3(new_n893), .A4(new_n891), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT107), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n892), .A2(new_n896), .ZN(new_n907));
  AOI22_X1  g482(.A1(new_n904), .A2(new_n906), .B1(new_n907), .B2(KEYINPUT43), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n902), .B1(new_n908), .B2(new_n871), .ZN(G397));
  INV_X1    g484(.A(G1384), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n831), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT45), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n484), .A2(G40), .A3(new_n475), .A4(new_n481), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n746), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(G1996), .A3(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT109), .ZN(new_n918));
  INV_X1    g493(.A(G2067), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n758), .B(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n915), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n915), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n922), .A2(G1996), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n918), .B(new_n921), .C1(new_n916), .C2(new_n923), .ZN(new_n924));
  XOR2_X1   g499(.A(new_n712), .B(new_n714), .Z(new_n925));
  AOI21_X1  g500(.A(new_n924), .B1(new_n915), .B2(new_n925), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n922), .A2(G1986), .A3(G290), .ZN(new_n927));
  XOR2_X1   g502(.A(new_n927), .B(KEYINPUT48), .Z(new_n928));
  AND2_X1   g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT126), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n923), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n932), .B1(KEYINPUT126), .B2(KEYINPUT46), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n923), .A2(new_n930), .A3(new_n931), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n915), .B1(new_n916), .B2(new_n920), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  XOR2_X1   g511(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n937));
  XOR2_X1   g512(.A(new_n936), .B(new_n937), .Z(new_n938));
  NAND2_X1  g513(.A1(new_n758), .A2(new_n919), .ZN(new_n939));
  OR3_X1    g514(.A1(new_n707), .A2(new_n711), .A3(new_n714), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n939), .B1(new_n924), .B2(new_n940), .ZN(new_n941));
  AOI211_X1 g516(.A(new_n929), .B(new_n938), .C1(new_n915), .C2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n910), .B1(new_n504), .B2(new_n513), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n914), .B1(new_n943), .B2(new_n912), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n831), .A2(KEYINPUT45), .A3(new_n910), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  XOR2_X1   g521(.A(KEYINPUT110), .B(G1971), .Z(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT111), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n914), .B1(new_n943), .B2(KEYINPUT50), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT50), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n831), .A2(new_n952), .A3(new_n910), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n950), .B1(G2090), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT112), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n949), .A2(KEYINPUT111), .ZN(new_n957));
  OR3_X1    g532(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n956), .B1(new_n955), .B2(new_n957), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(new_n959), .A3(G8), .ZN(new_n960));
  NAND2_X1  g535(.A1(G303), .A2(G8), .ZN(new_n961));
  XOR2_X1   g536(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n962));
  XOR2_X1   g537(.A(new_n961), .B(new_n962), .Z(new_n963));
  NAND2_X1  g538(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(G160), .A2(G40), .A3(new_n910), .A4(new_n831), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(G8), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n966), .B1(G1976), .B2(new_n689), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT52), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n967), .B(new_n968), .C1(G1976), .C2(new_n689), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT114), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n970), .A2(KEYINPUT49), .ZN(new_n971));
  NAND2_X1  g546(.A1(G305), .A2(G1981), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G1981), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n583), .A2(new_n590), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n971), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n972), .B(new_n975), .C1(new_n970), .C2(KEYINPUT49), .ZN(new_n978));
  INV_X1    g553(.A(new_n966), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n969), .B(new_n980), .C1(new_n968), .C2(new_n967), .ZN(new_n981));
  INV_X1    g556(.A(new_n513), .ZN(new_n982));
  AOI21_X1  g557(.A(G1384), .B1(new_n830), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n914), .B1(new_n983), .B2(KEYINPUT45), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n913), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n722), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n951), .A2(new_n953), .A3(new_n764), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n988), .A2(G8), .A3(G168), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n981), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n964), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n960), .A2(new_n963), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT63), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(G288), .A2(G1976), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n976), .B1(new_n980), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT115), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n979), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n997), .B1(new_n996), .B2(new_n995), .ZN(new_n998));
  INV_X1    g573(.A(new_n981), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n998), .B1(new_n992), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n993), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1002), .B1(new_n946), .B2(G2078), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n913), .A2(KEYINPUT53), .A3(new_n984), .A4(new_n792), .ZN(new_n1004));
  INV_X1    g579(.A(G1961), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n954), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1003), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(G171), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n1008), .B(KEYINPUT121), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n988), .A2(G8), .A3(G286), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT118), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n723), .B1(new_n913), .B2(new_n984), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n951), .A2(new_n953), .A3(new_n764), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1012), .B(G8), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(G286), .A2(G8), .ZN(new_n1016));
  XOR2_X1   g591(.A(new_n1016), .B(KEYINPUT119), .Z(new_n1017));
  AOI21_X1  g592(.A(new_n1011), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1012), .A2(new_n1011), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1019), .B1(new_n1016), .B2(new_n1011), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1020), .B1(new_n988), .B2(G8), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1010), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT120), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(KEYINPUT120), .B(new_n1010), .C1(new_n1018), .C2(new_n1021), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n1024), .A2(KEYINPUT62), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT62), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1009), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OR2_X1    g603(.A1(new_n989), .A2(KEYINPUT63), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n831), .A2(KEYINPUT50), .A3(new_n910), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n943), .A2(new_n952), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n914), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  XOR2_X1   g607(.A(KEYINPUT56), .B(G2072), .Z(new_n1033));
  OAI22_X1  g608(.A1(new_n1032), .A2(G1956), .B1(new_n946), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT57), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n573), .A2(new_n1035), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n568), .A2(new_n572), .A3(KEYINPUT57), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1034), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OR2_X1    g613(.A1(new_n946), .A2(new_n1033), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1039), .B(new_n1040), .C1(G1956), .C2(new_n1032), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT116), .B1(new_n965), .B2(G2067), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n911), .A2(new_n914), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(new_n1045), .A3(new_n919), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n954), .A2(new_n802), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1043), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n607), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1038), .B1(new_n1042), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1041), .A2(new_n1038), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT61), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g628(.A(KEYINPUT58), .B(G1341), .ZN(new_n1054));
  OAI22_X1  g629(.A1(new_n946), .A2(G1996), .B1(new_n1044), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n555), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1056), .B(KEYINPUT59), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1041), .A2(new_n1038), .A3(KEYINPUT61), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1053), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1048), .A2(KEYINPUT60), .ZN(new_n1060));
  OAI211_X1 g635(.A(KEYINPUT117), .B(new_n1049), .C1(new_n1060), .C2(new_n607), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT117), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1049), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n607), .B1(new_n1048), .B2(KEYINPUT60), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1061), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT60), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1059), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1061), .A2(new_n1065), .A3(KEYINPUT60), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1050), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1002), .B1(KEYINPUT123), .B2(new_n792), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(KEYINPUT123), .B2(new_n792), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1073), .B1(new_n911), .B2(new_n912), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n914), .A2(KEYINPUT122), .ZN(new_n1075));
  OR2_X1    g650(.A1(new_n914), .A2(KEYINPUT122), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1074), .A2(new_n945), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1077), .A2(new_n1003), .A3(new_n1006), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1071), .B1(new_n1078), .B2(G171), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1079), .B1(G171), .B2(new_n1007), .ZN(new_n1080));
  XNOR2_X1  g655(.A(new_n1080), .B(KEYINPUT125), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1077), .A2(new_n1003), .A3(G301), .A4(new_n1006), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT124), .ZN(new_n1083));
  XNOR2_X1  g658(.A(new_n1082), .B(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1071), .B1(new_n1009), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1081), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1028), .B(new_n1029), .C1(new_n1070), .C2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n949), .ZN(new_n1089));
  AOI211_X1 g664(.A(G2090), .B(new_n914), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1090));
  OAI21_X1  g665(.A(G8), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AOI211_X1 g666(.A(new_n981), .B(new_n992), .C1(new_n963), .C2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1001), .B1(new_n1088), .B2(new_n1092), .ZN(new_n1093));
  XOR2_X1   g668(.A(G290), .B(G1986), .Z(new_n1094));
  NOR2_X1   g669(.A1(new_n1094), .A2(new_n922), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n1095), .B(KEYINPUT108), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n926), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n942), .B1(new_n1093), .B2(new_n1097), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g673(.A1(G229), .A2(new_n461), .A3(G227), .A4(G401), .ZN(new_n1100));
  NAND2_X1  g674(.A1(new_n847), .A2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g675(.A1(new_n908), .A2(new_n1101), .ZN(G308));
  OR2_X1    g676(.A1(new_n908), .A2(new_n1101), .ZN(G225));
endmodule


