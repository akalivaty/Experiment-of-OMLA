//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(G8gat), .ZN(new_n206));
  INV_X1    g005(.A(G50gat), .ZN(new_n207));
  AND2_X1   g006(.A1(new_n207), .A2(G43gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT15), .B1(new_n207), .B2(G43gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(KEYINPUT83), .B(G36gat), .Z(new_n211));
  INV_X1    g010(.A(G29gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(G29gat), .A2(G36gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(KEYINPUT14), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n210), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n216), .B(KEYINPUT84), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n213), .B1(KEYINPUT86), .B2(new_n215), .ZN(new_n218));
  INV_X1    g017(.A(new_n210), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT15), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT85), .B(G43gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(G50gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n207), .A2(G43gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n220), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n215), .A2(KEYINPUT86), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n218), .A2(new_n219), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n217), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT17), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT17), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n217), .A2(new_n229), .A3(new_n226), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n206), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n227), .A2(new_n206), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT18), .ZN(new_n234));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n235), .B(KEYINPUT87), .Z(new_n236));
  NOR4_X1   g035(.A1(new_n231), .A2(new_n233), .A3(new_n234), .A4(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n230), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n229), .B1(new_n217), .B2(new_n226), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n232), .B1(new_n241), .B2(new_n206), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n234), .B1(new_n242), .B2(new_n236), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT89), .B1(new_n227), .B2(new_n206), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(new_n232), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n236), .B(KEYINPUT88), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(KEYINPUT13), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n238), .A2(new_n243), .A3(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(G169gat), .B(G197gat), .Z(new_n250));
  XNOR2_X1  g049(.A(G113gat), .B(G141gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT80), .B(KEYINPUT11), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n256), .B(KEYINPUT12), .Z(new_n257));
  NAND2_X1  g056(.A1(new_n249), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n257), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n238), .A2(new_n259), .A3(new_n243), .A4(new_n248), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(G8gat), .B(G36gat), .Z(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(G64gat), .ZN(new_n264));
  INV_X1    g063(.A(G92gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G226gat), .A2(G233gat), .ZN(new_n267));
  OR2_X1    g066(.A1(G183gat), .A2(G190gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(G183gat), .A2(G190gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(KEYINPUT24), .A3(new_n269), .ZN(new_n270));
  OR2_X1    g069(.A1(new_n269), .A2(KEYINPUT24), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(KEYINPUT65), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT25), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT23), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n275), .B1(G169gat), .B2(G176gat), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n270), .A2(new_n271), .A3(new_n276), .ZN(new_n277));
  AND2_X1   g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278));
  NOR2_X1   g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n278), .B1(KEYINPUT23), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n274), .A2(new_n277), .A3(new_n280), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n280), .A2(new_n270), .A3(new_n271), .A4(new_n276), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n282), .A2(new_n273), .A3(new_n272), .ZN(new_n283));
  OR2_X1    g082(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n285));
  AOI21_X1  g084(.A(G190gat), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G190gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n290));
  AND2_X1   g089(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n289), .B(new_n290), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n269), .ZN(new_n295));
  NOR3_X1   g094(.A1(new_n288), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n279), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n297), .B(KEYINPUT67), .C1(KEYINPUT26), .C2(new_n278), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT67), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n299), .B1(new_n300), .B2(new_n279), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n298), .B(new_n301), .C1(KEYINPUT26), .C2(new_n297), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n281), .A2(new_n283), .B1(new_n296), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n267), .B1(new_n303), .B2(KEYINPUT29), .ZN(new_n304));
  XNOR2_X1  g103(.A(G197gat), .B(G204gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT22), .ZN(new_n306));
  INV_X1    g105(.A(G211gat), .ZN(new_n307));
  INV_X1    g106(.A(G218gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G211gat), .B(G218gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(new_n305), .A3(new_n309), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n294), .A2(new_n295), .ZN(new_n316));
  INV_X1    g115(.A(new_n288), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n302), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  AND3_X1   g117(.A1(new_n282), .A2(new_n273), .A3(new_n272), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n282), .B1(new_n273), .B2(new_n272), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  XOR2_X1   g120(.A(new_n267), .B(KEYINPUT71), .Z(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  AND3_X1   g123(.A1(new_n304), .A2(new_n315), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT70), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n315), .B(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n322), .B1(new_n303), .B2(KEYINPUT29), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n321), .A2(G226gat), .A3(G233gat), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n266), .B1(new_n325), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n327), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT29), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n323), .B1(new_n321), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n303), .A2(new_n267), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n332), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n304), .A2(new_n315), .A3(new_n324), .ZN(new_n337));
  INV_X1    g136(.A(new_n266), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n331), .A2(KEYINPUT30), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT30), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n336), .A2(new_n337), .A3(new_n341), .A4(new_n338), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G227gat), .A2(G233gat), .ZN(new_n344));
  XOR2_X1   g143(.A(new_n344), .B(KEYINPUT64), .Z(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(G120gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(G113gat), .ZN(new_n348));
  INV_X1    g147(.A(G113gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G120gat), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT1), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  XOR2_X1   g150(.A(G127gat), .B(G134gat), .Z(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G134gat), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n354), .A2(KEYINPUT68), .A3(G127gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(G127gat), .B(G134gat), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT68), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n353), .B1(new_n358), .B2(new_n351), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n359), .B(new_n318), .C1(new_n319), .C2(new_n320), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n281), .A2(new_n283), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n359), .B1(new_n362), .B2(new_n318), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n346), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT33), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G15gat), .B(G43gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(G71gat), .B(G99gat), .ZN(new_n368));
  XOR2_X1   g167(.A(new_n367), .B(new_n368), .Z(new_n369));
  NAND2_X1  g168(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n364), .A2(KEYINPUT32), .ZN(new_n371));
  INV_X1    g170(.A(new_n359), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n321), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT34), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n373), .A2(new_n374), .A3(new_n345), .A4(new_n360), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(new_n344), .A3(new_n360), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT34), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n371), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n371), .B1(new_n377), .B2(new_n375), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n370), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n377), .A2(new_n375), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n382), .A2(KEYINPUT32), .A3(new_n364), .ZN(new_n383));
  INV_X1    g182(.A(new_n370), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n384), .A3(new_n378), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT73), .ZN(new_n387));
  XNOR2_X1  g186(.A(G155gat), .B(G162gat), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT2), .ZN(new_n389));
  INV_X1    g188(.A(G148gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(G141gat), .ZN(new_n391));
  INV_X1    g190(.A(G141gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(G148gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n388), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT72), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n391), .A2(new_n393), .A3(KEYINPUT72), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(G155gat), .A2(G162gat), .ZN(new_n400));
  INV_X1    g199(.A(G155gat), .ZN(new_n401));
  INV_X1    g200(.A(G162gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n400), .B1(new_n403), .B2(KEYINPUT2), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n395), .B1(new_n399), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT3), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n387), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n391), .A2(new_n393), .A3(KEYINPUT72), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT72), .B1(new_n391), .B2(new_n393), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n404), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n389), .ZN(new_n411));
  INV_X1    g210(.A(new_n388), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n410), .A2(new_n387), .A3(new_n413), .A4(new_n406), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n333), .B1(new_n407), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n315), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n416), .A2(KEYINPUT75), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT75), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n410), .A2(new_n406), .A3(new_n413), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT73), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT29), .B1(new_n421), .B2(new_n414), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n419), .B1(new_n422), .B2(new_n315), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n315), .A2(new_n333), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n405), .B1(new_n424), .B2(new_n406), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n418), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(G228gat), .A2(G233gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n416), .A2(new_n332), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n425), .B1(new_n430), .B2(KEYINPUT76), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n422), .A2(new_n327), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT76), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n428), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n429), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT77), .B1(new_n436), .B2(G22gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(G78gat), .B(G106gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT31), .B(G50gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(G22gat), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n429), .A2(new_n435), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n442), .B1(new_n429), .B2(new_n435), .ZN(new_n445));
  OAI22_X1  g244(.A1(new_n437), .A2(new_n441), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n436), .A2(G22gat), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n447), .A2(KEYINPUT77), .A3(new_n443), .A4(new_n440), .ZN(new_n448));
  AOI211_X1 g247(.A(new_n343), .B(new_n386), .C1(new_n446), .C2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n410), .A2(new_n413), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT3), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n372), .B(new_n451), .C1(new_n407), .C2(new_n415), .ZN(new_n452));
  NAND2_X1  g251(.A1(G225gat), .A2(G233gat), .ZN(new_n453));
  AND4_X1   g252(.A1(KEYINPUT4), .A2(new_n359), .A3(new_n410), .A4(new_n413), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT4), .B1(new_n405), .B2(new_n359), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n452), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT5), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n405), .B(new_n359), .ZN(new_n459));
  INV_X1    g258(.A(new_n453), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(KEYINPUT0), .B(G57gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n463), .B(G85gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(G1gat), .B(G29gat), .ZN(new_n465));
  XOR2_X1   g264(.A(new_n464), .B(new_n465), .Z(new_n466));
  NAND4_X1  g265(.A1(new_n452), .A2(new_n456), .A3(new_n458), .A4(new_n453), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n462), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT6), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n462), .A2(new_n467), .ZN(new_n471));
  INV_X1    g270(.A(new_n466), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT78), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT78), .ZN(new_n474));
  AOI211_X1 g273(.A(new_n474), .B(new_n466), .C1(new_n462), .C2(new_n467), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n470), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT79), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n471), .A2(KEYINPUT6), .A3(new_n472), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT79), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n470), .B(new_n479), .C1(new_n473), .C2(new_n475), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n477), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT35), .B1(new_n449), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n386), .ZN(new_n483));
  INV_X1    g282(.A(new_n343), .ZN(new_n484));
  INV_X1    g283(.A(new_n448), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT77), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n428), .A2(new_n427), .B1(new_n431), .B2(new_n434), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n486), .B1(new_n487), .B2(new_n442), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n488), .A2(new_n440), .B1(new_n447), .B2(new_n443), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n483), .B(new_n484), .C1(new_n485), .C2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT35), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n468), .A2(KEYINPUT74), .A3(new_n469), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n471), .A2(new_n472), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT74), .B1(new_n468), .B2(new_n469), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n478), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n490), .A2(new_n491), .A3(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n482), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n496), .A2(new_n484), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(new_n448), .A3(new_n446), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT69), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT36), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(KEYINPUT69), .A2(KEYINPUT36), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n386), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n381), .A2(new_n385), .A3(new_n502), .A4(new_n503), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT37), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n336), .A2(new_n509), .A3(new_n337), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(new_n266), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n509), .B1(new_n336), .B2(new_n337), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT38), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n334), .A2(new_n335), .A3(new_n332), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n315), .B1(new_n304), .B2(new_n324), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT37), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT38), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n516), .A2(new_n517), .A3(new_n266), .A4(new_n510), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n513), .A2(new_n339), .A3(new_n518), .ZN(new_n519));
  AND4_X1   g318(.A1(new_n478), .A2(new_n477), .A3(new_n519), .A4(new_n480), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n493), .A2(new_n474), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n471), .A2(KEYINPUT78), .A3(new_n472), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n452), .A2(new_n456), .ZN(new_n524));
  OR3_X1    g323(.A1(new_n524), .A2(KEYINPUT39), .A3(new_n453), .ZN(new_n525));
  OR2_X1    g324(.A1(new_n459), .A2(new_n460), .ZN(new_n526));
  OAI211_X1 g325(.A(KEYINPUT39), .B(new_n526), .C1(new_n524), .C2(new_n453), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(new_n466), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT40), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n525), .A2(KEYINPUT40), .A3(new_n466), .A4(new_n527), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n343), .A2(new_n523), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n532), .B1(new_n485), .B2(new_n489), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n501), .B(new_n508), .C1(new_n520), .C2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n262), .B1(new_n499), .B2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT91), .B(G64gat), .ZN(new_n536));
  INV_X1    g335(.A(G57gat), .ZN(new_n537));
  OR3_X1    g336(.A1(new_n536), .A2(KEYINPUT92), .A3(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G71gat), .B(G78gat), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT9), .ZN(new_n540));
  INV_X1    g339(.A(G71gat), .ZN(new_n541));
  INV_X1    g340(.A(G78gat), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n538), .A2(new_n539), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n537), .A2(G64gat), .ZN(new_n545));
  OAI211_X1 g344(.A(KEYINPUT92), .B(new_n545), .C1(new_n536), .C2(new_n537), .ZN(new_n546));
  INV_X1    g345(.A(new_n539), .ZN(new_n547));
  XNOR2_X1  g346(.A(G57gat), .B(G64gat), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n548), .A2(KEYINPUT90), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(KEYINPUT90), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n549), .A2(new_n543), .A3(new_n550), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n544), .A2(new_n546), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n206), .B1(new_n552), .B2(KEYINPUT21), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT93), .ZN(new_n554));
  XOR2_X1   g353(.A(G127gat), .B(G155gat), .Z(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(G183gat), .B(G211gat), .Z(new_n557));
  NAND2_X1  g356(.A1(G231gat), .A2(G233gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n556), .B(new_n559), .Z(new_n560));
  NOR2_X1   g359(.A1(new_n552), .A2(KEYINPUT21), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n560), .A2(new_n563), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(G190gat), .B(G218gat), .Z(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT98), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(KEYINPUT94), .A2(G85gat), .A3(G92gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT7), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT96), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(G85gat), .ZN(new_n576));
  NOR3_X1   g375(.A1(new_n576), .A2(new_n265), .A3(KEYINPUT95), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n577), .A2(KEYINPUT94), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n573), .B(KEYINPUT96), .ZN(new_n580));
  INV_X1    g379(.A(new_n578), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(G99gat), .A2(G106gat), .ZN(new_n583));
  AOI22_X1  g382(.A1(KEYINPUT8), .A2(new_n583), .B1(new_n576), .B2(new_n265), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n579), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT97), .ZN(new_n586));
  XOR2_X1   g385(.A(G99gat), .B(G106gat), .Z(new_n587));
  NAND3_X1  g386(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n585), .A2(new_n587), .ZN(new_n589));
  INV_X1    g388(.A(new_n587), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n579), .A2(new_n582), .A3(new_n590), .A4(new_n584), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n589), .A2(KEYINPUT97), .A3(new_n591), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n588), .B(new_n592), .C1(new_n239), .C2(new_n240), .ZN(new_n593));
  AND3_X1   g392(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n588), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n594), .B1(new_n595), .B2(new_n227), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n571), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  AOI211_X1 g399(.A(new_n571), .B(new_n598), .C1(new_n593), .C2(new_n596), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n569), .A2(new_n570), .ZN(new_n603));
  XOR2_X1   g402(.A(G134gat), .B(G162gat), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n605), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n607), .B1(new_n600), .B2(new_n601), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n589), .A2(new_n552), .A3(new_n591), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n611), .B1(new_n595), .B2(new_n552), .ZN(new_n612));
  NAND2_X1  g411(.A1(G230gat), .A2(G233gat), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n616), .A2(KEYINPUT99), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT10), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n611), .B(new_n618), .C1(new_n595), .C2(new_n552), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n595), .A2(KEYINPUT10), .A3(new_n552), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n614), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G120gat), .B(G148gat), .ZN(new_n623));
  INV_X1    g422(.A(G176gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n625), .B(G204gat), .Z(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n616), .A2(KEYINPUT99), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n617), .A2(new_n622), .A3(new_n627), .A4(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n627), .B1(new_n622), .B2(new_n615), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n567), .A2(new_n610), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n535), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n497), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(G1gat), .ZN(G1324gat));
  OAI21_X1  g437(.A(G8gat), .B1(new_n635), .B2(new_n484), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(KEYINPUT42), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT100), .B(G8gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n635), .A2(new_n484), .A3(new_n642), .ZN(new_n643));
  MUX2_X1   g442(.A(new_n640), .B(KEYINPUT42), .S(new_n643), .Z(G1325gat));
  INV_X1    g443(.A(G15gat), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n635), .A2(new_n645), .A3(new_n508), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n636), .A2(new_n483), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n646), .B1(new_n645), .B2(new_n647), .ZN(G1326gat));
  NAND2_X1  g447(.A1(new_n446), .A2(new_n448), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n635), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT43), .B(G22gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT101), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n650), .B(new_n652), .ZN(G1327gat));
  INV_X1    g452(.A(KEYINPUT103), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n534), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n477), .A2(new_n519), .A3(new_n478), .A4(new_n480), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n656), .A2(new_n649), .A3(new_n532), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n657), .A2(KEYINPUT103), .A3(new_n501), .A4(new_n508), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n499), .A2(new_n655), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n610), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT44), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n661), .B1(new_n499), .B2(new_n534), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n566), .B1(new_n664), .B2(new_n610), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT102), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n231), .A2(new_n233), .ZN(new_n668));
  INV_X1    g467(.A(new_n236), .ZN(new_n669));
  AOI21_X1  g468(.A(KEYINPUT18), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(new_n237), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n259), .B1(new_n671), .B2(new_n248), .ZN(new_n672));
  INV_X1    g471(.A(new_n260), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n667), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n258), .A2(KEYINPUT102), .A3(new_n260), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NOR4_X1   g476(.A1(new_n663), .A2(new_n666), .A3(new_n633), .A4(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(G29gat), .B1(new_n679), .B2(new_n496), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n535), .A2(new_n610), .A3(new_n632), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n681), .A2(new_n566), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n682), .A2(new_n212), .A3(new_n497), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT45), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n680), .A2(new_n684), .ZN(G1328gat));
  NAND3_X1  g484(.A1(new_n682), .A2(new_n343), .A3(new_n211), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(KEYINPUT46), .Z(new_n687));
  NOR2_X1   g486(.A1(new_n679), .A2(new_n484), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n687), .B1(new_n688), .B2(new_n211), .ZN(G1329gat));
  INV_X1    g488(.A(new_n508), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n221), .B1(new_n678), .B2(new_n690), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n682), .A2(new_n483), .A3(new_n221), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g493(.A(new_n649), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n678), .A2(G50gat), .A3(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n682), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n207), .B1(new_n697), .B2(new_n649), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g499(.A1(new_n567), .A2(new_n610), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n676), .A2(new_n632), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n659), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(KEYINPUT104), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT104), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n659), .A2(new_n705), .A3(new_n701), .A4(new_n702), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n496), .B(KEYINPUT105), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n704), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g508(.A1(new_n704), .A2(new_n706), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n710), .A2(new_n484), .ZN(new_n711));
  NOR2_X1   g510(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(KEYINPUT49), .B(G64gat), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n713), .B1(new_n711), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT106), .B(KEYINPUT107), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1333gat));
  OAI21_X1  g516(.A(new_n541), .B1(new_n710), .B2(new_n386), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n704), .A2(G71gat), .A3(new_n690), .A4(new_n706), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n719), .A2(KEYINPUT108), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n719), .A2(KEYINPUT108), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n718), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(KEYINPUT109), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n724), .B(new_n718), .C1(new_n720), .C2(new_n721), .ZN(new_n725));
  AND3_X1   g524(.A1(new_n723), .A2(KEYINPUT50), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT50), .B1(new_n723), .B2(new_n725), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(G1334gat));
  NOR2_X1   g527(.A1(new_n710), .A2(new_n649), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(new_n542), .ZN(G1335gat));
  NOR2_X1   g529(.A1(new_n663), .A2(new_n666), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n731), .A2(new_n702), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G85gat), .B1(new_n733), .B2(new_n496), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n659), .A2(new_n567), .A3(new_n610), .A4(new_n677), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT51), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT51), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n737), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT111), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n736), .A2(KEYINPUT110), .A3(KEYINPUT51), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n742), .B1(new_n741), .B2(new_n743), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n576), .B(new_n497), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n734), .B1(new_n747), .B2(new_n632), .ZN(G1336gat));
  NAND3_X1  g547(.A1(new_n732), .A2(KEYINPUT112), .A3(new_n343), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n731), .A2(new_n343), .A3(new_n702), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT112), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n749), .A2(G92gat), .A3(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n741), .A2(new_n743), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n633), .A2(new_n265), .A3(new_n343), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n753), .B(new_n754), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n750), .A2(G92gat), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n756), .B1(new_n737), .B2(new_n740), .ZN(new_n759));
  OAI21_X1  g558(.A(KEYINPUT52), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n760), .ZN(G1337gat));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n632), .A2(G99gat), .A3(new_n386), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n755), .A2(KEYINPUT111), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n764), .B1(new_n765), .B2(new_n744), .ZN(new_n766));
  INV_X1    g565(.A(G99gat), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n767), .B1(new_n732), .B2(new_n690), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n762), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n763), .B1(new_n745), .B2(new_n746), .ZN(new_n770));
  INV_X1    g569(.A(new_n768), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n770), .A2(new_n771), .A3(KEYINPUT113), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n769), .A2(new_n772), .ZN(G1338gat));
  NAND3_X1  g572(.A1(new_n731), .A2(new_n695), .A3(new_n702), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT53), .B1(new_n774), .B2(G106gat), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n632), .A2(G106gat), .A3(new_n649), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n775), .B1(new_n755), .B2(new_n777), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n774), .A2(KEYINPUT114), .A3(G106gat), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT114), .B1(new_n774), .B2(G106gat), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n777), .B1(new_n737), .B2(new_n740), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n778), .B1(new_n782), .B2(new_n783), .ZN(G1339gat));
  NAND2_X1  g583(.A1(new_n649), .A2(new_n483), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n245), .A2(new_n247), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n668), .A2(new_n669), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n256), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n260), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n609), .A2(new_n789), .ZN(new_n790));
  AOI211_X1 g589(.A(KEYINPUT54), .B(new_n614), .C1(new_n619), .C2(new_n620), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT115), .B1(new_n791), .B2(new_n627), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n621), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT115), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n794), .A2(new_n795), .A3(new_n626), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n619), .A2(new_n614), .A3(new_n620), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n622), .A2(KEYINPUT54), .A3(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n798), .B1(new_n797), .B2(new_n800), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n790), .B(new_n629), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n797), .A2(new_n800), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT55), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n630), .B1(new_n808), .B2(new_n801), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n809), .A2(KEYINPUT116), .A3(new_n790), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n808), .A2(new_n801), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n812), .A2(new_n676), .A3(new_n629), .ZN(new_n813));
  INV_X1    g612(.A(new_n789), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n633), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n610), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n567), .B1(new_n811), .B2(new_n816), .ZN(new_n817));
  NOR4_X1   g616(.A1(new_n567), .A2(new_n610), .A3(new_n633), .A4(new_n676), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n785), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n820), .A2(new_n497), .A3(new_n484), .ZN(new_n821));
  OAI21_X1  g620(.A(G113gat), .B1(new_n821), .B2(new_n262), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n707), .A2(new_n484), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(new_n817), .B2(new_n819), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n824), .A2(new_n649), .A3(new_n483), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n676), .A2(new_n349), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n822), .B1(new_n825), .B2(new_n826), .ZN(G1340gat));
  OR3_X1    g626(.A1(new_n825), .A2(G120gat), .A3(new_n632), .ZN(new_n828));
  OAI21_X1  g627(.A(G120gat), .B1(new_n821), .B2(new_n632), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(G1341gat));
  NOR2_X1   g629(.A1(new_n825), .A2(new_n567), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n566), .A2(G127gat), .ZN(new_n832));
  OAI22_X1  g631(.A1(new_n831), .A2(G127gat), .B1(new_n821), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT117), .ZN(G1342gat));
  NOR3_X1   g633(.A1(new_n825), .A2(G134gat), .A3(new_n609), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT56), .ZN(new_n836));
  OAI21_X1  g635(.A(G134gat), .B1(new_n821), .B2(new_n609), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(G1343gat));
  AOI22_X1  g637(.A1(new_n809), .A2(new_n261), .B1(new_n633), .B2(new_n814), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n806), .B(new_n810), .C1(new_n839), .C2(new_n610), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n818), .B1(new_n840), .B2(new_n567), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT57), .B1(new_n841), .B2(new_n649), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n817), .A2(new_n819), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n843), .A2(new_n844), .A3(new_n695), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n690), .A2(new_n496), .A3(new_n343), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n842), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(G141gat), .B1(new_n847), .B2(new_n262), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT58), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n690), .A2(new_n649), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n824), .A2(new_n392), .A3(new_n261), .A4(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n851), .A2(new_n852), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n848), .A2(new_n849), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n851), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n850), .ZN(new_n859));
  AOI211_X1 g658(.A(new_n823), .B(new_n859), .C1(new_n817), .C2(new_n819), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n860), .A2(KEYINPUT118), .A3(new_n392), .A4(new_n261), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n842), .A2(new_n845), .A3(new_n676), .A4(new_n846), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(G141gat), .ZN(new_n864));
  AOI211_X1 g663(.A(new_n856), .B(new_n849), .C1(new_n862), .C2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n864), .A2(new_n858), .A3(new_n861), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT119), .B1(new_n866), .B2(KEYINPUT58), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n855), .B1(new_n865), .B2(new_n867), .ZN(G1344gat));
  NAND3_X1  g667(.A1(new_n860), .A2(new_n390), .A3(new_n633), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n843), .A2(new_n695), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT57), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n804), .B1(new_n839), .B2(new_n610), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n873), .A2(new_n567), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n634), .A2(new_n262), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n844), .B(new_n695), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n633), .A3(new_n846), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n870), .B1(new_n878), .B2(G148gat), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n870), .B1(new_n847), .B2(new_n632), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(new_n390), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n869), .B1(new_n879), .B2(new_n881), .ZN(G1345gat));
  AOI21_X1  g681(.A(G155gat), .B1(new_n860), .B2(new_n566), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n847), .A2(new_n401), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n883), .B1(new_n884), .B2(new_n566), .ZN(G1346gat));
  AOI21_X1  g684(.A(G162gat), .B1(new_n860), .B2(new_n610), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n847), .A2(new_n402), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(new_n610), .ZN(G1347gat));
  NAND3_X1  g687(.A1(new_n820), .A2(new_n496), .A3(new_n343), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n889), .A2(KEYINPUT121), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(KEYINPUT121), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n677), .A2(G169gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n707), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n820), .A2(new_n343), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(G169gat), .B1(new_n895), .B2(new_n262), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT122), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n896), .A2(new_n897), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n893), .B1(new_n898), .B2(new_n899), .ZN(G1348gat));
  NOR3_X1   g699(.A1(new_n895), .A2(new_n624), .A3(new_n632), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n890), .A2(new_n633), .A3(new_n891), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n902), .B2(new_n624), .ZN(G1349gat));
  OR3_X1    g702(.A1(new_n895), .A2(KEYINPUT123), .A3(new_n567), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT123), .B1(new_n895), .B2(new_n567), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(G183gat), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n889), .B1(new_n284), .B2(new_n285), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n566), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT60), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT60), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n906), .A2(new_n911), .A3(new_n908), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(G1350gat));
  OAI21_X1  g712(.A(G190gat), .B1(new_n895), .B2(new_n609), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n914), .A2(KEYINPUT125), .A3(new_n915), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n914), .A2(KEYINPUT125), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n914), .A2(KEYINPUT125), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n917), .A2(KEYINPUT61), .A3(new_n918), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n890), .A2(new_n289), .A3(new_n610), .A4(new_n891), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT124), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n920), .A2(new_n921), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n916), .B(new_n919), .C1(new_n922), .C2(new_n923), .ZN(G1351gat));
  NOR3_X1   g723(.A1(new_n690), .A2(new_n484), .A3(new_n707), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n877), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(G197gat), .B1(new_n926), .B2(new_n262), .ZN(new_n927));
  AOI211_X1 g726(.A(new_n497), .B(new_n484), .C1(new_n817), .C2(new_n819), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n850), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n929), .A2(G197gat), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n927), .B1(new_n677), .B2(new_n930), .ZN(G1352gat));
  XNOR2_X1  g730(.A(KEYINPUT126), .B(G204gat), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n929), .A2(new_n632), .A3(new_n932), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT62), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n872), .A2(new_n633), .A3(new_n876), .A4(new_n925), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT127), .ZN(new_n936));
  OR2_X1    g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(new_n936), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n937), .A2(new_n932), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n934), .A2(new_n939), .ZN(G1353gat));
  INV_X1    g739(.A(new_n929), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n941), .A2(new_n307), .A3(new_n566), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n877), .A2(new_n566), .A3(new_n925), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n943), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n944));
  AOI21_X1  g743(.A(KEYINPUT63), .B1(new_n943), .B2(G211gat), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(G1354gat));
  OAI21_X1  g745(.A(G218gat), .B1(new_n926), .B2(new_n609), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n941), .A2(new_n308), .A3(new_n610), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(G1355gat));
endmodule


