

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U550 ( .A1(G651), .A2(n553), .ZN(n794) );
  NAND2_X2 U551 ( .A1(n611), .A2(n610), .ZN(n940) );
  NOR2_X2 U552 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X2 U553 ( .A1(n614), .A2(G8), .ZN(n707) );
  NOR2_X1 U554 ( .A1(n733), .A2(n732), .ZN(n744) );
  INV_X1 U555 ( .A(n612), .ZN(n614) );
  NAND2_X1 U556 ( .A1(G160), .A2(G40), .ZN(n710) );
  NOR2_X2 U557 ( .A1(n549), .A2(n548), .ZN(G160) );
  XNOR2_X1 U558 ( .A(n619), .B(n618), .ZN(n633) );
  INV_X1 U559 ( .A(KEYINPUT64), .ZN(n618) );
  NOR2_X1 U560 ( .A1(n940), .A2(n617), .ZN(n619) );
  AND2_X1 U561 ( .A1(n587), .A2(n586), .ZN(n711) );
  NOR2_X1 U562 ( .A1(n707), .A2(n689), .ZN(n513) );
  OR2_X1 U563 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U564 ( .A1(n682), .A2(n675), .ZN(n654) );
  XNOR2_X1 U565 ( .A(n600), .B(KEYINPUT95), .ZN(n629) );
  NOR2_X1 U566 ( .A1(n629), .A2(n926), .ZN(n630) );
  BUF_X1 U567 ( .A(n612), .Z(n646) );
  BUF_X1 U568 ( .A(n614), .Z(n652) );
  NOR2_X1 U569 ( .A1(G2084), .A2(n652), .ZN(n675) );
  OR2_X1 U570 ( .A1(n707), .A2(G1966), .ZN(n651) );
  XNOR2_X1 U571 ( .A(n651), .B(KEYINPUT93), .ZN(n682) );
  INV_X1 U572 ( .A(n928), .ZN(n689) );
  AND2_X1 U573 ( .A1(n690), .A2(n513), .ZN(n691) );
  NOR2_X2 U574 ( .A1(n588), .A2(n710), .ZN(n612) );
  INV_X1 U575 ( .A(G1384), .ZN(n586) );
  INV_X1 U576 ( .A(G2104), .ZN(n528) );
  AND2_X1 U577 ( .A1(n534), .A2(G2104), .ZN(n539) );
  INV_X1 U578 ( .A(KEYINPUT23), .ZN(n540) );
  XNOR2_X1 U579 ( .A(KEYINPUT107), .B(KEYINPUT40), .ZN(n763) );
  OR2_X1 U580 ( .A1(n538), .A2(n537), .ZN(n587) );
  XNOR2_X1 U581 ( .A(KEYINPUT7), .B(n527), .ZN(G168) );
  NOR2_X1 U582 ( .A1(G651), .A2(G543), .ZN(n798) );
  NAND2_X1 U583 ( .A1(n798), .A2(G89), .ZN(n514) );
  XNOR2_X1 U584 ( .A(n514), .B(KEYINPUT4), .ZN(n516) );
  XOR2_X1 U585 ( .A(KEYINPUT0), .B(G543), .Z(n553) );
  INV_X1 U586 ( .A(G651), .ZN(n520) );
  NOR2_X1 U587 ( .A1(n553), .A2(n520), .ZN(n797) );
  NAND2_X1 U588 ( .A1(G76), .A2(n797), .ZN(n515) );
  NAND2_X1 U589 ( .A1(n516), .A2(n515), .ZN(n519) );
  XOR2_X1 U590 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n517) );
  XNOR2_X1 U591 ( .A(KEYINPUT5), .B(n517), .ZN(n518) );
  XNOR2_X1 U592 ( .A(n519), .B(n518), .ZN(n526) );
  NOR2_X1 U593 ( .A1(G543), .A2(n520), .ZN(n521) );
  XOR2_X1 U594 ( .A(KEYINPUT1), .B(n521), .Z(n793) );
  NAND2_X1 U595 ( .A1(G63), .A2(n793), .ZN(n523) );
  NAND2_X1 U596 ( .A1(G51), .A2(n794), .ZN(n522) );
  NAND2_X1 U597 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U598 ( .A(KEYINPUT6), .B(n524), .Z(n525) );
  NAND2_X1 U599 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X2 U600 ( .A1(n528), .A2(G2105), .ZN(n903) );
  NAND2_X1 U601 ( .A1(G126), .A2(n903), .ZN(n532) );
  NAND2_X1 U602 ( .A1(G2105), .A2(G2104), .ZN(n530) );
  INV_X1 U603 ( .A(KEYINPUT66), .ZN(n529) );
  XNOR2_X2 U604 ( .A(n530), .B(n529), .ZN(n901) );
  NAND2_X1 U605 ( .A1(n901), .A2(G114), .ZN(n531) );
  NAND2_X1 U606 ( .A1(n532), .A2(n531), .ZN(n538) );
  NOR2_X1 U607 ( .A1(G2105), .A2(G2104), .ZN(n533) );
  XOR2_X1 U608 ( .A(KEYINPUT17), .B(n533), .Z(n716) );
  NAND2_X1 U609 ( .A1(G138), .A2(n716), .ZN(n536) );
  INV_X1 U610 ( .A(G2105), .ZN(n534) );
  BUF_X1 U611 ( .A(n539), .Z(n908) );
  NAND2_X1 U612 ( .A1(G102), .A2(n908), .ZN(n535) );
  NAND2_X1 U613 ( .A1(n536), .A2(n535), .ZN(n537) );
  INV_X1 U614 ( .A(n587), .ZN(G164) );
  NAND2_X1 U615 ( .A1(n903), .A2(G125), .ZN(n543) );
  NAND2_X1 U616 ( .A1(n539), .A2(G101), .ZN(n541) );
  XNOR2_X1 U617 ( .A(n541), .B(n540), .ZN(n542) );
  NAND2_X1 U618 ( .A1(n543), .A2(n542), .ZN(n545) );
  INV_X1 U619 ( .A(KEYINPUT65), .ZN(n544) );
  XNOR2_X1 U620 ( .A(n545), .B(n544), .ZN(n549) );
  NAND2_X1 U621 ( .A1(n716), .A2(G137), .ZN(n547) );
  NAND2_X1 U622 ( .A1(G113), .A2(n901), .ZN(n546) );
  NAND2_X1 U623 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U624 ( .A1(G49), .A2(n794), .ZN(n551) );
  NAND2_X1 U625 ( .A1(G74), .A2(G651), .ZN(n550) );
  NAND2_X1 U626 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U627 ( .A1(n793), .A2(n552), .ZN(n555) );
  NAND2_X1 U628 ( .A1(n553), .A2(G87), .ZN(n554) );
  NAND2_X1 U629 ( .A1(n555), .A2(n554), .ZN(G288) );
  NAND2_X1 U630 ( .A1(G64), .A2(n793), .ZN(n557) );
  NAND2_X1 U631 ( .A1(G52), .A2(n794), .ZN(n556) );
  NAND2_X1 U632 ( .A1(n557), .A2(n556), .ZN(n562) );
  NAND2_X1 U633 ( .A1(G77), .A2(n797), .ZN(n559) );
  NAND2_X1 U634 ( .A1(G90), .A2(n798), .ZN(n558) );
  NAND2_X1 U635 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U636 ( .A(KEYINPUT9), .B(n560), .Z(n561) );
  NOR2_X1 U637 ( .A1(n562), .A2(n561), .ZN(G171) );
  NAND2_X1 U638 ( .A1(G75), .A2(n797), .ZN(n564) );
  NAND2_X1 U639 ( .A1(G88), .A2(n798), .ZN(n563) );
  NAND2_X1 U640 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U641 ( .A1(G62), .A2(n793), .ZN(n566) );
  NAND2_X1 U642 ( .A1(G50), .A2(n794), .ZN(n565) );
  NAND2_X1 U643 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U644 ( .A1(n568), .A2(n567), .ZN(G166) );
  INV_X1 U645 ( .A(G166), .ZN(G303) );
  XOR2_X1 U646 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U647 ( .A1(G86), .A2(n798), .ZN(n570) );
  NAND2_X1 U648 ( .A1(G61), .A2(n793), .ZN(n569) );
  NAND2_X1 U649 ( .A1(n570), .A2(n569), .ZN(n573) );
  NAND2_X1 U650 ( .A1(n797), .A2(G73), .ZN(n571) );
  XOR2_X1 U651 ( .A(KEYINPUT2), .B(n571), .Z(n572) );
  NOR2_X1 U652 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U653 ( .A1(n794), .A2(G48), .ZN(n574) );
  NAND2_X1 U654 ( .A1(n575), .A2(n574), .ZN(G305) );
  NAND2_X1 U655 ( .A1(n794), .A2(G47), .ZN(n584) );
  NAND2_X1 U656 ( .A1(n797), .A2(G72), .ZN(n576) );
  XOR2_X1 U657 ( .A(KEYINPUT67), .B(n576), .Z(n578) );
  NAND2_X1 U658 ( .A1(n798), .A2(G85), .ZN(n577) );
  NAND2_X1 U659 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U660 ( .A(KEYINPUT68), .B(n579), .ZN(n582) );
  NAND2_X1 U661 ( .A1(G60), .A2(n793), .ZN(n580) );
  XNOR2_X1 U662 ( .A(KEYINPUT69), .B(n580), .ZN(n581) );
  NOR2_X1 U663 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U664 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U665 ( .A(n585), .B(KEYINPUT70), .ZN(G290) );
  INV_X1 U666 ( .A(n711), .ZN(n588) );
  NOR2_X1 U667 ( .A1(G1976), .A2(G288), .ZN(n687) );
  NAND2_X1 U668 ( .A1(n687), .A2(KEYINPUT33), .ZN(n589) );
  NOR2_X1 U669 ( .A1(n707), .A2(n589), .ZN(n693) );
  NAND2_X1 U670 ( .A1(G65), .A2(n793), .ZN(n591) );
  NAND2_X1 U671 ( .A1(G53), .A2(n794), .ZN(n590) );
  NAND2_X1 U672 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U673 ( .A1(G78), .A2(n797), .ZN(n593) );
  NAND2_X1 U674 ( .A1(G91), .A2(n798), .ZN(n592) );
  NAND2_X1 U675 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U676 ( .A1(n595), .A2(n594), .ZN(n926) );
  NAND2_X1 U677 ( .A1(G1956), .A2(n652), .ZN(n596) );
  XNOR2_X1 U678 ( .A(n596), .B(KEYINPUT94), .ZN(n599) );
  NAND2_X1 U679 ( .A1(n646), .A2(G2072), .ZN(n597) );
  XOR2_X1 U680 ( .A(KEYINPUT27), .B(n597), .Z(n598) );
  NAND2_X1 U681 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U682 ( .A1(n926), .A2(n629), .ZN(n638) );
  INV_X1 U683 ( .A(n638), .ZN(n628) );
  NAND2_X1 U684 ( .A1(G81), .A2(n798), .ZN(n601) );
  XOR2_X1 U685 ( .A(KEYINPUT73), .B(n601), .Z(n602) );
  XNOR2_X1 U686 ( .A(n602), .B(KEYINPUT12), .ZN(n604) );
  NAND2_X1 U687 ( .A1(G68), .A2(n797), .ZN(n603) );
  NAND2_X1 U688 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U689 ( .A(KEYINPUT13), .B(n605), .ZN(n611) );
  NAND2_X1 U690 ( .A1(G56), .A2(n793), .ZN(n606) );
  XOR2_X1 U691 ( .A(KEYINPUT14), .B(n606), .Z(n609) );
  NAND2_X1 U692 ( .A1(n794), .A2(G43), .ZN(n607) );
  XOR2_X1 U693 ( .A(KEYINPUT74), .B(n607), .Z(n608) );
  AND2_X1 U694 ( .A1(n612), .A2(G1996), .ZN(n613) );
  XNOR2_X1 U695 ( .A(n613), .B(KEYINPUT26), .ZN(n616) );
  AND2_X1 U696 ( .A1(n614), .A2(G1341), .ZN(n615) );
  NAND2_X1 U697 ( .A1(G66), .A2(n793), .ZN(n621) );
  NAND2_X1 U698 ( .A1(G54), .A2(n794), .ZN(n620) );
  NAND2_X1 U699 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U700 ( .A1(G79), .A2(n797), .ZN(n623) );
  NAND2_X1 U701 ( .A1(G92), .A2(n798), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U703 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U704 ( .A(n626), .B(KEYINPUT15), .ZN(n941) );
  NAND2_X1 U705 ( .A1(n633), .A2(n941), .ZN(n627) );
  OR2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n632) );
  XOR2_X1 U707 ( .A(n630), .B(KEYINPUT28), .Z(n631) );
  AND2_X1 U708 ( .A1(n632), .A2(n631), .ZN(n643) );
  NOR2_X1 U709 ( .A1(n633), .A2(n941), .ZN(n634) );
  XOR2_X1 U710 ( .A(n634), .B(KEYINPUT96), .Z(n641) );
  AND2_X1 U711 ( .A1(n646), .A2(G2067), .ZN(n635) );
  XNOR2_X1 U712 ( .A(n635), .B(KEYINPUT97), .ZN(n637) );
  NAND2_X1 U713 ( .A1(n652), .A2(G1348), .ZN(n636) );
  NAND2_X1 U714 ( .A1(n637), .A2(n636), .ZN(n639) );
  AND2_X1 U715 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U716 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U717 ( .A1(n643), .A2(n642), .ZN(n645) );
  XOR2_X1 U718 ( .A(KEYINPUT98), .B(KEYINPUT29), .Z(n644) );
  XNOR2_X1 U719 ( .A(n645), .B(n644), .ZN(n650) );
  XNOR2_X1 U720 ( .A(G2078), .B(KEYINPUT25), .ZN(n981) );
  NOR2_X1 U721 ( .A1(n652), .A2(n981), .ZN(n648) );
  INV_X1 U722 ( .A(G1961), .ZN(n952) );
  NOR2_X1 U723 ( .A1(n646), .A2(n952), .ZN(n647) );
  NOR2_X1 U724 ( .A1(n648), .A2(n647), .ZN(n658) );
  NAND2_X1 U725 ( .A1(G171), .A2(n658), .ZN(n649) );
  NAND2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n678) );
  INV_X1 U727 ( .A(KEYINPUT99), .ZN(n653) );
  XNOR2_X1 U728 ( .A(n654), .B(n653), .ZN(n655) );
  NAND2_X1 U729 ( .A1(n655), .A2(G8), .ZN(n656) );
  XNOR2_X1 U730 ( .A(n656), .B(KEYINPUT30), .ZN(n657) );
  NOR2_X1 U731 ( .A1(n657), .A2(G168), .ZN(n660) );
  NOR2_X1 U732 ( .A1(G171), .A2(n658), .ZN(n659) );
  NOR2_X1 U733 ( .A1(n660), .A2(n659), .ZN(n662) );
  INV_X1 U734 ( .A(KEYINPUT31), .ZN(n661) );
  XNOR2_X1 U735 ( .A(n662), .B(n661), .ZN(n677) );
  INV_X1 U736 ( .A(G8), .ZN(n667) );
  NOR2_X1 U737 ( .A1(G1971), .A2(n707), .ZN(n664) );
  NOR2_X1 U738 ( .A1(G2090), .A2(n652), .ZN(n663) );
  NOR2_X1 U739 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U740 ( .A1(n665), .A2(G303), .ZN(n666) );
  OR2_X1 U741 ( .A1(n667), .A2(n666), .ZN(n669) );
  AND2_X1 U742 ( .A1(n677), .A2(n669), .ZN(n668) );
  NAND2_X1 U743 ( .A1(n678), .A2(n668), .ZN(n673) );
  INV_X1 U744 ( .A(n669), .ZN(n671) );
  AND2_X1 U745 ( .A1(G286), .A2(G8), .ZN(n670) );
  OR2_X1 U746 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U747 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U748 ( .A(n674), .B(KEYINPUT32), .ZN(n685) );
  NAND2_X1 U749 ( .A1(G8), .A2(n675), .ZN(n676) );
  XNOR2_X1 U750 ( .A(n676), .B(KEYINPUT92), .ZN(n680) );
  NAND2_X1 U751 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U752 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U753 ( .A1(n682), .A2(n681), .ZN(n683) );
  INV_X1 U754 ( .A(n683), .ZN(n684) );
  NAND2_X1 U755 ( .A1(n685), .A2(n684), .ZN(n695) );
  NOR2_X1 U756 ( .A1(G1971), .A2(G303), .ZN(n686) );
  NOR2_X1 U757 ( .A1(n687), .A2(n686), .ZN(n932) );
  XNOR2_X1 U758 ( .A(KEYINPUT100), .B(n932), .ZN(n688) );
  NAND2_X1 U759 ( .A1(n695), .A2(n688), .ZN(n690) );
  NAND2_X1 U760 ( .A1(G1976), .A2(G288), .ZN(n928) );
  NOR2_X1 U761 ( .A1(KEYINPUT33), .A2(n691), .ZN(n692) );
  NOR2_X1 U762 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U763 ( .A(G1981), .B(G305), .Z(n936) );
  NAND2_X1 U764 ( .A1(n694), .A2(n936), .ZN(n703) );
  INV_X1 U765 ( .A(n707), .ZN(n700) );
  INV_X1 U766 ( .A(n695), .ZN(n698) );
  NAND2_X1 U767 ( .A1(G166), .A2(G8), .ZN(n696) );
  NOR2_X1 U768 ( .A1(G2090), .A2(n696), .ZN(n697) );
  NOR2_X1 U769 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U770 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U771 ( .A(n701), .B(KEYINPUT101), .ZN(n702) );
  NAND2_X1 U772 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U773 ( .A(n704), .B(KEYINPUT102), .ZN(n709) );
  NOR2_X1 U774 ( .A1(G1981), .A2(G305), .ZN(n705) );
  XOR2_X1 U775 ( .A(n705), .B(KEYINPUT24), .Z(n706) );
  NOR2_X1 U776 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U777 ( .A1(n709), .A2(n708), .ZN(n733) );
  NOR2_X1 U778 ( .A1(n711), .A2(n710), .ZN(n759) );
  NAND2_X1 U779 ( .A1(G107), .A2(n901), .ZN(n712) );
  XOR2_X1 U780 ( .A(KEYINPUT89), .B(n712), .Z(n714) );
  NAND2_X1 U781 ( .A1(n903), .A2(G119), .ZN(n713) );
  NAND2_X1 U782 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U783 ( .A(KEYINPUT90), .B(n715), .ZN(n719) );
  BUF_X1 U784 ( .A(n716), .Z(n907) );
  NAND2_X1 U785 ( .A1(G131), .A2(n907), .ZN(n717) );
  XNOR2_X1 U786 ( .A(KEYINPUT91), .B(n717), .ZN(n718) );
  NOR2_X1 U787 ( .A1(n719), .A2(n718), .ZN(n721) );
  NAND2_X1 U788 ( .A1(n908), .A2(G95), .ZN(n720) );
  NAND2_X1 U789 ( .A1(n721), .A2(n720), .ZN(n898) );
  NAND2_X1 U790 ( .A1(G1991), .A2(n898), .ZN(n730) );
  NAND2_X1 U791 ( .A1(G129), .A2(n903), .ZN(n723) );
  NAND2_X1 U792 ( .A1(G141), .A2(n907), .ZN(n722) );
  NAND2_X1 U793 ( .A1(n723), .A2(n722), .ZN(n726) );
  NAND2_X1 U794 ( .A1(n908), .A2(G105), .ZN(n724) );
  XOR2_X1 U795 ( .A(KEYINPUT38), .B(n724), .Z(n725) );
  NOR2_X1 U796 ( .A1(n726), .A2(n725), .ZN(n728) );
  NAND2_X1 U797 ( .A1(G117), .A2(n901), .ZN(n727) );
  NAND2_X1 U798 ( .A1(n728), .A2(n727), .ZN(n892) );
  NAND2_X1 U799 ( .A1(G1996), .A2(n892), .ZN(n729) );
  NAND2_X1 U800 ( .A1(n730), .A2(n729), .ZN(n1016) );
  NAND2_X1 U801 ( .A1(n759), .A2(n1016), .ZN(n747) );
  XNOR2_X1 U802 ( .A(G1986), .B(G290), .ZN(n947) );
  NAND2_X1 U803 ( .A1(n759), .A2(n947), .ZN(n731) );
  NAND2_X1 U804 ( .A1(n747), .A2(n731), .ZN(n732) );
  NAND2_X1 U805 ( .A1(G140), .A2(n907), .ZN(n735) );
  NAND2_X1 U806 ( .A1(G104), .A2(n908), .ZN(n734) );
  NAND2_X1 U807 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U808 ( .A(KEYINPUT34), .B(n736), .ZN(n741) );
  NAND2_X1 U809 ( .A1(G128), .A2(n903), .ZN(n738) );
  NAND2_X1 U810 ( .A1(G116), .A2(n901), .ZN(n737) );
  NAND2_X1 U811 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U812 ( .A(n739), .B(KEYINPUT35), .Z(n740) );
  NOR2_X1 U813 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U814 ( .A(KEYINPUT36), .B(n742), .Z(n743) );
  XOR2_X1 U815 ( .A(KEYINPUT88), .B(n743), .Z(n893) );
  XNOR2_X1 U816 ( .A(KEYINPUT37), .B(G2067), .ZN(n746) );
  NOR2_X1 U817 ( .A1(n893), .A2(n746), .ZN(n1021) );
  NAND2_X1 U818 ( .A1(n1021), .A2(n759), .ZN(n754) );
  NAND2_X1 U819 ( .A1(n744), .A2(n754), .ZN(n745) );
  XNOR2_X1 U820 ( .A(KEYINPUT103), .B(n745), .ZN(n762) );
  NAND2_X1 U821 ( .A1(n893), .A2(n746), .ZN(n1019) );
  NOR2_X1 U822 ( .A1(G1996), .A2(n892), .ZN(n1008) );
  INV_X1 U823 ( .A(n747), .ZN(n750) );
  NOR2_X1 U824 ( .A1(G1986), .A2(G290), .ZN(n748) );
  NOR2_X1 U825 ( .A1(G1991), .A2(n898), .ZN(n1012) );
  NOR2_X1 U826 ( .A1(n748), .A2(n1012), .ZN(n749) );
  NOR2_X1 U827 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U828 ( .A1(n1008), .A2(n751), .ZN(n752) );
  XNOR2_X1 U829 ( .A(KEYINPUT104), .B(n752), .ZN(n753) );
  XNOR2_X1 U830 ( .A(n753), .B(KEYINPUT39), .ZN(n755) );
  NAND2_X1 U831 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U832 ( .A1(n1019), .A2(n756), .ZN(n757) );
  XOR2_X1 U833 ( .A(KEYINPUT105), .B(n757), .Z(n758) );
  NAND2_X1 U834 ( .A1(n759), .A2(n758), .ZN(n760) );
  XOR2_X1 U835 ( .A(n760), .B(KEYINPUT106), .Z(n761) );
  NOR2_X1 U836 ( .A1(n762), .A2(n761), .ZN(n764) );
  XNOR2_X1 U837 ( .A(n764), .B(n763), .ZN(G329) );
  AND2_X1 U838 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U839 ( .A(G132), .ZN(G219) );
  INV_X1 U840 ( .A(G120), .ZN(G236) );
  INV_X1 U841 ( .A(G69), .ZN(G235) );
  INV_X1 U842 ( .A(G108), .ZN(G238) );
  NAND2_X1 U843 ( .A1(G7), .A2(G661), .ZN(n765) );
  XNOR2_X1 U844 ( .A(n765), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U845 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n767) );
  INV_X1 U846 ( .A(G223), .ZN(n845) );
  NAND2_X1 U847 ( .A1(G567), .A2(n845), .ZN(n766) );
  XNOR2_X1 U848 ( .A(n767), .B(n766), .ZN(G234) );
  INV_X1 U849 ( .A(G860), .ZN(n775) );
  OR2_X1 U850 ( .A1(n940), .A2(n775), .ZN(G153) );
  XNOR2_X1 U851 ( .A(G171), .B(KEYINPUT75), .ZN(G301) );
  INV_X1 U852 ( .A(G868), .ZN(n815) );
  NAND2_X1 U853 ( .A1(n941), .A2(n815), .ZN(n769) );
  NAND2_X1 U854 ( .A1(G868), .A2(G301), .ZN(n768) );
  NAND2_X1 U855 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U856 ( .A(n770), .B(KEYINPUT76), .ZN(G284) );
  NOR2_X1 U857 ( .A1(G286), .A2(n815), .ZN(n771) );
  XNOR2_X1 U858 ( .A(n771), .B(KEYINPUT79), .ZN(n773) );
  NAND2_X1 U859 ( .A1(n926), .A2(n815), .ZN(n772) );
  NAND2_X1 U860 ( .A1(n773), .A2(n772), .ZN(n774) );
  XOR2_X1 U861 ( .A(KEYINPUT80), .B(n774), .Z(G297) );
  NAND2_X1 U862 ( .A1(n775), .A2(G559), .ZN(n776) );
  INV_X1 U863 ( .A(n941), .ZN(n791) );
  NAND2_X1 U864 ( .A1(n776), .A2(n791), .ZN(n777) );
  XNOR2_X1 U865 ( .A(n777), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U866 ( .A1(G868), .A2(n940), .ZN(n780) );
  NAND2_X1 U867 ( .A1(n791), .A2(G868), .ZN(n778) );
  NOR2_X1 U868 ( .A1(G559), .A2(n778), .ZN(n779) );
  NOR2_X1 U869 ( .A1(n780), .A2(n779), .ZN(G282) );
  NAND2_X1 U870 ( .A1(G123), .A2(n903), .ZN(n781) );
  XNOR2_X1 U871 ( .A(n781), .B(KEYINPUT18), .ZN(n784) );
  NAND2_X1 U872 ( .A1(G135), .A2(n907), .ZN(n782) );
  XOR2_X1 U873 ( .A(KEYINPUT81), .B(n782), .Z(n783) );
  NAND2_X1 U874 ( .A1(n784), .A2(n783), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n908), .A2(G99), .ZN(n786) );
  NAND2_X1 U876 ( .A1(G111), .A2(n901), .ZN(n785) );
  NAND2_X1 U877 ( .A1(n786), .A2(n785), .ZN(n787) );
  NOR2_X1 U878 ( .A1(n788), .A2(n787), .ZN(n1018) );
  XNOR2_X1 U879 ( .A(G2096), .B(n1018), .ZN(n790) );
  INV_X1 U880 ( .A(G2100), .ZN(n789) );
  NAND2_X1 U881 ( .A1(n790), .A2(n789), .ZN(G156) );
  NAND2_X1 U882 ( .A1(n791), .A2(G559), .ZN(n804) );
  XNOR2_X1 U883 ( .A(n940), .B(n804), .ZN(n792) );
  NOR2_X1 U884 ( .A1(n792), .A2(G860), .ZN(n803) );
  NAND2_X1 U885 ( .A1(G67), .A2(n793), .ZN(n796) );
  NAND2_X1 U886 ( .A1(G55), .A2(n794), .ZN(n795) );
  NAND2_X1 U887 ( .A1(n796), .A2(n795), .ZN(n802) );
  NAND2_X1 U888 ( .A1(G80), .A2(n797), .ZN(n800) );
  NAND2_X1 U889 ( .A1(G93), .A2(n798), .ZN(n799) );
  NAND2_X1 U890 ( .A1(n800), .A2(n799), .ZN(n801) );
  NOR2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n814) );
  XNOR2_X1 U892 ( .A(n803), .B(n814), .ZN(G145) );
  XOR2_X1 U893 ( .A(KEYINPUT83), .B(n804), .Z(n812) );
  XNOR2_X1 U894 ( .A(KEYINPUT19), .B(KEYINPUT82), .ZN(n806) );
  XNOR2_X1 U895 ( .A(G288), .B(G166), .ZN(n805) );
  XNOR2_X1 U896 ( .A(n806), .B(n805), .ZN(n807) );
  XNOR2_X1 U897 ( .A(n814), .B(n807), .ZN(n809) );
  XNOR2_X1 U898 ( .A(G305), .B(n926), .ZN(n808) );
  XNOR2_X1 U899 ( .A(n809), .B(n808), .ZN(n810) );
  XOR2_X1 U900 ( .A(G290), .B(n810), .Z(n811) );
  XNOR2_X1 U901 ( .A(n940), .B(n811), .ZN(n872) );
  XNOR2_X1 U902 ( .A(n812), .B(n872), .ZN(n813) );
  NAND2_X1 U903 ( .A1(n813), .A2(G868), .ZN(n817) );
  NAND2_X1 U904 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U905 ( .A1(n817), .A2(n816), .ZN(n818) );
  XOR2_X1 U906 ( .A(KEYINPUT84), .B(n818), .Z(G295) );
  NAND2_X1 U907 ( .A1(G2078), .A2(G2084), .ZN(n819) );
  XOR2_X1 U908 ( .A(KEYINPUT20), .B(n819), .Z(n820) );
  NAND2_X1 U909 ( .A1(G2090), .A2(n820), .ZN(n821) );
  XNOR2_X1 U910 ( .A(KEYINPUT21), .B(n821), .ZN(n822) );
  NAND2_X1 U911 ( .A1(n822), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U912 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  XNOR2_X1 U913 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U914 ( .A1(G235), .A2(G236), .ZN(n823) );
  XNOR2_X1 U915 ( .A(n823), .B(KEYINPUT87), .ZN(n824) );
  NOR2_X1 U916 ( .A1(G238), .A2(n824), .ZN(n825) );
  NAND2_X1 U917 ( .A1(G57), .A2(n825), .ZN(n849) );
  NAND2_X1 U918 ( .A1(n849), .A2(G567), .ZN(n832) );
  NOR2_X1 U919 ( .A1(G219), .A2(G220), .ZN(n827) );
  XNOR2_X1 U920 ( .A(KEYINPUT22), .B(KEYINPUT85), .ZN(n826) );
  XNOR2_X1 U921 ( .A(n827), .B(n826), .ZN(n828) );
  NOR2_X1 U922 ( .A1(n828), .A2(G218), .ZN(n829) );
  NAND2_X1 U923 ( .A1(G96), .A2(n829), .ZN(n830) );
  XNOR2_X1 U924 ( .A(KEYINPUT86), .B(n830), .ZN(n850) );
  NAND2_X1 U925 ( .A1(n850), .A2(G2106), .ZN(n831) );
  NAND2_X1 U926 ( .A1(n832), .A2(n831), .ZN(n851) );
  NAND2_X1 U927 ( .A1(G661), .A2(G483), .ZN(n833) );
  NOR2_X1 U928 ( .A1(n851), .A2(n833), .ZN(n848) );
  NAND2_X1 U929 ( .A1(n848), .A2(G36), .ZN(G176) );
  XNOR2_X1 U930 ( .A(G2427), .B(G2451), .ZN(n843) );
  XOR2_X1 U931 ( .A(G2430), .B(G2443), .Z(n835) );
  XNOR2_X1 U932 ( .A(KEYINPUT109), .B(G2435), .ZN(n834) );
  XNOR2_X1 U933 ( .A(n835), .B(n834), .ZN(n839) );
  XOR2_X1 U934 ( .A(G2438), .B(G2454), .Z(n837) );
  XNOR2_X1 U935 ( .A(G1348), .B(G1341), .ZN(n836) );
  XNOR2_X1 U936 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U937 ( .A(n839), .B(n838), .Z(n841) );
  XNOR2_X1 U938 ( .A(KEYINPUT108), .B(G2446), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n841), .B(n840), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(n844) );
  NAND2_X1 U941 ( .A1(n844), .A2(G14), .ZN(n921) );
  XOR2_X1 U942 ( .A(KEYINPUT110), .B(n921), .Z(G401) );
  NAND2_X1 U943 ( .A1(G2106), .A2(n845), .ZN(G217) );
  AND2_X1 U944 ( .A1(G15), .A2(G2), .ZN(n846) );
  NAND2_X1 U945 ( .A1(G661), .A2(n846), .ZN(G259) );
  NAND2_X1 U946 ( .A1(G3), .A2(G1), .ZN(n847) );
  NAND2_X1 U947 ( .A1(n848), .A2(n847), .ZN(G188) );
  XNOR2_X1 U948 ( .A(G96), .B(KEYINPUT111), .ZN(G221) );
  NOR2_X1 U950 ( .A1(n850), .A2(n849), .ZN(G325) );
  INV_X1 U951 ( .A(G325), .ZN(G261) );
  INV_X1 U952 ( .A(n851), .ZN(G319) );
  XOR2_X1 U953 ( .A(G2096), .B(KEYINPUT43), .Z(n853) );
  XNOR2_X1 U954 ( .A(G2072), .B(KEYINPUT42), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U956 ( .A(n854), .B(G2678), .Z(n856) );
  XNOR2_X1 U957 ( .A(G2067), .B(G2090), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U959 ( .A(KEYINPUT112), .B(G2100), .Z(n858) );
  XNOR2_X1 U960 ( .A(G2078), .B(G2084), .ZN(n857) );
  XNOR2_X1 U961 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U962 ( .A(n860), .B(n859), .ZN(G227) );
  XOR2_X1 U963 ( .A(G1971), .B(G1956), .Z(n862) );
  XNOR2_X1 U964 ( .A(G1986), .B(G1976), .ZN(n861) );
  XNOR2_X1 U965 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U966 ( .A(G1966), .B(G1981), .Z(n864) );
  XNOR2_X1 U967 ( .A(G1991), .B(G1996), .ZN(n863) );
  XNOR2_X1 U968 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U969 ( .A(n866), .B(n865), .Z(n868) );
  XNOR2_X1 U970 ( .A(KEYINPUT113), .B(G2474), .ZN(n867) );
  XNOR2_X1 U971 ( .A(n868), .B(n867), .ZN(n869) );
  XNOR2_X1 U972 ( .A(KEYINPUT41), .B(n869), .ZN(n870) );
  XNOR2_X1 U973 ( .A(n870), .B(n952), .ZN(G229) );
  XOR2_X1 U974 ( .A(G171), .B(G286), .Z(n871) );
  XNOR2_X1 U975 ( .A(n941), .B(n871), .ZN(n873) );
  XNOR2_X1 U976 ( .A(n873), .B(n872), .ZN(n874) );
  NOR2_X1 U977 ( .A1(G37), .A2(n874), .ZN(G397) );
  NAND2_X1 U978 ( .A1(G124), .A2(n903), .ZN(n875) );
  XNOR2_X1 U979 ( .A(n875), .B(KEYINPUT44), .ZN(n876) );
  XNOR2_X1 U980 ( .A(n876), .B(KEYINPUT114), .ZN(n878) );
  NAND2_X1 U981 ( .A1(G100), .A2(n908), .ZN(n877) );
  NAND2_X1 U982 ( .A1(n878), .A2(n877), .ZN(n882) );
  NAND2_X1 U983 ( .A1(n907), .A2(G136), .ZN(n880) );
  NAND2_X1 U984 ( .A1(G112), .A2(n901), .ZN(n879) );
  NAND2_X1 U985 ( .A1(n880), .A2(n879), .ZN(n881) );
  NOR2_X1 U986 ( .A1(n882), .A2(n881), .ZN(G162) );
  NAND2_X1 U987 ( .A1(G139), .A2(n907), .ZN(n884) );
  NAND2_X1 U988 ( .A1(G103), .A2(n908), .ZN(n883) );
  NAND2_X1 U989 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U990 ( .A(KEYINPUT117), .B(n885), .Z(n890) );
  NAND2_X1 U991 ( .A1(G127), .A2(n903), .ZN(n887) );
  NAND2_X1 U992 ( .A1(G115), .A2(n901), .ZN(n886) );
  NAND2_X1 U993 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U994 ( .A(KEYINPUT47), .B(n888), .Z(n889) );
  NOR2_X1 U995 ( .A1(n890), .A2(n889), .ZN(n1003) );
  XOR2_X1 U996 ( .A(G164), .B(n1003), .Z(n891) );
  XNOR2_X1 U997 ( .A(n892), .B(n891), .ZN(n897) );
  XOR2_X1 U998 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n895) );
  XNOR2_X1 U999 ( .A(n893), .B(n1018), .ZN(n894) );
  XNOR2_X1 U1000 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U1001 ( .A(n897), .B(n896), .ZN(n900) );
  XNOR2_X1 U1002 ( .A(n898), .B(G162), .ZN(n899) );
  XNOR2_X1 U1003 ( .A(n900), .B(n899), .ZN(n916) );
  NAND2_X1 U1004 ( .A1(n901), .A2(G118), .ZN(n902) );
  XNOR2_X1 U1005 ( .A(n902), .B(KEYINPUT116), .ZN(n906) );
  NAND2_X1 U1006 ( .A1(G130), .A2(n903), .ZN(n904) );
  XOR2_X1 U1007 ( .A(KEYINPUT115), .B(n904), .Z(n905) );
  NAND2_X1 U1008 ( .A1(n906), .A2(n905), .ZN(n913) );
  NAND2_X1 U1009 ( .A1(G142), .A2(n907), .ZN(n910) );
  NAND2_X1 U1010 ( .A1(G106), .A2(n908), .ZN(n909) );
  NAND2_X1 U1011 ( .A1(n910), .A2(n909), .ZN(n911) );
  XOR2_X1 U1012 ( .A(KEYINPUT45), .B(n911), .Z(n912) );
  NOR2_X1 U1013 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1014 ( .A(G160), .B(n914), .ZN(n915) );
  XNOR2_X1 U1015 ( .A(n916), .B(n915), .ZN(n917) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n917), .ZN(n918) );
  XNOR2_X1 U1017 ( .A(KEYINPUT118), .B(n918), .ZN(G395) );
  NOR2_X1 U1018 ( .A1(G227), .A2(G229), .ZN(n919) );
  XOR2_X1 U1019 ( .A(KEYINPUT49), .B(n919), .Z(n920) );
  NAND2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n924) );
  NOR2_X1 U1021 ( .A1(G397), .A2(G395), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(KEYINPUT119), .B(n922), .ZN(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(G319), .A2(n925), .ZN(G225) );
  INV_X1 U1025 ( .A(G225), .ZN(G308) );
  INV_X1 U1026 ( .A(n926), .ZN(G299) );
  INV_X1 U1027 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1028 ( .A(G16), .B(KEYINPUT56), .ZN(n951) );
  NAND2_X1 U1029 ( .A1(G1971), .A2(G303), .ZN(n927) );
  NAND2_X1 U1030 ( .A1(n928), .A2(n927), .ZN(n934) );
  XOR2_X1 U1031 ( .A(G171), .B(G1961), .Z(n930) );
  XNOR2_X1 U1032 ( .A(G299), .B(G1956), .ZN(n929) );
  NOR2_X1 U1033 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1034 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n949) );
  XNOR2_X1 U1036 ( .A(G1966), .B(G168), .ZN(n935) );
  XNOR2_X1 U1037 ( .A(n935), .B(KEYINPUT124), .ZN(n937) );
  NAND2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n939) );
  XOR2_X1 U1039 ( .A(KEYINPUT125), .B(KEYINPUT57), .Z(n938) );
  XNOR2_X1 U1040 ( .A(n939), .B(n938), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(G1341), .B(n940), .ZN(n943) );
  XNOR2_X1 U1042 ( .A(G1348), .B(n941), .ZN(n942) );
  NOR2_X1 U1043 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n977) );
  INV_X1 U1048 ( .A(G16), .ZN(n975) );
  XNOR2_X1 U1049 ( .A(G5), .B(n952), .ZN(n972) );
  XOR2_X1 U1050 ( .A(G1966), .B(G21), .Z(n962) );
  XNOR2_X1 U1051 ( .A(G1348), .B(KEYINPUT59), .ZN(n953) );
  XNOR2_X1 U1052 ( .A(n953), .B(G4), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(G1981), .B(G6), .ZN(n955) );
  XNOR2_X1 U1054 ( .A(G1341), .B(G19), .ZN(n954) );
  NOR2_X1 U1055 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n959) );
  XNOR2_X1 U1057 ( .A(G20), .B(G1956), .ZN(n958) );
  NOR2_X1 U1058 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1059 ( .A(n960), .B(KEYINPUT60), .ZN(n961) );
  NAND2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1061 ( .A(KEYINPUT126), .B(n963), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(G1976), .B(G23), .ZN(n965) );
  XNOR2_X1 U1063 ( .A(G1971), .B(G22), .ZN(n964) );
  NOR2_X1 U1064 ( .A1(n965), .A2(n964), .ZN(n967) );
  XOR2_X1 U1065 ( .A(G1986), .B(G24), .Z(n966) );
  NAND2_X1 U1066 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1067 ( .A(KEYINPUT58), .B(n968), .ZN(n969) );
  NOR2_X1 U1068 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1070 ( .A(KEYINPUT61), .B(n973), .Z(n974) );
  NAND2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n1001) );
  XOR2_X1 U1073 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n996) );
  XNOR2_X1 U1074 ( .A(G2090), .B(G35), .ZN(n991) );
  XOR2_X1 U1075 ( .A(G1991), .B(G25), .Z(n978) );
  NAND2_X1 U1076 ( .A1(n978), .A2(G28), .ZN(n988) );
  XNOR2_X1 U1077 ( .A(G2067), .B(G26), .ZN(n980) );
  XNOR2_X1 U1078 ( .A(G33), .B(G2072), .ZN(n979) );
  NOR2_X1 U1079 ( .A1(n980), .A2(n979), .ZN(n986) );
  XOR2_X1 U1080 ( .A(n981), .B(G27), .Z(n984) );
  INV_X1 U1081 ( .A(G1996), .ZN(n982) );
  XOR2_X1 U1082 ( .A(n982), .B(G32), .Z(n983) );
  NOR2_X1 U1083 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1084 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1085 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1086 ( .A(KEYINPUT53), .B(n989), .ZN(n990) );
  NOR2_X1 U1087 ( .A1(n991), .A2(n990), .ZN(n994) );
  XOR2_X1 U1088 ( .A(G2084), .B(G34), .Z(n992) );
  XNOR2_X1 U1089 ( .A(KEYINPUT54), .B(n992), .ZN(n993) );
  NAND2_X1 U1090 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1091 ( .A(n996), .B(n995), .ZN(n997) );
  INV_X1 U1092 ( .A(G29), .ZN(n1029) );
  NAND2_X1 U1093 ( .A1(n997), .A2(n1029), .ZN(n998) );
  NAND2_X1 U1094 ( .A1(G11), .A2(n998), .ZN(n999) );
  XOR2_X1 U1095 ( .A(KEYINPUT123), .B(n999), .Z(n1000) );
  NOR2_X1 U1096 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1097 ( .A(n1002), .B(KEYINPUT127), .ZN(n1031) );
  XOR2_X1 U1098 ( .A(G2072), .B(n1003), .Z(n1005) );
  XOR2_X1 U1099 ( .A(G164), .B(G2078), .Z(n1004) );
  NOR2_X1 U1100 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1101 ( .A(KEYINPUT50), .B(n1006), .ZN(n1014) );
  XOR2_X1 U1102 ( .A(G2090), .B(G162), .Z(n1007) );
  NOR2_X1 U1103 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1104 ( .A(KEYINPUT51), .B(n1009), .Z(n1010) );
  XOR2_X1 U1105 ( .A(KEYINPUT120), .B(n1010), .Z(n1011) );
  NOR2_X1 U1106 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1107 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1108 ( .A1(n1016), .A2(n1015), .ZN(n1024) );
  XOR2_X1 U1109 ( .A(G160), .B(G2084), .Z(n1017) );
  NOR2_X1 U1110 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  NAND2_X1 U1111 ( .A1(n1020), .A2(n1019), .ZN(n1022) );
  NOR2_X1 U1112 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1113 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1114 ( .A(KEYINPUT121), .B(n1025), .ZN(n1026) );
  XOR2_X1 U1115 ( .A(KEYINPUT52), .B(n1026), .Z(n1027) );
  NOR2_X1 U1116 ( .A1(KEYINPUT55), .A2(n1027), .ZN(n1028) );
  NOR2_X1 U1117 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NOR2_X1 U1118 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1119 ( .A(KEYINPUT62), .B(n1032), .ZN(G311) );
  INV_X1 U1120 ( .A(G311), .ZN(G150) );
endmodule

