//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 0 0 1 1 1 0 0 0 1 0 0 0 0 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 1 0 1 0 1 0 1 1 1 1 0 1 1 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G116), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT67), .B(G119), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G116), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT5), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n187), .A2(KEYINPUT67), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT67), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G119), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT5), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n192), .A2(new_n194), .A3(new_n195), .A4(G116), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n196), .A2(G113), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT2), .B(G113), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  AOI22_X1  g013(.A1(new_n191), .A2(new_n197), .B1(new_n199), .B2(new_n190), .ZN(new_n200));
  INV_X1    g014(.A(G104), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT77), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT77), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G104), .ZN(new_n204));
  AOI21_X1  g018(.A(G107), .B1(new_n202), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G107), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(G104), .ZN(new_n207));
  OAI21_X1  g021(.A(G101), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT80), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OAI211_X1 g024(.A(KEYINPUT80), .B(G101), .C1(new_n205), .C2(new_n207), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NOR3_X1   g026(.A1(new_n201), .A2(KEYINPUT3), .A3(G107), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n203), .A2(G104), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n201), .A2(KEYINPUT77), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n206), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n213), .B1(new_n216), .B2(KEYINPUT3), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n202), .A2(new_n204), .A3(G107), .ZN(new_n218));
  INV_X1    g032(.A(G101), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n200), .A2(new_n212), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n192), .A2(new_n194), .ZN(new_n225));
  INV_X1    g039(.A(G116), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n224), .B(new_n198), .C1(new_n227), .C2(new_n188), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n199), .B1(new_n190), .B2(KEYINPUT66), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n213), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n218), .B(new_n231), .C1(new_n205), .C2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G101), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n231), .B1(new_n205), .B2(new_n232), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT4), .B1(new_n236), .B2(new_n220), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n230), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n219), .A2(KEYINPUT4), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n233), .A2(KEYINPUT78), .A3(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(KEYINPUT78), .B1(new_n233), .B2(new_n239), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n223), .B1(new_n238), .B2(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(G110), .B(G122), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n223), .B(new_n244), .C1(new_n238), .C2(new_n242), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(KEYINPUT6), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT6), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n243), .A2(new_n249), .A3(new_n245), .ZN(new_n250));
  INV_X1    g064(.A(G146), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G143), .ZN(new_n252));
  INV_X1    g066(.A(G143), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G146), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  XOR2_X1   g069(.A(KEYINPUT65), .B(G128), .Z(new_n256));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n257), .B1(G143), .B2(new_n251), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n255), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n252), .A2(new_n254), .A3(new_n257), .A4(G128), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AND2_X1   g075(.A1(KEYINPUT0), .A2(G128), .ZN(new_n262));
  OR2_X1    g076(.A1(new_n255), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(KEYINPUT0), .A2(G128), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n255), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT75), .B(G125), .ZN(new_n267));
  MUX2_X1   g081(.A(new_n261), .B(new_n266), .S(new_n267), .Z(new_n268));
  INV_X1    g082(.A(G953), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G224), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n268), .B(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n248), .A2(new_n250), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT84), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n248), .A2(KEYINPUT84), .A3(new_n250), .A4(new_n271), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OR3_X1    g090(.A1(new_n261), .A2(KEYINPUT86), .A3(new_n267), .ZN(new_n277));
  INV_X1    g091(.A(new_n266), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n267), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT86), .B1(new_n261), .B2(new_n267), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n270), .A2(KEYINPUT7), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT87), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT7), .B1(new_n270), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n284), .B1(new_n283), .B2(new_n270), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n281), .A2(new_n282), .B1(new_n268), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n212), .A2(new_n222), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n287), .B(new_n200), .ZN(new_n288));
  XNOR2_X1  g102(.A(KEYINPUT85), .B(KEYINPUT8), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n244), .B(new_n289), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n286), .B(new_n247), .C1(new_n288), .C2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G902), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n276), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(G210), .B1(G237), .B2(G902), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT88), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n293), .B1(new_n274), .B2(new_n275), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n296), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n298), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(KEYINPUT88), .A3(new_n296), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G214), .B1(G237), .B2(G902), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT89), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT89), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n302), .A2(new_n303), .A3(new_n308), .A4(new_n305), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G221), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT9), .B(G234), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n311), .B1(new_n313), .B2(new_n292), .ZN(new_n314));
  INV_X1    g128(.A(G469), .ZN(new_n315));
  XNOR2_X1  g129(.A(G110), .B(G140), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n269), .A2(G227), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n316), .B(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT10), .ZN(new_n320));
  INV_X1    g134(.A(G128), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n255), .B1(new_n258), .B2(new_n321), .ZN(new_n322));
  AOI22_X1  g136(.A1(new_n217), .A2(new_n221), .B1(new_n260), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT81), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n212), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n324), .B1(new_n212), .B2(new_n323), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n320), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n212), .A2(KEYINPUT10), .A3(new_n261), .A4(new_n222), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT4), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n329), .B1(new_n217), .B2(new_n221), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n278), .B1(new_n330), .B2(new_n234), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n233), .A2(new_n239), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT78), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n233), .A2(KEYINPUT78), .A3(new_n239), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n331), .A2(new_n336), .A3(KEYINPUT79), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT79), .B1(new_n331), .B2(new_n336), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n327), .B(new_n328), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT82), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT11), .ZN(new_n342));
  INV_X1    g156(.A(G134), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n342), .B1(new_n343), .B2(G137), .ZN(new_n344));
  INV_X1    g158(.A(G137), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(KEYINPUT11), .A3(G134), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n343), .A2(G137), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(KEYINPUT64), .A3(G131), .ZN(new_n349));
  NAND2_X1  g163(.A1(KEYINPUT64), .A2(G131), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n344), .A2(new_n346), .A3(new_n350), .A4(new_n347), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT68), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n349), .A2(KEYINPUT68), .A3(new_n351), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT79), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n266), .B1(new_n235), .B2(new_n237), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n358), .B1(new_n359), .B2(new_n242), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n331), .A2(new_n336), .A3(KEYINPUT79), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n362), .A2(KEYINPUT82), .A3(new_n327), .A4(new_n328), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n341), .A2(new_n357), .A3(new_n363), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n362), .A2(new_n356), .A3(new_n327), .A4(new_n328), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n319), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n319), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n259), .A2(new_n260), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n287), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n369), .B1(new_n325), .B2(new_n326), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n352), .A2(KEYINPUT12), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(KEYINPUT12), .B1(new_n370), .B2(new_n357), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n367), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n315), .B(new_n292), .C1(new_n366), .C2(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n315), .A2(new_n292), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n365), .A2(new_n319), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n365), .B1(new_n374), .B2(new_n373), .ZN(new_n380));
  AOI22_X1  g194(.A1(new_n364), .A2(new_n379), .B1(new_n380), .B2(new_n318), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n378), .B1(new_n381), .B2(G469), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n314), .B1(new_n377), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT83), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI211_X1 g199(.A(KEYINPUT83), .B(new_n314), .C1(new_n377), .C2(new_n382), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT94), .ZN(new_n387));
  NOR2_X1   g201(.A1(G475), .A2(G902), .ZN(new_n388));
  AOI21_X1  g202(.A(KEYINPUT20), .B1(new_n388), .B2(KEYINPUT93), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n389), .B1(KEYINPUT93), .B2(new_n388), .ZN(new_n390));
  NOR2_X1   g204(.A1(G237), .A2(G953), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G214), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n253), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(G143), .A3(G214), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT90), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(KEYINPUT18), .A3(G131), .ZN(new_n398));
  OR2_X1    g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(G125), .B(G140), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n251), .ZN(new_n401));
  NOR2_X1   g215(.A1(G125), .A2(G140), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n402), .B1(new_n267), .B2(G140), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n401), .B1(new_n404), .B2(new_n251), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n396), .A2(new_n398), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n399), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT16), .ZN(new_n408));
  INV_X1    g222(.A(G140), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n267), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  OAI211_X1 g224(.A(G146), .B(new_n410), .C1(new_n403), .C2(new_n408), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT19), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n400), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n413), .B1(new_n404), .B2(new_n412), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n411), .B1(new_n414), .B2(G146), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT91), .B1(new_n395), .B2(G131), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n395), .A2(G131), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT91), .ZN(new_n418));
  INV_X1    g232(.A(G131), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n393), .A2(new_n418), .A3(new_n419), .A4(new_n394), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n416), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n407), .B1(new_n415), .B2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(G113), .B(G122), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n423), .B(new_n201), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT17), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n416), .A2(new_n427), .A3(new_n417), .A4(new_n420), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n410), .B1(new_n403), .B2(new_n408), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n251), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n395), .A2(KEYINPUT17), .A3(G131), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n428), .A2(new_n430), .A3(new_n411), .A4(new_n431), .ZN(new_n432));
  XOR2_X1   g246(.A(new_n424), .B(KEYINPUT92), .Z(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n407), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n390), .B1(new_n426), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n388), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n436), .B1(new_n426), .B2(new_n434), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT20), .ZN(new_n438));
  OAI22_X1  g252(.A1(new_n387), .A2(new_n435), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n435), .A2(new_n387), .ZN(new_n440));
  OR2_X1    g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(G234), .A2(G237), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n442), .A2(G952), .A3(new_n269), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n442), .A2(G902), .A3(G953), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(G898), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n434), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n424), .B1(new_n432), .B2(new_n407), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n292), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT95), .B(G475), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT96), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n226), .A2(G122), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n226), .A2(G122), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n453), .B(new_n454), .C1(new_n455), .C2(KEYINPUT14), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n455), .A2(KEYINPUT14), .ZN(new_n457));
  INV_X1    g271(.A(new_n454), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT96), .B1(new_n454), .B2(KEYINPUT14), .ZN(new_n460));
  OAI211_X1 g274(.A(G107), .B(new_n456), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n458), .A2(new_n455), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n206), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n256), .A2(G143), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n253), .A2(G128), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n464), .A2(new_n343), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n343), .B1(new_n464), .B2(new_n465), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n461), .B(new_n463), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n464), .ZN(new_n470));
  XOR2_X1   g284(.A(new_n465), .B(KEYINPUT13), .Z(new_n471));
  OAI21_X1  g285(.A(G134), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n462), .B(new_n206), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n466), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G217), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n312), .A2(new_n476), .A3(G953), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n469), .A2(new_n474), .A3(new_n477), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n292), .ZN(new_n482));
  INV_X1    g296(.A(G478), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n483), .A2(KEYINPUT15), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n481), .B(new_n292), .C1(KEYINPUT15), .C2(new_n483), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n441), .A2(new_n447), .A3(new_n452), .A4(new_n488), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n385), .A2(new_n386), .A3(new_n489), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n310), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT29), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n354), .A2(new_n266), .A3(new_n355), .ZN(new_n493));
  INV_X1    g307(.A(new_n230), .ZN(new_n494));
  INV_X1    g308(.A(new_n347), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n343), .A2(G137), .ZN(new_n496));
  OAI21_X1  g310(.A(G131), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n261), .B(new_n497), .C1(G131), .C2(new_n348), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n493), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT28), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT28), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n493), .A2(new_n494), .A3(new_n501), .A4(new_n498), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n497), .B1(new_n348), .B2(G131), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n368), .A2(new_n504), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n352), .A2(new_n266), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n230), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  XOR2_X1   g322(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n509));
  NAND2_X1  g323(.A1(new_n391), .A2(G210), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n509), .B(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT26), .B(G101), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n511), .B(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n492), .B1(new_n508), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n493), .A2(KEYINPUT30), .A3(new_n498), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT30), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n516), .B1(new_n505), .B2(new_n506), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(new_n517), .A3(new_n230), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n499), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n519), .A2(KEYINPUT72), .A3(new_n513), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT72), .B1(new_n519), .B2(new_n513), .ZN(new_n521));
  NOR3_X1   g335(.A1(new_n514), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n493), .A2(new_n498), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n503), .B1(new_n494), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n513), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT29), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n292), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(G472), .B1(new_n522), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT71), .B(KEYINPUT32), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n518), .A2(KEYINPUT70), .A3(new_n499), .A4(new_n525), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT31), .ZN(new_n531));
  OR2_X1    g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n531), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n532), .A2(new_n533), .B1(new_n508), .B2(new_n513), .ZN(new_n534));
  NOR2_X1   g348(.A1(G472), .A2(G902), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n529), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n508), .A2(new_n513), .ZN(new_n538));
  INV_X1    g352(.A(new_n533), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n530), .A2(new_n531), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(KEYINPUT32), .A3(new_n535), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n528), .A2(new_n537), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n476), .B1(G234), .B2(new_n292), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT25), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT76), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n189), .A2(G128), .ZN(new_n548));
  OR2_X1    g362(.A1(new_n548), .A2(KEYINPUT73), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n256), .A2(G119), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(KEYINPUT73), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT24), .B(G110), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT23), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n555), .B1(new_n189), .B2(G128), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n556), .B(new_n548), .C1(new_n550), .C2(new_n555), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n554), .B1(G110), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(new_n411), .A3(new_n401), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n430), .A2(new_n411), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT74), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n557), .A2(new_n561), .A3(G110), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n561), .B1(new_n557), .B2(G110), .ZN(new_n563));
  OAI221_X1 g377(.A(new_n560), .B1(new_n553), .B2(new_n552), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT22), .B(G137), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n269), .A2(G221), .A3(G234), .ZN(new_n566));
  XOR2_X1   g380(.A(new_n565), .B(new_n566), .Z(new_n567));
  NAND3_X1  g381(.A1(new_n559), .A2(new_n564), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n567), .B1(new_n559), .B2(new_n564), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n547), .B1(new_n571), .B2(new_n292), .ZN(new_n572));
  INV_X1    g386(.A(new_n547), .ZN(new_n573));
  NOR4_X1   g387(.A1(new_n569), .A2(new_n570), .A3(G902), .A4(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n545), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n545), .A2(G902), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n544), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n491), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(G101), .ZN(G3));
  NAND2_X1  g395(.A1(new_n377), .A2(new_n382), .ZN(new_n582));
  INV_X1    g396(.A(new_n314), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT83), .ZN(new_n585));
  OAI21_X1  g399(.A(G472), .B1(new_n534), .B2(G902), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n586), .B1(new_n534), .B2(new_n536), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(new_n578), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n383), .A2(new_n384), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n585), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT97), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n585), .A2(new_n588), .A3(KEYINPUT97), .A4(new_n589), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT99), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT98), .B1(new_n300), .B2(new_n296), .ZN(new_n596));
  AOI211_X1 g410(.A(new_n297), .B(new_n293), .C1(new_n274), .C2(new_n275), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n305), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n295), .A2(KEYINPUT98), .A3(new_n297), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n595), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n298), .A2(KEYINPUT98), .A3(new_n301), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n596), .A2(new_n597), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n601), .A2(new_n602), .A3(KEYINPUT99), .A4(new_n305), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n452), .B1(new_n439), .B2(new_n440), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n483), .A2(new_n292), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n608), .B1(new_n482), .B2(G478), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n481), .B(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n609), .B1(new_n611), .B2(G478), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n606), .A2(new_n613), .A3(new_n446), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n594), .A2(new_n604), .A3(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT34), .B(G104), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G6));
  AND2_X1   g431(.A1(new_n437), .A2(new_n438), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n437), .A2(new_n438), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  AND4_X1   g435(.A1(new_n447), .A2(new_n621), .A3(new_n452), .A4(new_n487), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n594), .A2(new_n604), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT35), .B(G107), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G9));
  INV_X1    g439(.A(KEYINPUT100), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n559), .A2(new_n626), .A3(new_n564), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n567), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n629), .A2(KEYINPUT36), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n626), .B1(new_n559), .B2(new_n564), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n628), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n631), .B1(new_n628), .B2(new_n632), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n576), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n575), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n587), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n491), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT37), .B(G110), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G12));
  INV_X1    g457(.A(new_n443), .ZN(new_n644));
  INV_X1    g458(.A(new_n444), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n644), .B1(new_n645), .B2(G900), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n452), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n621), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n648), .A2(new_n488), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n543), .A2(new_n638), .A3(new_n649), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n385), .A2(new_n386), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n604), .A2(new_n651), .A3(KEYINPUT101), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n543), .A2(new_n638), .A3(new_n649), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n585), .A2(new_n589), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n600), .A2(new_n603), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G128), .ZN(G30));
  XNOR2_X1  g473(.A(new_n646), .B(KEYINPUT39), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n585), .A2(new_n589), .A3(new_n660), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n661), .A2(KEYINPUT40), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT38), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n304), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n302), .A2(KEYINPUT38), .A3(new_n303), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n519), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n667), .A2(new_n513), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n523), .A2(new_n494), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n499), .A2(new_n513), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n292), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g485(.A(G472), .B1(new_n668), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n537), .A2(new_n542), .A3(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n606), .A2(new_n488), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n639), .A2(new_n305), .A3(new_n673), .A4(new_n674), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n662), .A2(new_n666), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n676), .B1(KEYINPUT40), .B2(new_n661), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G143), .ZN(G45));
  NAND3_X1  g492(.A1(new_n605), .A2(new_n612), .A3(new_n646), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n543), .A2(new_n638), .A3(new_n680), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n385), .A2(new_n386), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n604), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G146), .ZN(G48));
  NOR2_X1   g498(.A1(new_n366), .A2(new_n376), .ZN(new_n685));
  OAI21_X1  g499(.A(G469), .B1(new_n685), .B2(G902), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n583), .A3(new_n377), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n687), .A2(new_n544), .A3(new_n578), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n688), .A2(new_n600), .A3(new_n603), .A4(new_n614), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT41), .B(G113), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G15));
  NAND4_X1  g505(.A1(new_n688), .A2(new_n600), .A3(new_n603), .A4(new_n622), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G116), .ZN(G18));
  NOR3_X1   g507(.A1(new_n544), .A2(new_n489), .A3(new_n639), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n686), .A2(new_n583), .A3(new_n377), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n694), .A2(new_n600), .A3(new_n603), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT102), .B(G119), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G21));
  AND2_X1   g512(.A1(new_n575), .A2(new_n577), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n524), .A2(new_n513), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n700), .B1(new_n539), .B2(new_n540), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n535), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n699), .A2(new_n586), .A3(new_n702), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n687), .A2(new_n703), .A3(new_n446), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n704), .A2(new_n600), .A3(new_n603), .A4(new_n674), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G122), .ZN(G24));
  NAND3_X1  g520(.A1(new_n638), .A2(new_n586), .A3(new_n702), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT103), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n679), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n605), .A2(new_n612), .A3(KEYINPUT103), .A4(new_n646), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  AND4_X1   g526(.A1(new_n600), .A2(new_n712), .A3(new_n695), .A4(new_n603), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT104), .B(G125), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G27));
  AOI21_X1  g529(.A(new_n306), .B1(new_n302), .B2(new_n303), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n579), .A2(new_n716), .A3(new_n383), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n711), .A2(KEYINPUT42), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n528), .A2(new_n542), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT32), .B1(new_n541), .B2(new_n535), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n721), .A2(new_n711), .A3(new_n578), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(new_n716), .A3(new_n383), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n717), .A2(new_n718), .B1(new_n723), .B2(KEYINPUT42), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G131), .ZN(G33));
  NAND4_X1  g539(.A1(new_n579), .A2(new_n716), .A3(new_n383), .A4(new_n649), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G134), .ZN(G36));
  NAND3_X1  g541(.A1(new_n441), .A2(new_n452), .A3(new_n612), .ZN(new_n728));
  XOR2_X1   g542(.A(new_n728), .B(KEYINPUT43), .Z(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n587), .A3(new_n638), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n716), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n732), .B1(KEYINPUT105), .B2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n377), .ZN(new_n735));
  OR2_X1    g549(.A1(new_n381), .A2(KEYINPUT45), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n381), .A2(KEYINPUT45), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n736), .A2(G469), .A3(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n378), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT46), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n735), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n742), .B1(new_n741), .B2(new_n740), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n743), .A2(new_n583), .A3(new_n660), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n734), .B(new_n744), .C1(KEYINPUT105), .C2(new_n733), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G137), .ZN(G39));
  NAND4_X1  g560(.A1(new_n716), .A2(new_n544), .A3(new_n578), .A4(new_n680), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n743), .A2(KEYINPUT47), .A3(new_n583), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(KEYINPUT47), .B1(new_n743), .B2(new_n583), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n748), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G140), .ZN(G42));
  INV_X1    g567(.A(G952), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n269), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n729), .A2(new_n443), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n703), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(new_n604), .A3(new_n695), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n695), .A2(new_n716), .ZN(new_n759));
  NOR4_X1   g573(.A1(new_n759), .A2(new_n578), .A3(new_n644), .A4(new_n673), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n606), .A2(new_n613), .ZN(new_n761));
  AOI211_X1 g575(.A(new_n754), .B(G953), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n759), .A2(new_n756), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT112), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n763), .B(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT48), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n721), .A2(new_n578), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n766), .B1(new_n765), .B2(new_n767), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n758), .B(new_n762), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n743), .A2(new_n583), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT47), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n686), .A2(new_n377), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n314), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n774), .A2(new_n749), .A3(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n716), .A3(new_n757), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n687), .A2(new_n305), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n779), .B1(new_n666), .B2(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n780), .A2(new_n664), .A3(new_n779), .A4(new_n665), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n757), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n784));
  OR3_X1    g598(.A1(new_n781), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n784), .B1(new_n781), .B2(new_n783), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n707), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n606), .A2(new_n613), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  AOI22_X1  g604(.A1(new_n765), .A2(new_n788), .B1(new_n760), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n778), .A2(new_n787), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n770), .B1(new_n771), .B2(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n778), .A2(new_n787), .A3(new_n791), .A4(KEYINPUT51), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n794), .A2(KEYINPUT113), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(KEYINPUT113), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n793), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT114), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n793), .B(new_n799), .C1(new_n795), .C2(new_n796), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n592), .A2(new_n310), .A3(new_n593), .A4(new_n614), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n487), .B(KEYINPUT108), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n803), .A2(new_n446), .A3(new_n605), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n592), .A2(new_n310), .A3(new_n593), .A4(new_n804), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n310), .B(new_n490), .C1(new_n579), .C2(new_n640), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT108), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n487), .B(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(KEYINPUT109), .B1(new_n808), .B2(new_n648), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT109), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n803), .A2(new_n810), .A3(new_n621), .A4(new_n647), .ZN(new_n811));
  AND4_X1   g625(.A1(new_n543), .A2(new_n809), .A3(new_n811), .A4(new_n638), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(new_n585), .A3(new_n589), .A4(new_n716), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n712), .A2(new_n716), .A3(new_n383), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n813), .A2(new_n726), .A3(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n802), .A2(new_n805), .A3(new_n806), .A4(new_n815), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n604), .B(new_n688), .C1(new_n614), .C2(new_n622), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n724), .A2(new_n817), .A3(new_n696), .A4(new_n705), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n713), .B1(new_n652), .B2(new_n657), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n600), .A2(new_n603), .A3(new_n674), .ZN(new_n821));
  AND4_X1   g635(.A1(new_n383), .A2(new_n639), .A3(new_n646), .A4(new_n673), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n821), .A2(new_n822), .B1(new_n604), .B2(new_n682), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n820), .A2(KEYINPUT52), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT52), .B1(new_n820), .B2(new_n823), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n819), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(KEYINPUT54), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n827), .A2(new_n828), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n832));
  INV_X1    g646(.A(new_n713), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n658), .A2(new_n823), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT52), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n824), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n816), .A2(new_n828), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT110), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n705), .A2(new_n689), .A3(new_n692), .A4(new_n696), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n717), .A2(new_n718), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n723), .A2(KEYINPUT42), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n839), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n705), .A2(new_n696), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(KEYINPUT110), .A3(new_n724), .A4(new_n817), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n837), .A2(new_n838), .A3(new_n844), .A4(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n831), .A2(new_n832), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n830), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n755), .B1(new_n801), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n699), .A2(new_n305), .A3(new_n583), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n606), .B(new_n612), .C1(new_n851), .C2(KEYINPUT106), .ZN(new_n852));
  AOI211_X1 g666(.A(new_n673), .B(new_n852), .C1(KEYINPUT106), .C2(new_n851), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n775), .B(KEYINPUT49), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n853), .A2(new_n854), .A3(new_n666), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT107), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n850), .A2(new_n856), .ZN(G75));
  NOR2_X1   g671(.A1(new_n269), .A2(G952), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n292), .B1(new_n831), .B2(new_n847), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n860), .A2(G210), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n248), .A2(new_n250), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(KEYINPUT115), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n271), .B(KEYINPUT55), .Z(new_n864));
  XNOR2_X1  g678(.A(new_n863), .B(new_n864), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n865), .A2(KEYINPUT56), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n859), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n860), .A2(G210), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT116), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT56), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n870), .B1(new_n869), .B2(new_n868), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n867), .B1(new_n871), .B2(new_n865), .ZN(G51));
  INV_X1    g686(.A(new_n738), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n825), .A2(new_n826), .ZN(new_n874));
  AND4_X1   g688(.A1(new_n802), .A2(new_n805), .A3(new_n806), .A4(new_n815), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n875), .A2(new_n844), .A3(KEYINPUT53), .A4(new_n846), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT53), .B1(new_n837), .B2(new_n819), .ZN(new_n878));
  OAI211_X1 g692(.A(G902), .B(new_n873), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT118), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n831), .A2(new_n847), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(KEYINPUT118), .A3(G902), .A4(new_n873), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(KEYINPUT54), .B1(new_n877), .B2(new_n878), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n848), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n378), .B(KEYINPUT57), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n685), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT117), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n884), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n887), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(new_n885), .B2(new_n848), .ZN(new_n892));
  OAI21_X1  g706(.A(KEYINPUT117), .B1(new_n892), .B2(new_n685), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n858), .B1(new_n890), .B2(new_n893), .ZN(G54));
  NAND3_X1  g708(.A1(new_n860), .A2(KEYINPUT58), .A3(G475), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n426), .A2(new_n434), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n895), .A2(new_n897), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n898), .A2(new_n899), .A3(new_n858), .ZN(G60));
  INV_X1    g714(.A(new_n611), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n607), .B(KEYINPUT59), .Z(new_n902));
  AOI21_X1  g716(.A(new_n901), .B1(new_n849), .B2(new_n902), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n886), .A2(new_n901), .A3(new_n902), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n903), .A2(new_n858), .A3(new_n904), .ZN(G63));
  NAND2_X1  g719(.A1(G217), .A2(G902), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT60), .Z(new_n907));
  NAND2_X1  g721(.A1(new_n882), .A2(new_n907), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n571), .B(KEYINPUT119), .Z(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n910), .B(new_n859), .C1(new_n636), .C2(new_n908), .ZN(new_n911));
  XNOR2_X1  g725(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OR2_X1    g727(.A1(new_n908), .A2(new_n636), .ZN(new_n914));
  OR2_X1    g728(.A1(KEYINPUT120), .A2(KEYINPUT61), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n914), .A2(new_n859), .A3(new_n910), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n913), .A2(new_n916), .ZN(G66));
  INV_X1    g731(.A(G224), .ZN(new_n918));
  OAI21_X1  g732(.A(G953), .B1(new_n445), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n802), .A2(new_n805), .A3(new_n806), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n920), .A2(new_n840), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n919), .B1(new_n921), .B2(G953), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n863), .B1(G898), .B2(new_n269), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n922), .B(new_n923), .ZN(G69));
  NAND2_X1  g738(.A1(new_n515), .A2(new_n517), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n414), .B(KEYINPUT121), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n761), .B1(new_n606), .B2(new_n808), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT123), .Z(new_n929));
  NAND3_X1  g743(.A1(new_n929), .A2(new_n579), .A3(new_n716), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n745), .B(new_n752), .C1(new_n661), .C2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n820), .A2(new_n683), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT122), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n820), .A2(KEYINPUT122), .A3(new_n683), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n934), .A2(new_n677), .A3(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT62), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n934), .A2(KEYINPUT62), .A3(new_n677), .A4(new_n935), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n931), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n927), .B1(new_n940), .B2(G953), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n744), .A2(new_n821), .A3(new_n767), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n724), .A2(new_n726), .ZN(new_n943));
  AND4_X1   g757(.A1(new_n745), .A2(new_n752), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n944), .A2(new_n269), .A3(new_n934), .A4(new_n935), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n927), .B1(G900), .B2(G953), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n269), .B1(G227), .B2(G900), .ZN(new_n947));
  AOI22_X1  g761(.A1(new_n945), .A2(new_n946), .B1(KEYINPUT124), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n941), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n947), .A2(KEYINPUT124), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n949), .B(new_n950), .Z(G72));
  NAND2_X1  g765(.A1(new_n940), .A2(new_n921), .ZN(new_n952));
  XOR2_X1   g766(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n953));
  NAND2_X1  g767(.A1(G472), .A2(G902), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT126), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n668), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT127), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n520), .A2(new_n521), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(new_n513), .B2(new_n519), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n829), .A2(new_n955), .A3(new_n961), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n944), .A2(new_n921), .A3(new_n934), .A4(new_n935), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n956), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n519), .A2(new_n525), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n858), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n958), .A2(new_n959), .A3(new_n962), .A4(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n962), .ZN(new_n968));
  INV_X1    g782(.A(new_n668), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n952), .B2(new_n956), .ZN(new_n970));
  OAI21_X1  g784(.A(KEYINPUT127), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n967), .A2(new_n971), .ZN(G57));
endmodule


