//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 0 1 1 0 1 0 0 0 1 1 1 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 0 1 0 0 1 1 0 1 0 0 1 1 1 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n815, new_n816, new_n817, new_n818, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n983, new_n984, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1037, new_n1038,
    new_n1039;
  INV_X1    g000(.A(G43gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(G50gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(G50gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n204), .A2(KEYINPUT15), .A3(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT15), .ZN(new_n208));
  OR2_X1    g007(.A1(KEYINPUT88), .A2(G50gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(KEYINPUT88), .A2(G50gat), .ZN(new_n210));
  AOI21_X1  g009(.A(G43gat), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n208), .B1(new_n211), .B2(new_n203), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT14), .B(G29gat), .ZN(new_n213));
  INV_X1    g012(.A(G36gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT14), .ZN(new_n216));
  NOR3_X1   g015(.A1(new_n216), .A2(new_n214), .A3(G29gat), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n207), .B1(new_n212), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n217), .B1(new_n214), .B2(new_n213), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(new_n206), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT17), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G15gat), .B(G22gat), .ZN(new_n224));
  INV_X1    g023(.A(G1gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT16), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(G1gat), .B2(new_n224), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G8gat), .ZN(new_n229));
  INV_X1    g028(.A(G8gat), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n227), .B(new_n230), .C1(G1gat), .C2(new_n224), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n210), .ZN(new_n234));
  NOR2_X1   g033(.A1(KEYINPUT88), .A2(G50gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n202), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT15), .B1(new_n236), .B2(new_n204), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n206), .B1(new_n237), .B2(new_n221), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT17), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n219), .A2(new_n207), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n223), .A2(new_n233), .A3(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n220), .A2(new_n222), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(new_n232), .ZN(new_n244));
  NAND2_X1  g043(.A1(G229gat), .A2(G233gat), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n242), .A2(KEYINPUT18), .A3(new_n244), .A4(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n245), .B(KEYINPUT13), .Z(new_n247));
  NOR2_X1   g046(.A1(new_n243), .A2(new_n232), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n232), .A2(new_n238), .A3(new_n240), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G113gat), .B(G141gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(G197gat), .ZN(new_n254));
  XOR2_X1   g053(.A(KEYINPUT11), .B(G169gat), .Z(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(KEYINPUT12), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n242), .A2(new_n244), .A3(new_n245), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT90), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT18), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n259), .B1(new_n258), .B2(new_n260), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n252), .B(new_n257), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT89), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n246), .A2(new_n250), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n264), .B1(new_n246), .B2(new_n250), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n258), .A2(new_n260), .ZN(new_n267));
  NOR3_X1   g066(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n263), .B1(new_n268), .B2(new_n257), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G78gat), .B(G106gat), .ZN(new_n271));
  INV_X1    g070(.A(G50gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(G22gat), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(G228gat), .A2(G233gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(G155gat), .A2(G162gat), .ZN(new_n278));
  OR2_X1    g077(.A1(G155gat), .A2(G162gat), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n278), .B1(new_n279), .B2(KEYINPUT2), .ZN(new_n280));
  AND2_X1   g079(.A1(G141gat), .A2(G148gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(G141gat), .A2(G148gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT77), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n280), .A2(new_n283), .A3(KEYINPUT77), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT75), .B1(new_n281), .B2(new_n282), .ZN(new_n289));
  INV_X1    g088(.A(G141gat), .ZN(new_n290));
  INV_X1    g089(.A(G148gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT75), .ZN(new_n293));
  NAND2_X1  g092(.A1(G141gat), .A2(G148gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT2), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n289), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT76), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n279), .A2(new_n278), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n298), .B1(new_n297), .B2(new_n299), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n288), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G211gat), .ZN(new_n304));
  INV_X1    g103(.A(G218gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G211gat), .A2(G218gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT72), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n306), .A2(new_n310), .A3(new_n307), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G197gat), .B(G204gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT22), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n307), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n309), .A2(new_n316), .A3(new_n311), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT29), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT82), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT3), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT29), .B1(new_n318), .B2(new_n319), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT82), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n303), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT3), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n288), .B(new_n328), .C1(new_n300), .C2(new_n301), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n320), .B1(new_n329), .B2(new_n321), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n277), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n320), .A2(KEYINPUT81), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT81), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n321), .B1(new_n318), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n328), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n277), .B1(new_n335), .B2(new_n302), .ZN(new_n336));
  INV_X1    g135(.A(new_n330), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n331), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n340), .B1(new_n331), .B2(new_n338), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n275), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n336), .A2(new_n337), .ZN(new_n344));
  INV_X1    g143(.A(new_n326), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n328), .B1(new_n325), .B2(KEYINPUT82), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n302), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n276), .B1(new_n347), .B2(new_n337), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n339), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n331), .A2(new_n338), .A3(new_n340), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(new_n350), .A3(new_n274), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n343), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n302), .A2(KEYINPUT3), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT1), .ZN(new_n354));
  XNOR2_X1  g153(.A(G127gat), .B(G134gat), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT70), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(G134gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(G127gat), .ZN(new_n359));
  INV_X1    g158(.A(G127gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(G134gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n362), .A2(KEYINPUT70), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n357), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(G113gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(G120gat), .ZN(new_n366));
  XOR2_X1   g165(.A(KEYINPUT69), .B(G120gat), .Z(new_n367));
  OAI21_X1  g166(.A(new_n366), .B1(new_n367), .B2(new_n365), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G120gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(G113gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT68), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n366), .A2(new_n371), .A3(KEYINPUT68), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n374), .A2(new_n354), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n362), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n369), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n353), .A2(new_n329), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(G225gat), .A2(G233gat), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n381), .B1(new_n302), .B2(new_n378), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n297), .A2(new_n299), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT76), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI22_X1  g185(.A1(new_n364), .A2(new_n368), .B1(new_n376), .B2(new_n362), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n386), .A2(KEYINPUT4), .A3(new_n288), .A4(new_n387), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n379), .A2(new_n380), .A3(new_n382), .A4(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT5), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n302), .A2(new_n378), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n386), .A2(new_n288), .A3(new_n387), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n380), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n390), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n389), .A2(new_n395), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n382), .A2(new_n388), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n397), .A2(new_n390), .A3(new_n380), .A4(new_n379), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  XOR2_X1   g198(.A(G1gat), .B(G29gat), .Z(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G57gat), .B(G85gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n399), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT6), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  AND2_X1   g208(.A1(new_n396), .A2(new_n398), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT6), .B1(new_n410), .B2(new_n404), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n406), .A2(KEYINPUT79), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n406), .A2(KEYINPUT79), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n409), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT30), .ZN(new_n416));
  NAND2_X1  g215(.A1(G169gat), .A2(G176gat), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT66), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(G169gat), .ZN(new_n422));
  INV_X1    g221(.A(G176gat), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT23), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT23), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n425), .B1(G169gat), .B2(G176gat), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n421), .A2(KEYINPUT25), .A3(new_n424), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(G183gat), .A2(G190gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT24), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT24), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n430), .A2(G183gat), .A3(G190gat), .ZN(new_n431));
  INV_X1    g230(.A(G183gat), .ZN(new_n432));
  INV_X1    g231(.A(G190gat), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n429), .A2(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT67), .B1(new_n427), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n429), .A2(new_n431), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n436), .B1(G183gat), .B2(G190gat), .ZN(new_n437));
  AND3_X1   g236(.A1(new_n424), .A2(new_n426), .A3(KEYINPUT25), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT67), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n437), .A2(new_n438), .A3(new_n439), .A4(new_n421), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT25), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT65), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n443), .A2(new_n432), .A3(new_n433), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n442), .A2(new_n444), .B1(new_n429), .B2(new_n431), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n424), .A2(new_n426), .A3(new_n417), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n441), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n435), .A2(new_n440), .A3(new_n447), .ZN(new_n448));
  NOR3_X1   g247(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n417), .ZN(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT27), .B(G183gat), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n452), .A2(KEYINPUT28), .A3(new_n433), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT28), .B1(new_n452), .B2(new_n433), .ZN(new_n454));
  OAI221_X1 g253(.A(new_n428), .B1(new_n449), .B2(new_n451), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n448), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(G226gat), .A2(G233gat), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT29), .B1(new_n448), .B2(new_n455), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n459), .B(new_n320), .C1(new_n458), .C2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT74), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n456), .A2(new_n321), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n457), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT74), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n464), .A2(new_n465), .A3(new_n320), .A4(new_n459), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n460), .A2(new_n458), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n459), .A2(KEYINPUT73), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT73), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n456), .A2(new_n469), .A3(new_n458), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n467), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n462), .B(new_n466), .C1(new_n471), .C2(new_n320), .ZN(new_n472));
  XNOR2_X1  g271(.A(G8gat), .B(G36gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(G64gat), .B(G92gat), .ZN(new_n474));
  XOR2_X1   g273(.A(new_n473), .B(new_n474), .Z(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n416), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n472), .A2(new_n476), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n469), .B1(new_n456), .B2(new_n458), .ZN(new_n479));
  AOI211_X1 g278(.A(KEYINPUT73), .B(new_n457), .C1(new_n448), .C2(new_n455), .ZN(new_n480));
  OAI22_X1  g279(.A1(new_n479), .A2(new_n480), .B1(new_n458), .B2(new_n460), .ZN(new_n481));
  INV_X1    g280(.A(new_n320), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n481), .A2(new_n482), .B1(new_n461), .B2(KEYINPUT74), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n483), .A2(KEYINPUT30), .A3(new_n475), .A4(new_n466), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n477), .A2(new_n478), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n352), .B1(new_n415), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n456), .A2(new_n387), .ZN(new_n488));
  NAND2_X1  g287(.A1(G227gat), .A2(G233gat), .ZN(new_n489));
  XOR2_X1   g288(.A(new_n489), .B(KEYINPUT64), .Z(new_n490));
  NAND3_X1  g289(.A1(new_n378), .A2(new_n448), .A3(new_n455), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n488), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT33), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  XOR2_X1   g293(.A(G15gat), .B(G43gat), .Z(new_n495));
  XNOR2_X1  g294(.A(G71gat), .B(G99gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n495), .B(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT34), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n488), .A2(new_n491), .ZN(new_n500));
  INV_X1    g299(.A(new_n490), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n500), .A2(new_n499), .A3(new_n501), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n498), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n497), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n506), .B1(new_n492), .B2(new_n493), .ZN(new_n507));
  INV_X1    g306(.A(new_n504), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n507), .B1(new_n508), .B2(new_n502), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n492), .A2(KEYINPUT32), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n505), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n511), .B1(new_n505), .B2(new_n509), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT71), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT36), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n505), .A2(new_n509), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n510), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n512), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n516), .A2(new_n517), .ZN(new_n522));
  NAND2_X1  g321(.A1(KEYINPUT71), .A2(KEYINPUT36), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n487), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n472), .A2(new_n476), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n472), .A2(KEYINPUT37), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n475), .B1(new_n483), .B2(new_n466), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT37), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n475), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n528), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n527), .B1(new_n532), .B2(KEYINPUT38), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT84), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n399), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n396), .A2(new_n398), .A3(KEYINPUT84), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n535), .A2(new_n405), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n408), .B1(new_n411), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT86), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT38), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n540), .B(new_n476), .C1(new_n472), .C2(KEYINPUT37), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n464), .B(new_n320), .C1(new_n479), .C2(new_n480), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n464), .A2(new_n459), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n542), .A2(KEYINPUT85), .B1(new_n482), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n468), .A2(new_n470), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT85), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n545), .A2(new_n546), .A3(new_n320), .A4(new_n464), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n530), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n539), .B1(new_n541), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n531), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n478), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n542), .A2(KEYINPUT85), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n543), .A2(new_n482), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(new_n547), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT37), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n551), .A2(KEYINPUT86), .A3(new_n540), .A4(new_n555), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n533), .A2(new_n538), .A3(new_n549), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n343), .A2(new_n351), .ZN(new_n558));
  XOR2_X1   g357(.A(KEYINPUT83), .B(KEYINPUT39), .Z(new_n559));
  INV_X1    g358(.A(new_n379), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n382), .A2(new_n388), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n394), .B(new_n559), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n380), .B1(new_n397), .B2(new_n379), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n391), .A2(new_n392), .A3(new_n380), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT39), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n562), .B(new_n404), .C1(new_n563), .C2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT40), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n394), .B1(new_n560), .B2(new_n561), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n569), .A2(KEYINPUT39), .A3(new_n564), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n570), .A2(KEYINPUT40), .A3(new_n404), .A4(new_n562), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  AND3_X1   g371(.A1(new_n396), .A2(KEYINPUT84), .A3(new_n398), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT84), .B1(new_n396), .B2(new_n398), .ZN(new_n574));
  NOR3_X1   g373(.A1(new_n573), .A2(new_n574), .A3(new_n404), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n558), .B1(new_n576), .B2(new_n485), .ZN(new_n577));
  AND3_X1   g376(.A1(new_n557), .A2(KEYINPUT87), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT87), .B1(new_n557), .B2(new_n577), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n526), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n515), .A2(new_n352), .A3(new_n486), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n407), .B1(new_n399), .B2(new_n405), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n582), .B1(KEYINPUT79), .B2(new_n406), .ZN(new_n583));
  INV_X1    g382(.A(new_n414), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n408), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(KEYINPUT35), .B1(new_n581), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT35), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n574), .A2(new_n404), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n582), .B1(new_n588), .B2(new_n536), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n587), .B1(new_n589), .B2(new_n408), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NOR3_X1   g390(.A1(new_n521), .A2(new_n558), .A3(new_n485), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n586), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n270), .B1(new_n580), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT94), .ZN(new_n596));
  INV_X1    g395(.A(G64gat), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n597), .A2(G57gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(G57gat), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT9), .ZN(new_n600));
  NAND2_X1  g399(.A1(G71gat), .A2(G78gat), .ZN(new_n601));
  AOI22_X1  g400(.A1(new_n598), .A2(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT91), .B1(G71gat), .B2(G78gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(new_n601), .ZN(new_n604));
  NAND3_X1  g403(.A1(KEYINPUT91), .A2(G71gat), .A3(G78gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT92), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n604), .A2(KEYINPUT92), .A3(new_n605), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n602), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OR2_X1    g409(.A1(G71gat), .A2(G78gat), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n602), .A2(new_n601), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT93), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n599), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n601), .A2(new_n600), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n604), .A2(KEYINPUT92), .A3(new_n605), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT92), .B1(new_n604), .B2(new_n605), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT93), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n602), .A2(new_n601), .A3(new_n611), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n613), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT21), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n596), .B1(new_n624), .B2(new_n233), .ZN(new_n625));
  AOI211_X1 g424(.A(KEYINPUT94), .B(new_n232), .C1(new_n623), .C2(KEYINPUT21), .ZN(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n627));
  INV_X1    g426(.A(G155gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  OR3_X1    g428(.A1(new_n625), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n629), .B1(new_n625), .B2(new_n626), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(G183gat), .B(G211gat), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n620), .B1(new_n619), .B2(new_n621), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT21), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AND2_X1   g438(.A1(G231gat), .A2(G233gat), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n360), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n641), .A2(new_n360), .A3(new_n642), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n634), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n645), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n647), .A2(new_n643), .A3(new_n633), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n632), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n633), .B1(new_n647), .B2(new_n643), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n644), .A2(new_n634), .A3(new_n645), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n650), .A2(new_n651), .A3(new_n630), .A4(new_n631), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT7), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(KEYINPUT97), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT97), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(KEYINPUT7), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n654), .A2(new_n656), .A3(G85gat), .A4(G92gat), .ZN(new_n657));
  INV_X1    g456(.A(G85gat), .ZN(new_n658));
  INV_X1    g457(.A(G92gat), .ZN(new_n659));
  OAI211_X1 g458(.A(KEYINPUT97), .B(new_n653), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(G99gat), .A2(G106gat), .ZN(new_n661));
  AOI22_X1  g460(.A1(KEYINPUT8), .A2(new_n661), .B1(new_n658), .B2(new_n659), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n657), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(G99gat), .ZN(new_n664));
  INV_X1    g463(.A(G106gat), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n663), .A2(new_n661), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n661), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n657), .A2(new_n668), .A3(new_n660), .A4(new_n662), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  AND2_X1   g470(.A1(G232gat), .A2(G233gat), .ZN(new_n672));
  AOI22_X1  g471(.A1(new_n243), .A2(new_n671), .B1(KEYINPUT41), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n223), .A2(new_n241), .A3(new_n670), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(G190gat), .B(G218gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n676), .B(new_n677), .Z(new_n678));
  XOR2_X1   g477(.A(new_n675), .B(new_n678), .Z(new_n679));
  XOR2_X1   g478(.A(G134gat), .B(G162gat), .Z(new_n680));
  NOR2_X1   g479(.A1(new_n672), .A2(KEYINPUT41), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g481(.A(KEYINPUT95), .B(KEYINPUT96), .Z(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n679), .B(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n649), .A2(new_n652), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(KEYINPUT100), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT100), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n649), .A2(new_n652), .A3(new_n688), .A4(new_n685), .ZN(new_n689));
  AND4_X1   g488(.A1(new_n619), .A2(new_n667), .A3(new_n621), .A4(new_n669), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n690), .B1(new_n623), .B2(new_n670), .ZN(new_n691));
  NAND2_X1  g490(.A1(G230gat), .A2(G233gat), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(G120gat), .B(G148gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(G176gat), .B(G204gat), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n695), .B(new_n696), .Z(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n670), .B1(new_n635), .B2(new_n636), .ZN(new_n700));
  INV_X1    g499(.A(new_n690), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT10), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n623), .A2(KEYINPUT10), .A3(new_n671), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n692), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(KEYINPUT101), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n623), .A2(KEYINPUT10), .A3(new_n671), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(new_n691), .B2(KEYINPUT10), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT101), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n708), .A2(new_n709), .A3(new_n692), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n694), .B1(new_n706), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n705), .B1(new_n711), .B2(new_n697), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n595), .A2(new_n687), .A3(new_n689), .A4(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n714), .A2(new_n415), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(new_n225), .ZN(G1324gat));
  OR2_X1    g515(.A1(new_n714), .A2(new_n486), .ZN(new_n717));
  XOR2_X1   g516(.A(KEYINPUT16), .B(G8gat), .Z(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  AOI22_X1  g519(.A1(new_n720), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n717), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n717), .A2(new_n719), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT42), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n722), .A2(KEYINPUT102), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(KEYINPUT102), .B1(new_n722), .B2(new_n723), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n721), .B1(new_n724), .B2(new_n725), .ZN(G1325gat));
  INV_X1    g525(.A(new_n525), .ZN(new_n727));
  OAI21_X1  g526(.A(G15gat), .B1(new_n714), .B2(new_n727), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n521), .A2(G15gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n714), .B2(new_n729), .ZN(G1326gat));
  NOR2_X1   g529(.A1(new_n714), .A2(new_n352), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT103), .ZN(new_n732));
  XNOR2_X1  g531(.A(KEYINPUT43), .B(G22gat), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1327gat));
  NAND2_X1  g533(.A1(new_n580), .A2(KEYINPUT105), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n587), .B1(new_n592), .B2(new_n415), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n581), .A2(new_n590), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n586), .A2(new_n593), .A3(KEYINPUT106), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT105), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n742), .B(new_n526), .C1(new_n578), .C2(new_n579), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n735), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n685), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT44), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n747));
  AOI211_X1 g546(.A(new_n747), .B(new_n685), .C1(new_n580), .C2(new_n594), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n649), .A2(new_n652), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n712), .B(KEYINPUT104), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n751), .A2(new_n752), .A3(new_n270), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(G29gat), .B1(new_n754), .B2(new_n415), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n751), .A2(new_n685), .A3(new_n712), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n595), .A2(new_n756), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n757), .A2(G29gat), .A3(new_n415), .ZN(new_n758));
  XOR2_X1   g557(.A(new_n758), .B(KEYINPUT45), .Z(new_n759));
  NAND2_X1  g558(.A1(new_n755), .A2(new_n759), .ZN(G1328gat));
  OAI21_X1  g559(.A(G36gat), .B1(new_n754), .B2(new_n486), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n757), .A2(G36gat), .A3(new_n486), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT46), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(G1329gat));
  NAND4_X1  g563(.A1(new_n749), .A2(G43gat), .A3(new_n525), .A4(new_n753), .ZN(new_n765));
  OR2_X1    g564(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n595), .A2(new_n515), .A3(new_n756), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n767), .A2(new_n202), .B1(KEYINPUT107), .B2(KEYINPUT47), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n765), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n766), .B1(new_n765), .B2(new_n768), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n769), .A2(new_n770), .ZN(G1330gat));
  NAND2_X1  g570(.A1(new_n743), .A2(new_n741), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT87), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n537), .A2(new_n411), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n531), .B1(new_n472), .B2(new_n476), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n530), .B1(new_n483), .B2(new_n466), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT38), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n527), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n774), .A2(new_n777), .A3(new_n409), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n556), .A2(new_n549), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n537), .A2(new_n568), .A3(new_n571), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n352), .B1(new_n486), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n773), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n557), .A2(new_n577), .A3(KEYINPUT87), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n742), .B1(new_n786), .B2(new_n526), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n745), .B1(new_n772), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n747), .ZN(new_n789));
  INV_X1    g588(.A(new_n748), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n789), .A2(new_n558), .A3(new_n790), .A4(new_n753), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n234), .A2(new_n235), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT108), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n757), .A2(new_n352), .A3(new_n793), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n795), .B1(new_n791), .B2(new_n793), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT48), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n794), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  AOI221_X4 g597(.A(new_n795), .B1(KEYINPUT108), .B2(KEYINPUT48), .C1(new_n791), .C2(new_n793), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n798), .A2(new_n799), .ZN(G1331gat));
  AND4_X1   g599(.A1(new_n270), .A2(new_n687), .A3(new_n689), .A4(new_n752), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n744), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n415), .B(KEYINPUT109), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g605(.A1(new_n803), .A2(new_n485), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n807), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n808));
  XOR2_X1   g607(.A(KEYINPUT49), .B(G64gat), .Z(new_n809));
  OAI21_X1  g608(.A(new_n808), .B1(new_n807), .B2(new_n809), .ZN(G1333gat));
  OAI21_X1  g609(.A(G71gat), .B1(new_n802), .B2(new_n727), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n521), .A2(G71gat), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n811), .B1(new_n802), .B2(new_n812), .ZN(new_n813));
  XOR2_X1   g612(.A(new_n813), .B(KEYINPUT50), .Z(G1334gat));
  OR3_X1    g613(.A1(new_n802), .A2(KEYINPUT111), .A3(new_n352), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT111), .B1(new_n802), .B2(new_n352), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g616(.A(KEYINPUT110), .B(G78gat), .ZN(new_n818));
  XOR2_X1   g617(.A(new_n817), .B(new_n818), .Z(G1335gat));
  NOR2_X1   g618(.A1(new_n751), .A2(new_n269), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n712), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n749), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(G85gat), .B1(new_n823), .B2(new_n415), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n745), .B(new_n820), .C1(new_n772), .C2(new_n787), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT51), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n744), .A2(KEYINPUT51), .A3(new_n745), .A4(new_n820), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n829), .A2(new_n658), .A3(new_n585), .A4(new_n712), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n824), .A2(new_n830), .ZN(G1336gat));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n749), .A2(new_n485), .A3(new_n822), .ZN(new_n833));
  XOR2_X1   g632(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n834));
  NAND2_X1  g633(.A1(new_n825), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n828), .ZN(new_n836));
  INV_X1    g635(.A(new_n752), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n837), .A2(G92gat), .A3(new_n486), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n833), .A2(G92gat), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n833), .A2(G92gat), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n829), .A2(new_n838), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n832), .ZN(new_n842));
  OAI22_X1  g641(.A1(new_n832), .A2(new_n839), .B1(new_n840), .B2(new_n842), .ZN(G1337gat));
  OAI21_X1  g642(.A(G99gat), .B1(new_n823), .B2(new_n727), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n829), .A2(new_n664), .A3(new_n515), .A4(new_n712), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(G1338gat));
  NOR4_X1   g645(.A1(new_n746), .A2(new_n352), .A3(new_n748), .A4(new_n821), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n352), .A2(G106gat), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n752), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n849), .B1(new_n835), .B2(new_n828), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT113), .ZN(new_n851));
  OAI22_X1  g650(.A1(new_n847), .A2(new_n665), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT53), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n829), .A2(new_n752), .A3(new_n848), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n855), .B(new_n856), .C1(new_n665), .C2(new_n847), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n854), .A2(new_n857), .ZN(G1339gat));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n859), .B1(new_n708), .B2(new_n692), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n693), .B(new_n707), .C1(new_n691), .C2(KEYINPUT10), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n697), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n706), .A2(new_n859), .A3(new_n710), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n863), .A3(KEYINPUT55), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n705), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT55), .B1(new_n862), .B2(new_n863), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n248), .A2(new_n249), .A3(new_n247), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n245), .B1(new_n242), .B2(new_n244), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n256), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n263), .A2(new_n869), .ZN(new_n870));
  NOR4_X1   g669(.A1(new_n865), .A2(new_n866), .A3(new_n685), .A4(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n712), .A2(new_n263), .A3(new_n869), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n864), .A2(new_n269), .A3(new_n705), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(new_n874), .B2(new_n866), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n685), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n750), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n687), .A2(new_n270), .A3(new_n689), .A4(new_n713), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n880), .A2(new_n804), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n881), .A2(new_n592), .ZN(new_n882));
  AOI21_X1  g681(.A(G113gat), .B1(new_n882), .B2(new_n269), .ZN(new_n883));
  INV_X1    g682(.A(new_n879), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n884), .B1(new_n750), .B2(new_n877), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n558), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n415), .A2(new_n485), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n515), .A3(new_n887), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n888), .A2(new_n365), .A3(new_n270), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n883), .A2(new_n889), .ZN(G1340gat));
  OAI21_X1  g689(.A(G120gat), .B1(new_n888), .B2(new_n837), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n713), .A2(new_n367), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n882), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT114), .ZN(G1341gat));
  OAI21_X1  g694(.A(G127gat), .B1(new_n888), .B2(new_n750), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n882), .A2(new_n360), .A3(new_n751), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  XOR2_X1   g697(.A(new_n898), .B(KEYINPUT115), .Z(G1342gat));
  NAND3_X1  g698(.A1(new_n882), .A2(new_n358), .A3(new_n745), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n900), .A2(KEYINPUT56), .ZN(new_n901));
  OAI21_X1  g700(.A(G134gat), .B1(new_n888), .B2(new_n685), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(KEYINPUT56), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(G1343gat));
  NAND2_X1  g703(.A1(new_n727), .A2(new_n887), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n880), .A2(new_n558), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT57), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n352), .A2(new_n908), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  AND3_X1   g710(.A1(new_n864), .A2(new_n269), .A3(new_n705), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT55), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n706), .A2(new_n859), .A3(new_n710), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n704), .A2(KEYINPUT54), .A3(new_n861), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n698), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n913), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(KEYINPUT116), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT116), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n866), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n912), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n745), .B1(new_n921), .B2(new_n873), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n872), .B1(new_n922), .B2(KEYINPUT117), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT117), .ZN(new_n924));
  AOI211_X1 g723(.A(new_n924), .B(new_n745), .C1(new_n921), .C2(new_n873), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n750), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n911), .B1(new_n926), .B2(new_n879), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n909), .B1(new_n927), .B2(KEYINPUT118), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT118), .ZN(new_n929));
  AOI211_X1 g728(.A(new_n929), .B(new_n911), .C1(new_n926), .C2(new_n879), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n269), .B(new_n906), .C1(new_n928), .C2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT121), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n862), .A2(new_n863), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n919), .B1(new_n933), .B2(new_n913), .ZN(new_n934));
  AOI211_X1 g733(.A(KEYINPUT116), .B(KEYINPUT55), .C1(new_n862), .C2(new_n863), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n874), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(new_n873), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n685), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n871), .B1(new_n938), .B2(new_n924), .ZN(new_n939));
  INV_X1    g738(.A(new_n925), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n751), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n910), .B1(new_n941), .B2(new_n884), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(new_n929), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n927), .A2(KEYINPUT118), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n943), .A2(new_n944), .A3(new_n909), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT121), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n945), .A2(new_n946), .A3(new_n269), .A4(new_n906), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n932), .A2(G141gat), .A3(new_n947), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n525), .A2(new_n352), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n881), .A2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT120), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n485), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n881), .A2(KEYINPUT120), .A3(new_n949), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n270), .A2(G141gat), .ZN(new_n955));
  AOI21_X1  g754(.A(KEYINPUT58), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n948), .A2(new_n956), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n931), .A2(G141gat), .ZN(new_n958));
  INV_X1    g757(.A(new_n950), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n270), .A2(new_n485), .A3(G141gat), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT119), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n959), .A2(KEYINPUT119), .A3(new_n960), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(KEYINPUT58), .B1(new_n958), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n957), .A2(new_n966), .ZN(G1344gat));
  NAND3_X1  g766(.A1(new_n954), .A2(new_n291), .A3(new_n712), .ZN(new_n968));
  AOI22_X1  g767(.A1(new_n942), .A2(new_n929), .B1(new_n908), .B2(new_n907), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n905), .B1(new_n969), .B2(new_n944), .ZN(new_n970));
  AOI211_X1 g769(.A(KEYINPUT59), .B(new_n291), .C1(new_n970), .C2(new_n712), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT59), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n885), .A2(new_n908), .A3(new_n352), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n750), .B1(new_n922), .B2(new_n871), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(new_n879), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT57), .B1(new_n975), .B2(new_n558), .ZN(new_n976));
  OAI211_X1 g775(.A(new_n712), .B(new_n906), .C1(new_n973), .C2(new_n976), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n972), .B1(new_n977), .B2(G148gat), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n968), .B1(new_n971), .B2(new_n978), .ZN(G1345gat));
  NAND3_X1  g778(.A1(new_n954), .A2(new_n628), .A3(new_n751), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n970), .A2(new_n751), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n980), .B1(new_n981), .B2(new_n628), .ZN(G1346gat));
  AOI21_X1  g781(.A(G162gat), .B1(new_n954), .B2(new_n745), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n745), .A2(G162gat), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n983), .B1(new_n970), .B2(new_n984), .ZN(G1347gat));
  NOR2_X1   g784(.A1(new_n885), .A2(new_n585), .ZN(new_n986));
  AND4_X1   g785(.A1(new_n352), .A2(new_n986), .A3(new_n485), .A4(new_n515), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n987), .A2(new_n422), .A3(new_n269), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n988), .B(KEYINPUT122), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n804), .A2(new_n486), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(new_n515), .ZN(new_n991));
  XNOR2_X1  g790(.A(new_n991), .B(KEYINPUT123), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n992), .A2(new_n886), .ZN(new_n993));
  OAI21_X1  g792(.A(G169gat), .B1(new_n993), .B2(new_n270), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n989), .A2(new_n994), .ZN(G1348gat));
  NAND4_X1  g794(.A1(new_n992), .A2(G176gat), .A3(new_n752), .A4(new_n886), .ZN(new_n996));
  AND2_X1   g795(.A1(new_n996), .A2(KEYINPUT124), .ZN(new_n997));
  AOI21_X1  g796(.A(G176gat), .B1(new_n987), .B2(new_n712), .ZN(new_n998));
  NOR2_X1   g797(.A1(new_n996), .A2(KEYINPUT124), .ZN(new_n999));
  NOR3_X1   g798(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(G1349gat));
  OAI21_X1  g799(.A(KEYINPUT125), .B1(new_n993), .B2(new_n750), .ZN(new_n1001));
  INV_X1    g800(.A(KEYINPUT125), .ZN(new_n1002));
  NAND4_X1  g801(.A1(new_n992), .A2(new_n1002), .A3(new_n751), .A4(new_n886), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n1001), .A2(G183gat), .A3(new_n1003), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n987), .A2(new_n452), .A3(new_n751), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1006), .A2(KEYINPUT60), .ZN(new_n1007));
  INV_X1    g806(.A(KEYINPUT60), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n1004), .A2(new_n1008), .A3(new_n1005), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1007), .A2(new_n1009), .ZN(G1350gat));
  NAND3_X1  g809(.A1(new_n987), .A2(new_n433), .A3(new_n745), .ZN(new_n1011));
  OAI21_X1  g810(.A(G190gat), .B1(new_n993), .B2(new_n685), .ZN(new_n1012));
  AND2_X1   g811(.A1(new_n1012), .A2(KEYINPUT61), .ZN(new_n1013));
  NOR2_X1   g812(.A1(new_n1012), .A2(KEYINPUT61), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n1011), .B1(new_n1013), .B2(new_n1014), .ZN(G1351gat));
  AND3_X1   g814(.A1(new_n986), .A2(new_n485), .A3(new_n949), .ZN(new_n1016));
  AOI21_X1  g815(.A(G197gat), .B1(new_n1016), .B2(new_n269), .ZN(new_n1017));
  NOR2_X1   g816(.A1(new_n973), .A2(new_n976), .ZN(new_n1018));
  XNOR2_X1  g817(.A(new_n1018), .B(KEYINPUT126), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n990), .A2(new_n727), .ZN(new_n1020));
  INV_X1    g819(.A(new_n1020), .ZN(new_n1021));
  AND3_X1   g820(.A1(new_n1021), .A2(G197gat), .A3(new_n269), .ZN(new_n1022));
  AOI21_X1  g821(.A(new_n1017), .B1(new_n1019), .B2(new_n1022), .ZN(G1352gat));
  NAND2_X1  g822(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1024));
  OAI21_X1  g823(.A(G204gat), .B1(new_n1024), .B2(new_n837), .ZN(new_n1025));
  INV_X1    g824(.A(G204gat), .ZN(new_n1026));
  NAND3_X1  g825(.A1(new_n1016), .A2(new_n1026), .A3(new_n712), .ZN(new_n1027));
  XOR2_X1   g826(.A(new_n1027), .B(KEYINPUT62), .Z(new_n1028));
  NAND2_X1  g827(.A1(new_n1025), .A2(new_n1028), .ZN(G1353gat));
  NAND3_X1  g828(.A1(new_n1016), .A2(new_n304), .A3(new_n751), .ZN(new_n1030));
  OAI211_X1 g829(.A(new_n751), .B(new_n1021), .C1(new_n973), .C2(new_n976), .ZN(new_n1031));
  OR2_X1    g830(.A1(new_n1031), .A2(KEYINPUT127), .ZN(new_n1032));
  AOI21_X1  g831(.A(new_n304), .B1(new_n1031), .B2(KEYINPUT127), .ZN(new_n1033));
  AND3_X1   g832(.A1(new_n1032), .A2(KEYINPUT63), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g833(.A(KEYINPUT63), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1035));
  OAI21_X1  g834(.A(new_n1030), .B1(new_n1034), .B2(new_n1035), .ZN(G1354gat));
  AOI21_X1  g835(.A(G218gat), .B1(new_n1016), .B2(new_n745), .ZN(new_n1037));
  INV_X1    g836(.A(new_n1024), .ZN(new_n1038));
  NOR2_X1   g837(.A1(new_n685), .A2(new_n305), .ZN(new_n1039));
  AOI21_X1  g838(.A(new_n1037), .B1(new_n1038), .B2(new_n1039), .ZN(G1355gat));
endmodule


