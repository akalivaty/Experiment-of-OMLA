

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U553 ( .A(n652), .B(n651), .ZN(n658) );
  OR2_X1 U554 ( .A1(n756), .A2(n755), .ZN(n768) );
  AND2_X1 U555 ( .A1(n717), .A2(n520), .ZN(n756) );
  BUF_X1 U556 ( .A(n723), .Z(n724) );
  NOR2_X2 U557 ( .A1(G2105), .A2(G2104), .ZN(n526) );
  NOR2_X1 U558 ( .A1(n673), .A2(n980), .ZN(n602) );
  NAND2_X1 U559 ( .A1(n732), .A2(n733), .ZN(n673) );
  NAND2_X1 U560 ( .A1(G8), .A2(n673), .ZN(n716) );
  XNOR2_X1 U561 ( .A(n606), .B(n605), .ZN(n641) );
  INV_X1 U562 ( .A(KEYINPUT96), .ZN(n605) );
  INV_X1 U563 ( .A(KEYINPUT102), .ZN(n688) );
  NOR2_X1 U564 ( .A1(n687), .A2(n686), .ZN(n689) );
  XNOR2_X1 U565 ( .A(KEYINPUT32), .B(KEYINPUT106), .ZN(n681) );
  NAND2_X1 U566 ( .A1(n518), .A2(G8), .ZN(n682) );
  XNOR2_X1 U567 ( .A(n712), .B(KEYINPUT107), .ZN(n717) );
  XOR2_X1 U568 ( .A(n680), .B(KEYINPUT105), .Z(n518) );
  XNOR2_X1 U569 ( .A(n682), .B(n681), .ZN(n705) );
  OR2_X1 U570 ( .A1(n783), .A2(n645), .ZN(n519) );
  OR2_X1 U571 ( .A1(n716), .A2(n715), .ZN(n520) );
  OR2_X1 U572 ( .A1(n716), .A2(n702), .ZN(n521) );
  INV_X1 U573 ( .A(n989), .ZN(n783) );
  NOR2_X2 U574 ( .A1(n540), .A2(n539), .ZN(G160) );
  AND2_X1 U575 ( .A1(n753), .A2(n752), .ZN(n522) );
  AND2_X1 U576 ( .A1(n521), .A2(n913), .ZN(n523) );
  INV_X1 U577 ( .A(KEYINPUT99), .ZN(n659) );
  NOR2_X1 U578 ( .A1(n641), .A2(n642), .ZN(n608) );
  XNOR2_X1 U579 ( .A(n662), .B(KEYINPUT30), .ZN(n663) );
  XNOR2_X1 U580 ( .A(n689), .B(n688), .ZN(n706) );
  XNOR2_X1 U581 ( .A(n610), .B(KEYINPUT70), .ZN(n611) );
  XNOR2_X1 U582 ( .A(n612), .B(n611), .ZN(n614) );
  INV_X1 U583 ( .A(KEYINPUT17), .ZN(n525) );
  NAND2_X1 U584 ( .A1(n754), .A2(n522), .ZN(n755) );
  NOR2_X1 U585 ( .A1(n626), .A2(n625), .ZN(n628) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n578) );
  XOR2_X1 U587 ( .A(n628), .B(n627), .Z(n989) );
  NOR2_X2 U588 ( .A1(G651), .A2(G543), .ZN(n809) );
  NAND2_X1 U589 ( .A1(n1003), .A2(G137), .ZN(n538) );
  NOR2_X1 U590 ( .A1(n559), .A2(n558), .ZN(G171) );
  INV_X1 U591 ( .A(G2104), .ZN(n529) );
  NOR2_X2 U592 ( .A1(G2105), .A2(n529), .ZN(n723) );
  NAND2_X1 U593 ( .A1(n723), .A2(G102), .ZN(n524) );
  XNOR2_X1 U594 ( .A(n524), .B(KEYINPUT86), .ZN(n528) );
  XNOR2_X2 U595 ( .A(n526), .B(n525), .ZN(n1003) );
  NAND2_X1 U596 ( .A1(G138), .A2(n1003), .ZN(n527) );
  NAND2_X1 U597 ( .A1(n528), .A2(n527), .ZN(n533) );
  AND2_X1 U598 ( .A1(n529), .A2(G2105), .ZN(n999) );
  NAND2_X1 U599 ( .A1(G126), .A2(n999), .ZN(n531) );
  AND2_X1 U600 ( .A1(G2105), .A2(G2104), .ZN(n1000) );
  NAND2_X1 U601 ( .A1(G114), .A2(n1000), .ZN(n530) );
  NAND2_X1 U602 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U603 ( .A1(n533), .A2(n532), .ZN(G164) );
  NAND2_X1 U604 ( .A1(n1000), .A2(G113), .ZN(n536) );
  NAND2_X1 U605 ( .A1(G101), .A2(n723), .ZN(n534) );
  XOR2_X1 U606 ( .A(KEYINPUT23), .B(n534), .Z(n535) );
  NAND2_X1 U607 ( .A1(n536), .A2(n535), .ZN(n540) );
  NAND2_X1 U608 ( .A1(G125), .A2(n999), .ZN(n537) );
  NAND2_X1 U609 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X2 U610 ( .A1(G651), .A2(n578), .ZN(n805) );
  NAND2_X1 U611 ( .A1(G53), .A2(n805), .ZN(n544) );
  INV_X1 U612 ( .A(G651), .ZN(n546) );
  NOR2_X1 U613 ( .A1(G543), .A2(n546), .ZN(n542) );
  XNOR2_X1 U614 ( .A(KEYINPUT65), .B(KEYINPUT1), .ZN(n541) );
  XNOR2_X2 U615 ( .A(n542), .B(n541), .ZN(n806) );
  NAND2_X1 U616 ( .A1(G65), .A2(n806), .ZN(n543) );
  NAND2_X1 U617 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U618 ( .A(KEYINPUT68), .B(n545), .ZN(n549) );
  NOR2_X2 U619 ( .A1(n578), .A2(n546), .ZN(n813) );
  NAND2_X1 U620 ( .A1(G78), .A2(n813), .ZN(n547) );
  XNOR2_X1 U621 ( .A(KEYINPUT67), .B(n547), .ZN(n548) );
  NOR2_X1 U622 ( .A1(n549), .A2(n548), .ZN(n551) );
  NAND2_X1 U623 ( .A1(n809), .A2(G91), .ZN(n550) );
  NAND2_X1 U624 ( .A1(n551), .A2(n550), .ZN(G299) );
  NAND2_X1 U625 ( .A1(G52), .A2(n805), .ZN(n553) );
  NAND2_X1 U626 ( .A1(G64), .A2(n806), .ZN(n552) );
  NAND2_X1 U627 ( .A1(n553), .A2(n552), .ZN(n559) );
  NAND2_X1 U628 ( .A1(n813), .A2(G77), .ZN(n554) );
  XNOR2_X1 U629 ( .A(n554), .B(KEYINPUT66), .ZN(n556) );
  NAND2_X1 U630 ( .A1(G90), .A2(n809), .ZN(n555) );
  NAND2_X1 U631 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U632 ( .A(KEYINPUT9), .B(n557), .Z(n558) );
  NAND2_X1 U633 ( .A1(n809), .A2(G89), .ZN(n560) );
  XNOR2_X1 U634 ( .A(n560), .B(KEYINPUT4), .ZN(n562) );
  NAND2_X1 U635 ( .A1(G76), .A2(n813), .ZN(n561) );
  NAND2_X1 U636 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U637 ( .A(n563), .B(KEYINPUT5), .ZN(n568) );
  NAND2_X1 U638 ( .A1(G51), .A2(n805), .ZN(n565) );
  NAND2_X1 U639 ( .A1(G63), .A2(n806), .ZN(n564) );
  NAND2_X1 U640 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U641 ( .A(KEYINPUT6), .B(n566), .Z(n567) );
  NAND2_X1 U642 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U643 ( .A(n569), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U644 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U645 ( .A1(G75), .A2(n813), .ZN(n570) );
  XNOR2_X1 U646 ( .A(n570), .B(KEYINPUT83), .ZN(n577) );
  NAND2_X1 U647 ( .A1(G50), .A2(n805), .ZN(n572) );
  NAND2_X1 U648 ( .A1(G62), .A2(n806), .ZN(n571) );
  NAND2_X1 U649 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U650 ( .A(KEYINPUT82), .B(n573), .Z(n575) );
  NAND2_X1 U651 ( .A1(n809), .A2(G88), .ZN(n574) );
  NAND2_X1 U652 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U653 ( .A1(n577), .A2(n576), .ZN(G166) );
  INV_X1 U654 ( .A(G166), .ZN(G303) );
  NAND2_X1 U655 ( .A1(G651), .A2(G74), .ZN(n583) );
  NAND2_X1 U656 ( .A1(G49), .A2(n805), .ZN(n580) );
  NAND2_X1 U657 ( .A1(G87), .A2(n578), .ZN(n579) );
  NAND2_X1 U658 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U659 ( .A1(n806), .A2(n581), .ZN(n582) );
  NAND2_X1 U660 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U661 ( .A(KEYINPUT79), .B(n584), .Z(G288) );
  NAND2_X1 U662 ( .A1(G73), .A2(n813), .ZN(n585) );
  XOR2_X1 U663 ( .A(KEYINPUT2), .B(n585), .Z(n591) );
  NAND2_X1 U664 ( .A1(n809), .A2(G86), .ZN(n586) );
  XNOR2_X1 U665 ( .A(n586), .B(KEYINPUT80), .ZN(n588) );
  NAND2_X1 U666 ( .A1(G61), .A2(n806), .ZN(n587) );
  NAND2_X1 U667 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U668 ( .A(KEYINPUT81), .B(n589), .Z(n590) );
  NOR2_X1 U669 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U670 ( .A1(n805), .A2(G48), .ZN(n592) );
  NAND2_X1 U671 ( .A1(n593), .A2(n592), .ZN(G305) );
  NAND2_X1 U672 ( .A1(G47), .A2(n805), .ZN(n595) );
  NAND2_X1 U673 ( .A1(G60), .A2(n806), .ZN(n594) );
  NAND2_X1 U674 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U675 ( .A1(G85), .A2(n809), .ZN(n597) );
  NAND2_X1 U676 ( .A1(G72), .A2(n813), .ZN(n596) );
  NAND2_X1 U677 ( .A1(n597), .A2(n596), .ZN(n598) );
  OR2_X1 U678 ( .A1(n599), .A2(n598), .ZN(G290) );
  NOR2_X1 U679 ( .A1(G164), .A2(G1384), .ZN(n732) );
  NAND2_X1 U680 ( .A1(G160), .A2(G40), .ZN(n600) );
  XNOR2_X1 U681 ( .A(n600), .B(KEYINPUT87), .ZN(n733) );
  INV_X1 U682 ( .A(G2072), .ZN(n980) );
  XOR2_X1 U683 ( .A(KEYINPUT27), .B(KEYINPUT95), .Z(n601) );
  XNOR2_X1 U684 ( .A(n602), .B(n601), .ZN(n604) );
  NAND2_X1 U685 ( .A1(n673), .A2(G1956), .ZN(n603) );
  NAND2_X1 U686 ( .A1(n604), .A2(n603), .ZN(n606) );
  INV_X1 U687 ( .A(G299), .ZN(n642) );
  XNOR2_X1 U688 ( .A(KEYINPUT97), .B(KEYINPUT28), .ZN(n607) );
  XNOR2_X1 U689 ( .A(n608), .B(n607), .ZN(n650) );
  NAND2_X1 U690 ( .A1(G43), .A2(n805), .ZN(n619) );
  NAND2_X1 U691 ( .A1(G56), .A2(n806), .ZN(n609) );
  XOR2_X1 U692 ( .A(KEYINPUT14), .B(n609), .Z(n617) );
  NAND2_X1 U693 ( .A1(G81), .A2(n809), .ZN(n612) );
  XOR2_X1 U694 ( .A(KEYINPUT12), .B(KEYINPUT71), .Z(n610) );
  NAND2_X1 U695 ( .A1(n813), .A2(G68), .ZN(n613) );
  NAND2_X1 U696 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U697 ( .A(KEYINPUT13), .B(n615), .Z(n616) );
  NOR2_X1 U698 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U699 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U700 ( .A(n620), .B(KEYINPUT72), .ZN(n987) );
  INV_X1 U701 ( .A(n673), .ZN(n654) );
  NAND2_X1 U702 ( .A1(G54), .A2(n805), .ZN(n622) );
  NAND2_X1 U703 ( .A1(G66), .A2(n806), .ZN(n621) );
  NAND2_X1 U704 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U705 ( .A1(G92), .A2(n809), .ZN(n624) );
  NAND2_X1 U706 ( .A1(G79), .A2(n813), .ZN(n623) );
  NAND2_X1 U707 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U708 ( .A(KEYINPUT74), .B(KEYINPUT15), .ZN(n627) );
  INV_X1 U709 ( .A(G1348), .ZN(n629) );
  OR2_X1 U710 ( .A1(n989), .A2(n629), .ZN(n630) );
  NAND2_X1 U711 ( .A1(KEYINPUT26), .A2(n630), .ZN(n631) );
  NOR2_X1 U712 ( .A1(n631), .A2(G1341), .ZN(n632) );
  NOR2_X1 U713 ( .A1(n654), .A2(n632), .ZN(n633) );
  NOR2_X1 U714 ( .A1(n987), .A2(n633), .ZN(n638) );
  NAND2_X1 U715 ( .A1(KEYINPUT26), .A2(G1996), .ZN(n635) );
  NAND2_X1 U716 ( .A1(n783), .A2(G2067), .ZN(n634) );
  NAND2_X1 U717 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U718 ( .A1(n654), .A2(n636), .ZN(n637) );
  NAND2_X1 U719 ( .A1(n638), .A2(n637), .ZN(n640) );
  NOR2_X1 U720 ( .A1(G1996), .A2(KEYINPUT26), .ZN(n639) );
  NOR2_X1 U721 ( .A1(n640), .A2(n639), .ZN(n648) );
  NAND2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U723 ( .A1(G1348), .A2(n673), .ZN(n644) );
  NAND2_X1 U724 ( .A1(G2067), .A2(n654), .ZN(n643) );
  NAND2_X1 U725 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U726 ( .A1(n646), .A2(n519), .ZN(n647) );
  OR2_X1 U727 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U728 ( .A1(n650), .A2(n649), .ZN(n652) );
  XOR2_X1 U729 ( .A(KEYINPUT29), .B(KEYINPUT98), .Z(n651) );
  XNOR2_X1 U730 ( .A(G2078), .B(KEYINPUT25), .ZN(n653) );
  XNOR2_X1 U731 ( .A(n653), .B(KEYINPUT94), .ZN(n893) );
  NOR2_X1 U732 ( .A1(n893), .A2(n673), .ZN(n656) );
  INV_X1 U733 ( .A(G1961), .ZN(n972) );
  NOR2_X1 U734 ( .A1(n654), .A2(n972), .ZN(n655) );
  NOR2_X1 U735 ( .A1(n656), .A2(n655), .ZN(n664) );
  NAND2_X1 U736 ( .A1(G171), .A2(n664), .ZN(n657) );
  NAND2_X1 U737 ( .A1(n658), .A2(n657), .ZN(n671) );
  NOR2_X1 U738 ( .A1(G1966), .A2(n716), .ZN(n686) );
  NOR2_X1 U739 ( .A1(G2084), .A2(n673), .ZN(n683) );
  NOR2_X1 U740 ( .A1(n686), .A2(n683), .ZN(n660) );
  XNOR2_X1 U741 ( .A(n660), .B(n659), .ZN(n661) );
  NAND2_X1 U742 ( .A1(n661), .A2(G8), .ZN(n662) );
  NOR2_X1 U743 ( .A1(G168), .A2(n663), .ZN(n667) );
  NOR2_X1 U744 ( .A1(G171), .A2(n664), .ZN(n665) );
  XNOR2_X1 U745 ( .A(n665), .B(KEYINPUT100), .ZN(n666) );
  NOR2_X1 U746 ( .A1(n667), .A2(n666), .ZN(n669) );
  XNOR2_X1 U747 ( .A(KEYINPUT31), .B(KEYINPUT101), .ZN(n668) );
  XNOR2_X1 U748 ( .A(n669), .B(n668), .ZN(n670) );
  NAND2_X1 U749 ( .A1(n671), .A2(n670), .ZN(n685) );
  NAND2_X1 U750 ( .A1(n685), .A2(G286), .ZN(n679) );
  NOR2_X1 U751 ( .A1(G1971), .A2(n716), .ZN(n672) );
  XOR2_X1 U752 ( .A(KEYINPUT103), .B(n672), .Z(n676) );
  NOR2_X1 U753 ( .A1(G2090), .A2(n673), .ZN(n674) );
  XNOR2_X1 U754 ( .A(KEYINPUT104), .B(n674), .ZN(n675) );
  NOR2_X1 U755 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U756 ( .A1(n677), .A2(G303), .ZN(n678) );
  NAND2_X1 U757 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U758 ( .A1(G8), .A2(n683), .ZN(n684) );
  NAND2_X1 U759 ( .A1(n685), .A2(n684), .ZN(n687) );
  NAND2_X1 U760 ( .A1(G1976), .A2(G288), .ZN(n922) );
  AND2_X1 U761 ( .A1(n706), .A2(n922), .ZN(n690) );
  NAND2_X1 U762 ( .A1(n705), .A2(n690), .ZN(n696) );
  INV_X1 U763 ( .A(n716), .ZN(n694) );
  INV_X1 U764 ( .A(n922), .ZN(n692) );
  NOR2_X1 U765 ( .A1(G1976), .A2(G288), .ZN(n701) );
  NOR2_X1 U766 ( .A1(G1971), .A2(G303), .ZN(n691) );
  NOR2_X1 U767 ( .A1(n701), .A2(n691), .ZN(n919) );
  NOR2_X1 U768 ( .A1(n692), .A2(n919), .ZN(n693) );
  NAND2_X1 U769 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U770 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U771 ( .A(n697), .B(KEYINPUT64), .ZN(n698) );
  INV_X1 U772 ( .A(n698), .ZN(n700) );
  INV_X1 U773 ( .A(KEYINPUT33), .ZN(n699) );
  NAND2_X1 U774 ( .A1(n700), .A2(n699), .ZN(n703) );
  NAND2_X1 U775 ( .A1(n701), .A2(KEYINPUT33), .ZN(n702) );
  XOR2_X1 U776 ( .A(G1981), .B(G305), .Z(n913) );
  NAND2_X1 U777 ( .A1(n703), .A2(n523), .ZN(n711) );
  NOR2_X1 U778 ( .A1(G2090), .A2(G303), .ZN(n704) );
  NAND2_X1 U779 ( .A1(G8), .A2(n704), .ZN(n708) );
  NAND2_X1 U780 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U781 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U782 ( .A1(n709), .A2(n716), .ZN(n710) );
  NAND2_X1 U783 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U784 ( .A1(G1981), .A2(G305), .ZN(n713) );
  XNOR2_X1 U785 ( .A(KEYINPUT93), .B(n713), .ZN(n714) );
  XNOR2_X1 U786 ( .A(KEYINPUT24), .B(n714), .ZN(n715) );
  XNOR2_X1 U787 ( .A(G2067), .B(KEYINPUT37), .ZN(n718) );
  XOR2_X1 U788 ( .A(n718), .B(KEYINPUT89), .Z(n763) );
  NAND2_X1 U789 ( .A1(n1000), .A2(G116), .ZN(n719) );
  XNOR2_X1 U790 ( .A(n719), .B(KEYINPUT90), .ZN(n721) );
  NAND2_X1 U791 ( .A1(G128), .A2(n999), .ZN(n720) );
  NAND2_X1 U792 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U793 ( .A(n722), .B(KEYINPUT35), .ZN(n729) );
  NAND2_X1 U794 ( .A1(G104), .A2(n724), .ZN(n726) );
  NAND2_X1 U795 ( .A1(G140), .A2(n1003), .ZN(n725) );
  NAND2_X1 U796 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U797 ( .A(KEYINPUT34), .B(n727), .Z(n728) );
  NAND2_X1 U798 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U799 ( .A(n730), .B(KEYINPUT36), .Z(n996) );
  OR2_X1 U800 ( .A1(n763), .A2(n996), .ZN(n731) );
  XOR2_X1 U801 ( .A(n731), .B(KEYINPUT91), .Z(n876) );
  INV_X1 U802 ( .A(n732), .ZN(n734) );
  NAND2_X1 U803 ( .A1(n734), .A2(n733), .ZN(n750) );
  OR2_X1 U804 ( .A1(n876), .A2(n750), .ZN(n754) );
  XNOR2_X1 U805 ( .A(G1986), .B(G290), .ZN(n921) );
  INV_X1 U806 ( .A(n750), .ZN(n765) );
  NAND2_X1 U807 ( .A1(n921), .A2(n765), .ZN(n735) );
  XNOR2_X1 U808 ( .A(n735), .B(KEYINPUT88), .ZN(n753) );
  NAND2_X1 U809 ( .A1(G105), .A2(n724), .ZN(n736) );
  XNOR2_X1 U810 ( .A(n736), .B(KEYINPUT38), .ZN(n743) );
  NAND2_X1 U811 ( .A1(G141), .A2(n1003), .ZN(n738) );
  NAND2_X1 U812 ( .A1(G117), .A2(n1000), .ZN(n737) );
  NAND2_X1 U813 ( .A1(n738), .A2(n737), .ZN(n741) );
  NAND2_X1 U814 ( .A1(n999), .A2(G129), .ZN(n739) );
  XOR2_X1 U815 ( .A(KEYINPUT92), .B(n739), .Z(n740) );
  NOR2_X1 U816 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U817 ( .A1(n743), .A2(n742), .ZN(n994) );
  AND2_X1 U818 ( .A1(n994), .A2(G1996), .ZN(n873) );
  NAND2_X1 U819 ( .A1(G95), .A2(n724), .ZN(n745) );
  NAND2_X1 U820 ( .A1(G131), .A2(n1003), .ZN(n744) );
  NAND2_X1 U821 ( .A1(n745), .A2(n744), .ZN(n749) );
  NAND2_X1 U822 ( .A1(G119), .A2(n999), .ZN(n747) );
  NAND2_X1 U823 ( .A1(G107), .A2(n1000), .ZN(n746) );
  NAND2_X1 U824 ( .A1(n747), .A2(n746), .ZN(n748) );
  OR2_X1 U825 ( .A1(n749), .A2(n748), .ZN(n1019) );
  AND2_X1 U826 ( .A1(n1019), .A2(G1991), .ZN(n868) );
  NOR2_X1 U827 ( .A1(n873), .A2(n868), .ZN(n751) );
  NOR2_X1 U828 ( .A1(n751), .A2(n750), .ZN(n759) );
  INV_X1 U829 ( .A(n759), .ZN(n752) );
  NOR2_X1 U830 ( .A1(G1996), .A2(n994), .ZN(n865) );
  NOR2_X1 U831 ( .A1(G1986), .A2(G290), .ZN(n757) );
  NOR2_X1 U832 ( .A1(G1991), .A2(n1019), .ZN(n867) );
  NOR2_X1 U833 ( .A1(n757), .A2(n867), .ZN(n758) );
  NOR2_X1 U834 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U835 ( .A1(n865), .A2(n760), .ZN(n761) );
  XNOR2_X1 U836 ( .A(n761), .B(KEYINPUT39), .ZN(n762) );
  NAND2_X1 U837 ( .A1(n762), .A2(n876), .ZN(n764) );
  NAND2_X1 U838 ( .A1(n996), .A2(n763), .ZN(n877) );
  NAND2_X1 U839 ( .A1(n764), .A2(n877), .ZN(n766) );
  NAND2_X1 U840 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U841 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U842 ( .A(n769), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U843 ( .A(G1341), .B(G2427), .ZN(n779) );
  XOR2_X1 U844 ( .A(G2451), .B(KEYINPUT109), .Z(n771) );
  XNOR2_X1 U845 ( .A(G1348), .B(G2443), .ZN(n770) );
  XNOR2_X1 U846 ( .A(n771), .B(n770), .ZN(n775) );
  XOR2_X1 U847 ( .A(G2438), .B(G2435), .Z(n773) );
  XNOR2_X1 U848 ( .A(G2430), .B(G2454), .ZN(n772) );
  XNOR2_X1 U849 ( .A(n773), .B(n772), .ZN(n774) );
  XOR2_X1 U850 ( .A(n775), .B(n774), .Z(n777) );
  XNOR2_X1 U851 ( .A(G2446), .B(KEYINPUT108), .ZN(n776) );
  XNOR2_X1 U852 ( .A(n777), .B(n776), .ZN(n778) );
  XNOR2_X1 U853 ( .A(n779), .B(n778), .ZN(n780) );
  AND2_X1 U854 ( .A1(n780), .A2(G14), .ZN(G401) );
  AND2_X1 U855 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U856 ( .A(G132), .ZN(G219) );
  INV_X1 U857 ( .A(G82), .ZN(G220) );
  NAND2_X1 U858 ( .A1(G7), .A2(G661), .ZN(n781) );
  XOR2_X1 U859 ( .A(n781), .B(KEYINPUT10), .Z(n1033) );
  NAND2_X1 U860 ( .A1(n1033), .A2(G567), .ZN(n782) );
  XOR2_X1 U861 ( .A(KEYINPUT11), .B(n782), .Z(G234) );
  INV_X1 U862 ( .A(G860), .ZN(n788) );
  OR2_X1 U863 ( .A1(n788), .A2(n987), .ZN(G153) );
  XNOR2_X1 U864 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U865 ( .A1(G868), .A2(G301), .ZN(n785) );
  INV_X1 U866 ( .A(G868), .ZN(n827) );
  NAND2_X1 U867 ( .A1(n783), .A2(n827), .ZN(n784) );
  NAND2_X1 U868 ( .A1(n785), .A2(n784), .ZN(G284) );
  NOR2_X1 U869 ( .A1(G868), .A2(G299), .ZN(n787) );
  NOR2_X1 U870 ( .A1(G286), .A2(n827), .ZN(n786) );
  NOR2_X1 U871 ( .A1(n787), .A2(n786), .ZN(G297) );
  NAND2_X1 U872 ( .A1(n788), .A2(G559), .ZN(n789) );
  NAND2_X1 U873 ( .A1(n789), .A2(n989), .ZN(n790) );
  XNOR2_X1 U874 ( .A(n790), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U875 ( .A1(n987), .A2(G868), .ZN(n793) );
  NAND2_X1 U876 ( .A1(n989), .A2(G868), .ZN(n791) );
  NOR2_X1 U877 ( .A1(G559), .A2(n791), .ZN(n792) );
  NOR2_X1 U878 ( .A1(n793), .A2(n792), .ZN(G282) );
  NAND2_X1 U879 ( .A1(G99), .A2(n724), .ZN(n795) );
  NAND2_X1 U880 ( .A1(G111), .A2(n1000), .ZN(n794) );
  NAND2_X1 U881 ( .A1(n795), .A2(n794), .ZN(n801) );
  NAND2_X1 U882 ( .A1(n999), .A2(G123), .ZN(n796) );
  XNOR2_X1 U883 ( .A(n796), .B(KEYINPUT18), .ZN(n798) );
  NAND2_X1 U884 ( .A1(G135), .A2(n1003), .ZN(n797) );
  NAND2_X1 U885 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U886 ( .A(KEYINPUT75), .B(n799), .Z(n800) );
  NOR2_X1 U887 ( .A1(n801), .A2(n800), .ZN(n995) );
  XNOR2_X1 U888 ( .A(n995), .B(G2096), .ZN(n802) );
  XNOR2_X1 U889 ( .A(n802), .B(KEYINPUT76), .ZN(n803) );
  INV_X1 U890 ( .A(G2100), .ZN(n977) );
  NAND2_X1 U891 ( .A1(n803), .A2(n977), .ZN(G156) );
  NAND2_X1 U892 ( .A1(n989), .A2(G559), .ZN(n804) );
  XNOR2_X1 U893 ( .A(n987), .B(n804), .ZN(n823) );
  NOR2_X1 U894 ( .A1(n823), .A2(G860), .ZN(n817) );
  NAND2_X1 U895 ( .A1(G55), .A2(n805), .ZN(n808) );
  NAND2_X1 U896 ( .A1(G67), .A2(n806), .ZN(n807) );
  NAND2_X1 U897 ( .A1(n808), .A2(n807), .ZN(n812) );
  NAND2_X1 U898 ( .A1(G93), .A2(n809), .ZN(n810) );
  XNOR2_X1 U899 ( .A(KEYINPUT77), .B(n810), .ZN(n811) );
  NOR2_X1 U900 ( .A1(n812), .A2(n811), .ZN(n815) );
  NAND2_X1 U901 ( .A1(n813), .A2(G80), .ZN(n814) );
  NAND2_X1 U902 ( .A1(n815), .A2(n814), .ZN(n826) );
  XOR2_X1 U903 ( .A(n826), .B(KEYINPUT78), .Z(n816) );
  XNOR2_X1 U904 ( .A(n817), .B(n816), .ZN(G145) );
  XOR2_X1 U905 ( .A(G299), .B(KEYINPUT19), .Z(n819) );
  XOR2_X1 U906 ( .A(G290), .B(G303), .Z(n818) );
  XNOR2_X1 U907 ( .A(n819), .B(n818), .ZN(n820) );
  XNOR2_X1 U908 ( .A(n820), .B(G288), .ZN(n821) );
  XNOR2_X1 U909 ( .A(n821), .B(n826), .ZN(n822) );
  XNOR2_X1 U910 ( .A(n822), .B(G305), .ZN(n988) );
  XOR2_X1 U911 ( .A(n988), .B(n823), .Z(n824) );
  NAND2_X1 U912 ( .A1(n824), .A2(G868), .ZN(n825) );
  XNOR2_X1 U913 ( .A(n825), .B(KEYINPUT84), .ZN(n829) );
  NAND2_X1 U914 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U915 ( .A1(n829), .A2(n828), .ZN(G295) );
  NAND2_X1 U916 ( .A1(G2078), .A2(G2084), .ZN(n830) );
  XOR2_X1 U917 ( .A(KEYINPUT20), .B(n830), .Z(n831) );
  NAND2_X1 U918 ( .A1(G2090), .A2(n831), .ZN(n833) );
  XOR2_X1 U919 ( .A(KEYINPUT21), .B(KEYINPUT85), .Z(n832) );
  XNOR2_X1 U920 ( .A(n833), .B(n832), .ZN(n834) );
  NAND2_X1 U921 ( .A1(G2072), .A2(n834), .ZN(G158) );
  XNOR2_X1 U922 ( .A(KEYINPUT69), .B(G57), .ZN(G237) );
  XNOR2_X1 U923 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U924 ( .A1(G108), .A2(G120), .ZN(n835) );
  NOR2_X1 U925 ( .A1(G237), .A2(n835), .ZN(n836) );
  NAND2_X1 U926 ( .A1(G69), .A2(n836), .ZN(n964) );
  NAND2_X1 U927 ( .A1(n964), .A2(G567), .ZN(n841) );
  NOR2_X1 U928 ( .A1(G220), .A2(G219), .ZN(n837) );
  XOR2_X1 U929 ( .A(KEYINPUT22), .B(n837), .Z(n838) );
  NOR2_X1 U930 ( .A1(G218), .A2(n838), .ZN(n839) );
  NAND2_X1 U931 ( .A1(G96), .A2(n839), .ZN(n965) );
  NAND2_X1 U932 ( .A1(n965), .A2(G2106), .ZN(n840) );
  NAND2_X1 U933 ( .A1(n841), .A2(n840), .ZN(n1032) );
  NAND2_X1 U934 ( .A1(G661), .A2(G483), .ZN(n842) );
  NOR2_X1 U935 ( .A1(n1032), .A2(n842), .ZN(n845) );
  NAND2_X1 U936 ( .A1(n845), .A2(G36), .ZN(G176) );
  NAND2_X1 U937 ( .A1(G2106), .A2(n1033), .ZN(G217) );
  AND2_X1 U938 ( .A1(G15), .A2(G2), .ZN(n843) );
  NAND2_X1 U939 ( .A1(G661), .A2(n843), .ZN(G259) );
  NAND2_X1 U940 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U941 ( .A1(n845), .A2(n844), .ZN(G188) );
  NAND2_X1 U943 ( .A1(G124), .A2(n999), .ZN(n846) );
  XOR2_X1 U944 ( .A(KEYINPUT111), .B(n846), .Z(n847) );
  XNOR2_X1 U945 ( .A(n847), .B(KEYINPUT44), .ZN(n849) );
  NAND2_X1 U946 ( .A1(G100), .A2(n724), .ZN(n848) );
  NAND2_X1 U947 ( .A1(n849), .A2(n848), .ZN(n853) );
  NAND2_X1 U948 ( .A1(G136), .A2(n1003), .ZN(n851) );
  NAND2_X1 U949 ( .A1(G112), .A2(n1000), .ZN(n850) );
  NAND2_X1 U950 ( .A1(n851), .A2(n850), .ZN(n852) );
  NOR2_X1 U951 ( .A1(n853), .A2(n852), .ZN(G162) );
  XOR2_X1 U952 ( .A(G164), .B(G2078), .Z(n862) );
  NAND2_X1 U953 ( .A1(G103), .A2(n724), .ZN(n855) );
  NAND2_X1 U954 ( .A1(G139), .A2(n1003), .ZN(n854) );
  NAND2_X1 U955 ( .A1(n855), .A2(n854), .ZN(n860) );
  NAND2_X1 U956 ( .A1(G127), .A2(n999), .ZN(n857) );
  NAND2_X1 U957 ( .A1(G115), .A2(n1000), .ZN(n856) );
  NAND2_X1 U958 ( .A1(n857), .A2(n856), .ZN(n858) );
  XOR2_X1 U959 ( .A(KEYINPUT47), .B(n858), .Z(n859) );
  NOR2_X1 U960 ( .A1(n860), .A2(n859), .ZN(n1018) );
  XOR2_X1 U961 ( .A(G2072), .B(n1018), .Z(n861) );
  NOR2_X1 U962 ( .A1(n862), .A2(n861), .ZN(n863) );
  XOR2_X1 U963 ( .A(KEYINPUT50), .B(n863), .Z(n882) );
  XOR2_X1 U964 ( .A(G2090), .B(G162), .Z(n864) );
  NOR2_X1 U965 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U966 ( .A(KEYINPUT51), .B(n866), .Z(n875) );
  NOR2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n871) );
  XOR2_X1 U968 ( .A(G2084), .B(G160), .Z(n869) );
  NOR2_X1 U969 ( .A1(n995), .A2(n869), .ZN(n870) );
  NAND2_X1 U970 ( .A1(n871), .A2(n870), .ZN(n872) );
  NOR2_X1 U971 ( .A1(n873), .A2(n872), .ZN(n874) );
  NAND2_X1 U972 ( .A1(n875), .A2(n874), .ZN(n879) );
  NAND2_X1 U973 ( .A1(n877), .A2(n876), .ZN(n878) );
  NOR2_X1 U974 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U975 ( .A(KEYINPUT119), .B(n880), .ZN(n881) );
  NOR2_X1 U976 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U977 ( .A(KEYINPUT52), .B(n883), .ZN(n885) );
  INV_X1 U978 ( .A(KEYINPUT55), .ZN(n884) );
  NAND2_X1 U979 ( .A1(n885), .A2(n884), .ZN(n886) );
  NAND2_X1 U980 ( .A1(n886), .A2(G29), .ZN(n962) );
  XNOR2_X1 U981 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n887) );
  XNOR2_X1 U982 ( .A(n887), .B(G34), .ZN(n888) );
  XNOR2_X1 U983 ( .A(G2084), .B(n888), .ZN(n904) );
  XNOR2_X1 U984 ( .A(G2090), .B(G35), .ZN(n902) );
  XOR2_X1 U985 ( .A(G1991), .B(G25), .Z(n889) );
  NAND2_X1 U986 ( .A1(n889), .A2(G28), .ZN(n890) );
  XNOR2_X1 U987 ( .A(n890), .B(KEYINPUT120), .ZN(n899) );
  XNOR2_X1 U988 ( .A(G1996), .B(G32), .ZN(n892) );
  XOR2_X1 U989 ( .A(G33), .B(n980), .Z(n891) );
  NOR2_X1 U990 ( .A1(n892), .A2(n891), .ZN(n897) );
  XOR2_X1 U991 ( .A(n893), .B(G27), .Z(n895) );
  XNOR2_X1 U992 ( .A(G26), .B(G2067), .ZN(n894) );
  NOR2_X1 U993 ( .A1(n895), .A2(n894), .ZN(n896) );
  NAND2_X1 U994 ( .A1(n897), .A2(n896), .ZN(n898) );
  NOR2_X1 U995 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U996 ( .A(KEYINPUT53), .B(n900), .ZN(n901) );
  NOR2_X1 U997 ( .A1(n902), .A2(n901), .ZN(n903) );
  NAND2_X1 U998 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U999 ( .A(KEYINPUT55), .B(n905), .Z(n907) );
  INV_X1 U1000 ( .A(G29), .ZN(n906) );
  NAND2_X1 U1001 ( .A1(n907), .A2(n906), .ZN(n908) );
  NAND2_X1 U1002 ( .A1(G11), .A2(n908), .ZN(n960) );
  INV_X1 U1003 ( .A(G16), .ZN(n956) );
  XOR2_X1 U1004 ( .A(n956), .B(KEYINPUT56), .Z(n929) );
  XOR2_X1 U1005 ( .A(G299), .B(G1956), .Z(n912) );
  XNOR2_X1 U1006 ( .A(G171), .B(n972), .ZN(n910) );
  XOR2_X1 U1007 ( .A(n989), .B(G1348), .Z(n909) );
  NOR2_X1 U1008 ( .A1(n910), .A2(n909), .ZN(n911) );
  NAND2_X1 U1009 ( .A1(n912), .A2(n911), .ZN(n917) );
  XNOR2_X1 U1010 ( .A(G168), .B(G1966), .ZN(n914) );
  NAND2_X1 U1011 ( .A1(n914), .A2(n913), .ZN(n915) );
  XOR2_X1 U1012 ( .A(KEYINPUT57), .B(n915), .Z(n916) );
  NOR2_X1 U1013 ( .A1(n917), .A2(n916), .ZN(n927) );
  NAND2_X1 U1014 ( .A1(G1971), .A2(G303), .ZN(n918) );
  NAND2_X1 U1015 ( .A1(n919), .A2(n918), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(n921), .A2(n920), .ZN(n923) );
  NAND2_X1 U1017 ( .A1(n923), .A2(n922), .ZN(n925) );
  XNOR2_X1 U1018 ( .A(G1341), .B(n987), .ZN(n924) );
  NOR2_X1 U1019 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1020 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1021 ( .A1(n929), .A2(n928), .ZN(n958) );
  XNOR2_X1 U1022 ( .A(G1986), .B(G24), .ZN(n934) );
  XNOR2_X1 U1023 ( .A(G1971), .B(G22), .ZN(n931) );
  XNOR2_X1 U1024 ( .A(G1976), .B(G23), .ZN(n930) );
  NOR2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1026 ( .A(KEYINPUT125), .B(n932), .ZN(n933) );
  NOR2_X1 U1027 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1028 ( .A(n935), .B(KEYINPUT58), .Z(n936) );
  XNOR2_X1 U1029 ( .A(KEYINPUT126), .B(n936), .ZN(n953) );
  XOR2_X1 U1030 ( .A(G1348), .B(KEYINPUT59), .Z(n937) );
  XNOR2_X1 U1031 ( .A(G4), .B(n937), .ZN(n945) );
  XOR2_X1 U1032 ( .A(G1341), .B(G19), .Z(n940) );
  XOR2_X1 U1033 ( .A(G20), .B(KEYINPUT122), .Z(n938) );
  XNOR2_X1 U1034 ( .A(n938), .B(G1956), .ZN(n939) );
  NAND2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n942) );
  XNOR2_X1 U1036 ( .A(G6), .B(G1981), .ZN(n941) );
  NOR2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(n943), .B(KEYINPUT123), .ZN(n944) );
  NOR2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(KEYINPUT60), .B(n946), .ZN(n948) );
  XOR2_X1 U1041 ( .A(G1961), .B(G5), .Z(n947) );
  NAND2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(G21), .B(G1966), .ZN(n949) );
  NOR2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1045 ( .A(KEYINPUT124), .B(n951), .Z(n952) );
  NOR2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(KEYINPUT61), .B(n954), .ZN(n955) );
  NAND2_X1 U1048 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1049 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1050 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1051 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1052 ( .A(KEYINPUT62), .B(n963), .Z(G311) );
  XNOR2_X1 U1053 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1054 ( .A(G120), .ZN(G236) );
  INV_X1 U1055 ( .A(G108), .ZN(G238) );
  INV_X1 U1056 ( .A(G96), .ZN(G221) );
  INV_X1 U1057 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(G325) );
  INV_X1 U1059 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U1060 ( .A(G1971), .B(G1976), .ZN(n976) );
  XOR2_X1 U1061 ( .A(G1966), .B(G1956), .Z(n967) );
  XNOR2_X1 U1062 ( .A(G1996), .B(G1981), .ZN(n966) );
  XNOR2_X1 U1063 ( .A(n967), .B(n966), .ZN(n971) );
  XOR2_X1 U1064 ( .A(KEYINPUT110), .B(KEYINPUT41), .Z(n969) );
  XNOR2_X1 U1065 ( .A(G1991), .B(G1986), .ZN(n968) );
  XNOR2_X1 U1066 ( .A(n969), .B(n968), .ZN(n970) );
  XOR2_X1 U1067 ( .A(n971), .B(n970), .Z(n974) );
  XOR2_X1 U1068 ( .A(n972), .B(G2474), .Z(n973) );
  XNOR2_X1 U1069 ( .A(n974), .B(n973), .ZN(n975) );
  XNOR2_X1 U1070 ( .A(n976), .B(n975), .ZN(G229) );
  XNOR2_X1 U1071 ( .A(n977), .B(G2096), .ZN(n979) );
  XNOR2_X1 U1072 ( .A(G2067), .B(G2090), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(n979), .B(n978), .ZN(n984) );
  XOR2_X1 U1074 ( .A(G2678), .B(KEYINPUT42), .Z(n982) );
  XOR2_X1 U1075 ( .A(n980), .B(KEYINPUT43), .Z(n981) );
  XNOR2_X1 U1076 ( .A(n982), .B(n981), .ZN(n983) );
  XOR2_X1 U1077 ( .A(n984), .B(n983), .Z(n986) );
  XNOR2_X1 U1078 ( .A(G2078), .B(G2084), .ZN(n985) );
  XNOR2_X1 U1079 ( .A(n986), .B(n985), .ZN(G227) );
  XOR2_X1 U1080 ( .A(n988), .B(n987), .Z(n991) );
  XOR2_X1 U1081 ( .A(G171), .B(n989), .Z(n990) );
  XNOR2_X1 U1082 ( .A(n991), .B(n990), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(n992), .B(G286), .ZN(n993) );
  NOR2_X1 U1084 ( .A1(G37), .A2(n993), .ZN(G397) );
  XNOR2_X1 U1085 ( .A(n995), .B(n994), .ZN(n998) );
  XOR2_X1 U1086 ( .A(G164), .B(n996), .Z(n997) );
  XNOR2_X1 U1087 ( .A(n998), .B(n997), .ZN(n1011) );
  NAND2_X1 U1088 ( .A1(G130), .A2(n999), .ZN(n1002) );
  NAND2_X1 U1089 ( .A1(G118), .A2(n1000), .ZN(n1001) );
  NAND2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1009) );
  NAND2_X1 U1091 ( .A1(G106), .A2(n724), .ZN(n1005) );
  NAND2_X1 U1092 ( .A1(G142), .A2(n1003), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1094 ( .A(KEYINPUT45), .B(n1006), .Z(n1007) );
  XNOR2_X1 U1095 ( .A(KEYINPUT112), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1097 ( .A(n1011), .B(n1010), .Z(n1013) );
  XNOR2_X1 U1098 ( .A(G160), .B(G162), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(n1013), .B(n1012), .ZN(n1017) );
  XOR2_X1 U1100 ( .A(KEYINPUT46), .B(KEYINPUT113), .Z(n1015) );
  XNOR2_X1 U1101 ( .A(KEYINPUT114), .B(KEYINPUT48), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(n1015), .B(n1014), .ZN(n1016) );
  XOR2_X1 U1103 ( .A(n1017), .B(n1016), .Z(n1021) );
  XOR2_X1 U1104 ( .A(n1019), .B(n1018), .Z(n1020) );
  XNOR2_X1 U1105 ( .A(n1021), .B(n1020), .ZN(n1022) );
  NOR2_X1 U1106 ( .A1(G37), .A2(n1022), .ZN(n1023) );
  XOR2_X1 U1107 ( .A(KEYINPUT115), .B(n1023), .Z(G395) );
  XNOR2_X1 U1108 ( .A(KEYINPUT117), .B(KEYINPUT49), .ZN(n1025) );
  NOR2_X1 U1109 ( .A1(G229), .A2(G227), .ZN(n1024) );
  XNOR2_X1 U1110 ( .A(n1025), .B(n1024), .ZN(n1029) );
  NOR2_X1 U1111 ( .A1(n1032), .A2(G401), .ZN(n1026) );
  XOR2_X1 U1112 ( .A(KEYINPUT116), .B(n1026), .Z(n1027) );
  NOR2_X1 U1113 ( .A1(G397), .A2(n1027), .ZN(n1028) );
  NAND2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NOR2_X1 U1115 ( .A1(n1030), .A2(G395), .ZN(n1031) );
  XOR2_X1 U1116 ( .A(n1031), .B(KEYINPUT118), .Z(G225) );
  INV_X1 U1117 ( .A(G225), .ZN(G308) );
  INV_X1 U1118 ( .A(n1032), .ZN(G319) );
  INV_X1 U1119 ( .A(n1033), .ZN(G223) );
endmodule

