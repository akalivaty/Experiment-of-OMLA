

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U554 ( .A(n723), .B(n722), .ZN(n725) );
  XNOR2_X2 U555 ( .A(n539), .B(KEYINPUT23), .ZN(n540) );
  XNOR2_X2 U556 ( .A(n538), .B(KEYINPUT64), .ZN(n563) );
  AND2_X2 U557 ( .A1(G2104), .A2(n541), .ZN(n538) );
  BUF_X1 U558 ( .A(n611), .Z(n550) );
  XNOR2_X1 U559 ( .A(n545), .B(n544), .ZN(n893) );
  XNOR2_X2 U560 ( .A(n754), .B(KEYINPUT105), .ZN(n766) );
  AND2_X2 U561 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X2 U562 ( .A(n742), .B(KEYINPUT99), .ZN(n765) );
  NOR2_X1 U563 ( .A1(G2105), .A2(G2104), .ZN(n545) );
  NOR2_X1 U564 ( .A1(G299), .A2(n730), .ZN(n727) );
  NOR2_X1 U565 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U566 ( .A1(n749), .A2(n748), .ZN(n751) );
  INV_X1 U567 ( .A(G2105), .ZN(n541) );
  INV_X1 U568 ( .A(KEYINPUT108), .ZN(n777) );
  OR2_X1 U569 ( .A1(n830), .A2(n829), .ZN(n831) );
  NOR2_X1 U570 ( .A1(n549), .A2(n548), .ZN(n699) );
  OR2_X1 U571 ( .A1(n826), .A2(n813), .ZN(n522) );
  NAND2_X1 U572 ( .A1(n966), .A2(G2067), .ZN(n708) );
  INV_X1 U573 ( .A(KEYINPUT27), .ZN(n722) );
  INV_X1 U574 ( .A(KEYINPUT102), .ZN(n726) );
  NOR2_X1 U575 ( .A1(n764), .A2(n743), .ZN(n745) );
  INV_X1 U576 ( .A(KEYINPUT31), .ZN(n750) );
  INV_X1 U577 ( .A(KEYINPUT107), .ZN(n772) );
  NAND2_X1 U578 ( .A1(n780), .A2(n700), .ZN(n720) );
  NAND2_X1 U579 ( .A1(G8), .A2(n720), .ZN(n826) );
  NAND2_X1 U580 ( .A1(n664), .A2(G66), .ZN(n610) );
  INV_X1 U581 ( .A(KEYINPUT1), .ZN(n523) );
  INV_X1 U582 ( .A(KEYINPUT17), .ZN(n544) );
  AND2_X1 U583 ( .A1(n814), .A2(n522), .ZN(n815) );
  XNOR2_X1 U584 ( .A(KEYINPUT15), .B(KEYINPUT72), .ZN(n617) );
  BUF_X1 U585 ( .A(n699), .Z(G160) );
  INV_X1 U586 ( .A(G651), .ZN(n533) );
  NOR2_X1 U587 ( .A1(G543), .A2(n533), .ZN(n524) );
  XNOR2_X2 U588 ( .A(n524), .B(n523), .ZN(n664) );
  NAND2_X1 U589 ( .A1(n664), .A2(G65), .ZN(n525) );
  XOR2_X1 U590 ( .A(KEYINPUT67), .B(n525), .Z(n531) );
  INV_X1 U591 ( .A(G543), .ZN(n526) );
  NAND2_X1 U592 ( .A1(KEYINPUT0), .A2(n526), .ZN(n529) );
  INV_X1 U593 ( .A(KEYINPUT0), .ZN(n527) );
  NAND2_X1 U594 ( .A1(n527), .A2(G543), .ZN(n528) );
  NAND2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n660) );
  NOR2_X1 U596 ( .A1(n660), .A2(G651), .ZN(n611) );
  NAND2_X1 U597 ( .A1(n611), .A2(G53), .ZN(n530) );
  NAND2_X1 U598 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U599 ( .A(KEYINPUT68), .B(n532), .Z(n537) );
  NOR2_X2 U600 ( .A1(G543), .A2(G651), .ZN(n656) );
  NAND2_X1 U601 ( .A1(G91), .A2(n656), .ZN(n535) );
  NOR2_X4 U602 ( .A1(n660), .A2(n533), .ZN(n652) );
  NAND2_X1 U603 ( .A1(G78), .A2(n652), .ZN(n534) );
  AND2_X1 U604 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U605 ( .A1(n537), .A2(n536), .ZN(G299) );
  NAND2_X1 U606 ( .A1(n563), .A2(G101), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(KEYINPUT65), .ZN(n543) );
  NOR2_X1 U608 ( .A1(G2104), .A2(n541), .ZN(n898) );
  NAND2_X1 U609 ( .A1(G125), .A2(n898), .ZN(n542) );
  NAND2_X1 U610 ( .A1(n543), .A2(n542), .ZN(n549) );
  NAND2_X1 U611 ( .A1(G137), .A2(n893), .ZN(n547) );
  AND2_X1 U612 ( .A1(G2105), .A2(G2104), .ZN(n899) );
  NAND2_X1 U613 ( .A1(G113), .A2(n899), .ZN(n546) );
  NAND2_X1 U614 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U615 ( .A(KEYINPUT74), .B(KEYINPUT6), .ZN(n554) );
  NAND2_X1 U616 ( .A1(G63), .A2(n664), .ZN(n552) );
  NAND2_X1 U617 ( .A1(G51), .A2(n550), .ZN(n551) );
  NAND2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(n561) );
  NAND2_X1 U620 ( .A1(n656), .A2(G89), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(KEYINPUT4), .ZN(n557) );
  NAND2_X1 U622 ( .A1(G76), .A2(n652), .ZN(n556) );
  NAND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(KEYINPUT73), .B(n558), .ZN(n559) );
  XNOR2_X1 U625 ( .A(KEYINPUT5), .B(n559), .ZN(n560) );
  NOR2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U627 ( .A(KEYINPUT7), .B(n562), .Z(G168) );
  XOR2_X1 U628 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U629 ( .A1(G138), .A2(n893), .ZN(n566) );
  INV_X1 U630 ( .A(n563), .ZN(n564) );
  INV_X1 U631 ( .A(n564), .ZN(n894) );
  NAND2_X1 U632 ( .A1(G102), .A2(n894), .ZN(n565) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n570) );
  NAND2_X1 U634 ( .A1(G126), .A2(n898), .ZN(n568) );
  NAND2_X1 U635 ( .A1(G114), .A2(n899), .ZN(n567) );
  NAND2_X1 U636 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U637 ( .A1(n570), .A2(n569), .ZN(G164) );
  NAND2_X1 U638 ( .A1(G60), .A2(n664), .ZN(n572) );
  NAND2_X1 U639 ( .A1(G47), .A2(n550), .ZN(n571) );
  NAND2_X1 U640 ( .A1(n572), .A2(n571), .ZN(n576) );
  NAND2_X1 U641 ( .A1(G85), .A2(n656), .ZN(n574) );
  NAND2_X1 U642 ( .A1(G72), .A2(n652), .ZN(n573) );
  NAND2_X1 U643 ( .A1(n574), .A2(n573), .ZN(n575) );
  OR2_X1 U644 ( .A1(n576), .A2(n575), .ZN(G290) );
  AND2_X1 U645 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U646 ( .A1(n898), .A2(G123), .ZN(n577) );
  XNOR2_X1 U647 ( .A(n577), .B(KEYINPUT18), .ZN(n579) );
  NAND2_X1 U648 ( .A1(G135), .A2(n893), .ZN(n578) );
  NAND2_X1 U649 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U650 ( .A(n580), .B(KEYINPUT77), .ZN(n582) );
  NAND2_X1 U651 ( .A1(G111), .A2(n899), .ZN(n581) );
  NAND2_X1 U652 ( .A1(n582), .A2(n581), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n894), .A2(G99), .ZN(n583) );
  XOR2_X1 U654 ( .A(KEYINPUT78), .B(n583), .Z(n584) );
  NOR2_X1 U655 ( .A1(n585), .A2(n584), .ZN(n1023) );
  XNOR2_X1 U656 ( .A(n1023), .B(G2096), .ZN(n586) );
  XNOR2_X1 U657 ( .A(n586), .B(KEYINPUT79), .ZN(n587) );
  OR2_X1 U658 ( .A1(G2100), .A2(n587), .ZN(G156) );
  INV_X1 U659 ( .A(G108), .ZN(G238) );
  INV_X1 U660 ( .A(G120), .ZN(G236) );
  INV_X1 U661 ( .A(G69), .ZN(G235) );
  INV_X1 U662 ( .A(G132), .ZN(G219) );
  INV_X1 U663 ( .A(G82), .ZN(G220) );
  NAND2_X1 U664 ( .A1(G64), .A2(n664), .ZN(n589) );
  NAND2_X1 U665 ( .A1(G52), .A2(n550), .ZN(n588) );
  NAND2_X1 U666 ( .A1(n589), .A2(n588), .ZN(n595) );
  NAND2_X1 U667 ( .A1(n656), .A2(G90), .ZN(n590) );
  XNOR2_X1 U668 ( .A(n590), .B(KEYINPUT66), .ZN(n592) );
  NAND2_X1 U669 ( .A1(G77), .A2(n652), .ZN(n591) );
  NAND2_X1 U670 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U671 ( .A(KEYINPUT9), .B(n593), .Z(n594) );
  NOR2_X1 U672 ( .A1(n595), .A2(n594), .ZN(G171) );
  NAND2_X1 U673 ( .A1(G7), .A2(G661), .ZN(n596) );
  XNOR2_X1 U674 ( .A(n596), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U675 ( .A(G223), .ZN(n849) );
  NAND2_X1 U676 ( .A1(n849), .A2(G567), .ZN(n597) );
  XOR2_X1 U677 ( .A(KEYINPUT11), .B(n597), .Z(G234) );
  NAND2_X1 U678 ( .A1(G56), .A2(n664), .ZN(n598) );
  XOR2_X1 U679 ( .A(KEYINPUT14), .B(n598), .Z(n599) );
  XNOR2_X1 U680 ( .A(n599), .B(KEYINPUT69), .ZN(n601) );
  NAND2_X1 U681 ( .A1(G43), .A2(n611), .ZN(n600) );
  NAND2_X1 U682 ( .A1(n601), .A2(n600), .ZN(n608) );
  NAND2_X1 U683 ( .A1(n656), .A2(G81), .ZN(n602) );
  XNOR2_X1 U684 ( .A(n602), .B(KEYINPUT12), .ZN(n604) );
  NAND2_X1 U685 ( .A1(G68), .A2(n652), .ZN(n603) );
  NAND2_X1 U686 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U687 ( .A(KEYINPUT13), .B(n605), .Z(n606) );
  XNOR2_X1 U688 ( .A(KEYINPUT70), .B(n606), .ZN(n607) );
  NOR2_X1 U689 ( .A1(n608), .A2(n607), .ZN(n964) );
  NAND2_X1 U690 ( .A1(n964), .A2(G860), .ZN(G153) );
  INV_X1 U691 ( .A(G171), .ZN(G301) );
  NAND2_X1 U692 ( .A1(G92), .A2(n656), .ZN(n609) );
  NAND2_X1 U693 ( .A1(n610), .A2(n609), .ZN(n616) );
  NAND2_X1 U694 ( .A1(G79), .A2(n652), .ZN(n613) );
  NAND2_X1 U695 ( .A1(G54), .A2(n611), .ZN(n612) );
  NAND2_X1 U696 ( .A1(n613), .A2(n612), .ZN(n614) );
  XOR2_X1 U697 ( .A(n614), .B(KEYINPUT71), .Z(n615) );
  NOR2_X1 U698 ( .A1(n616), .A2(n615), .ZN(n618) );
  XNOR2_X2 U699 ( .A(n618), .B(n617), .ZN(n966) );
  NOR2_X1 U700 ( .A1(n966), .A2(G868), .ZN(n620) );
  INV_X1 U701 ( .A(G868), .ZN(n627) );
  NOR2_X1 U702 ( .A1(n627), .A2(G301), .ZN(n619) );
  NOR2_X1 U703 ( .A1(n620), .A2(n619), .ZN(G284) );
  NOR2_X1 U704 ( .A1(G286), .A2(n627), .ZN(n622) );
  NOR2_X1 U705 ( .A1(G868), .A2(G299), .ZN(n621) );
  NOR2_X1 U706 ( .A1(n622), .A2(n621), .ZN(G297) );
  INV_X1 U707 ( .A(G559), .ZN(n623) );
  NOR2_X1 U708 ( .A1(G860), .A2(n623), .ZN(n624) );
  XNOR2_X1 U709 ( .A(KEYINPUT75), .B(n624), .ZN(n625) );
  INV_X1 U710 ( .A(n966), .ZN(n638) );
  NAND2_X1 U711 ( .A1(n625), .A2(n638), .ZN(n626) );
  XNOR2_X1 U712 ( .A(n626), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U713 ( .A1(n964), .A2(n627), .ZN(n628) );
  XOR2_X1 U714 ( .A(KEYINPUT76), .B(n628), .Z(n631) );
  NAND2_X1 U715 ( .A1(G868), .A2(n638), .ZN(n629) );
  NOR2_X1 U716 ( .A1(G559), .A2(n629), .ZN(n630) );
  NOR2_X1 U717 ( .A1(n631), .A2(n630), .ZN(G282) );
  NAND2_X1 U718 ( .A1(G67), .A2(n664), .ZN(n633) );
  NAND2_X1 U719 ( .A1(G55), .A2(n550), .ZN(n632) );
  NAND2_X1 U720 ( .A1(n633), .A2(n632), .ZN(n637) );
  NAND2_X1 U721 ( .A1(G93), .A2(n656), .ZN(n635) );
  NAND2_X1 U722 ( .A1(G80), .A2(n652), .ZN(n634) );
  NAND2_X1 U723 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U724 ( .A1(n637), .A2(n636), .ZN(n670) );
  NAND2_X1 U725 ( .A1(G559), .A2(n638), .ZN(n678) );
  XOR2_X1 U726 ( .A(n964), .B(n678), .Z(n639) );
  NOR2_X1 U727 ( .A1(G860), .A2(n639), .ZN(n640) );
  XNOR2_X1 U728 ( .A(n670), .B(n640), .ZN(G145) );
  NAND2_X1 U729 ( .A1(n550), .A2(G50), .ZN(n641) );
  XNOR2_X1 U730 ( .A(n641), .B(KEYINPUT82), .ZN(n643) );
  NAND2_X1 U731 ( .A1(G62), .A2(n664), .ZN(n642) );
  NAND2_X1 U732 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U733 ( .A(KEYINPUT83), .B(n644), .ZN(n649) );
  NAND2_X1 U734 ( .A1(G88), .A2(n656), .ZN(n646) );
  NAND2_X1 U735 ( .A1(G75), .A2(n652), .ZN(n645) );
  NAND2_X1 U736 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U737 ( .A(KEYINPUT84), .B(n647), .Z(n648) );
  NAND2_X1 U738 ( .A1(n649), .A2(n648), .ZN(G303) );
  INV_X1 U739 ( .A(G303), .ZN(G166) );
  NAND2_X1 U740 ( .A1(G61), .A2(n664), .ZN(n651) );
  NAND2_X1 U741 ( .A1(G48), .A2(n550), .ZN(n650) );
  NAND2_X1 U742 ( .A1(n651), .A2(n650), .ZN(n655) );
  NAND2_X1 U743 ( .A1(n652), .A2(G73), .ZN(n653) );
  XOR2_X1 U744 ( .A(KEYINPUT2), .B(n653), .Z(n654) );
  NOR2_X1 U745 ( .A1(n655), .A2(n654), .ZN(n658) );
  NAND2_X1 U746 ( .A1(n656), .A2(G86), .ZN(n657) );
  NAND2_X1 U747 ( .A1(n658), .A2(n657), .ZN(G305) );
  NAND2_X1 U748 ( .A1(G49), .A2(n550), .ZN(n659) );
  XNOR2_X1 U749 ( .A(n659), .B(KEYINPUT80), .ZN(n666) );
  NAND2_X1 U750 ( .A1(G74), .A2(G651), .ZN(n662) );
  NAND2_X1 U751 ( .A1(G87), .A2(n660), .ZN(n661) );
  NAND2_X1 U752 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U753 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U754 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U755 ( .A(KEYINPUT81), .B(n667), .Z(G288) );
  NOR2_X1 U756 ( .A1(G868), .A2(n670), .ZN(n668) );
  XNOR2_X1 U757 ( .A(n668), .B(KEYINPUT87), .ZN(n681) );
  XOR2_X1 U758 ( .A(G305), .B(G288), .Z(n669) );
  XNOR2_X1 U759 ( .A(n670), .B(n669), .ZN(n675) );
  XOR2_X1 U760 ( .A(KEYINPUT85), .B(KEYINPUT19), .Z(n672) );
  XNOR2_X1 U761 ( .A(n964), .B(KEYINPUT86), .ZN(n671) );
  XNOR2_X1 U762 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U763 ( .A(G290), .B(n673), .ZN(n674) );
  XNOR2_X1 U764 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U765 ( .A(G166), .B(n676), .ZN(n677) );
  XNOR2_X1 U766 ( .A(G299), .B(n677), .ZN(n918) );
  XOR2_X1 U767 ( .A(n918), .B(n678), .Z(n679) );
  NAND2_X1 U768 ( .A1(G868), .A2(n679), .ZN(n680) );
  NAND2_X1 U769 ( .A1(n681), .A2(n680), .ZN(G295) );
  XOR2_X1 U770 ( .A(KEYINPUT20), .B(KEYINPUT88), .Z(n683) );
  NAND2_X1 U771 ( .A1(G2084), .A2(G2078), .ZN(n682) );
  XNOR2_X1 U772 ( .A(n683), .B(n682), .ZN(n684) );
  NAND2_X1 U773 ( .A1(G2090), .A2(n684), .ZN(n685) );
  XNOR2_X1 U774 ( .A(KEYINPUT21), .B(n685), .ZN(n686) );
  NAND2_X1 U775 ( .A1(n686), .A2(G2072), .ZN(G158) );
  XOR2_X1 U776 ( .A(KEYINPUT89), .B(G44), .Z(n687) );
  XNOR2_X1 U777 ( .A(KEYINPUT3), .B(n687), .ZN(G218) );
  NOR2_X1 U778 ( .A1(G220), .A2(G219), .ZN(n688) );
  XOR2_X1 U779 ( .A(KEYINPUT22), .B(n688), .Z(n689) );
  NOR2_X1 U780 ( .A1(G218), .A2(n689), .ZN(n690) );
  NAND2_X1 U781 ( .A1(G96), .A2(n690), .ZN(n854) );
  NAND2_X1 U782 ( .A1(n854), .A2(G2106), .ZN(n696) );
  NOR2_X1 U783 ( .A1(G235), .A2(G236), .ZN(n691) );
  XNOR2_X1 U784 ( .A(KEYINPUT90), .B(n691), .ZN(n692) );
  NAND2_X1 U785 ( .A1(n692), .A2(G57), .ZN(n693) );
  NOR2_X1 U786 ( .A1(n693), .A2(G238), .ZN(n694) );
  XNOR2_X1 U787 ( .A(n694), .B(KEYINPUT91), .ZN(n855) );
  NAND2_X1 U788 ( .A1(n855), .A2(G567), .ZN(n695) );
  NAND2_X1 U789 ( .A1(n696), .A2(n695), .ZN(n856) );
  NAND2_X1 U790 ( .A1(G661), .A2(G483), .ZN(n697) );
  XNOR2_X1 U791 ( .A(KEYINPUT92), .B(n697), .ZN(n698) );
  NOR2_X1 U792 ( .A1(n856), .A2(n698), .ZN(n852) );
  NAND2_X1 U793 ( .A1(n852), .A2(G36), .ZN(G176) );
  NOR2_X1 U794 ( .A1(G164), .A2(G1384), .ZN(n780) );
  NAND2_X1 U795 ( .A1(n699), .A2(G40), .ZN(n779) );
  INV_X1 U796 ( .A(n779), .ZN(n700) );
  BUF_X2 U797 ( .A(n720), .Z(n755) );
  NAND2_X1 U798 ( .A1(G1348), .A2(n755), .ZN(n702) );
  INV_X1 U799 ( .A(n755), .ZN(n736) );
  NAND2_X1 U800 ( .A1(G2067), .A2(n736), .ZN(n701) );
  NAND2_X1 U801 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U802 ( .A1(n966), .A2(n703), .ZN(n719) );
  AND2_X1 U803 ( .A1(G1348), .A2(n966), .ZN(n963) );
  INV_X1 U804 ( .A(G1341), .ZN(n990) );
  NOR2_X1 U805 ( .A1(KEYINPUT101), .A2(n990), .ZN(n704) );
  NOR2_X1 U806 ( .A1(n963), .A2(n704), .ZN(n705) );
  NAND2_X1 U807 ( .A1(n705), .A2(KEYINPUT26), .ZN(n706) );
  NAND2_X1 U808 ( .A1(n706), .A2(n755), .ZN(n707) );
  NAND2_X1 U809 ( .A1(n707), .A2(n964), .ZN(n717) );
  NAND2_X1 U810 ( .A1(KEYINPUT26), .A2(G1996), .ZN(n709) );
  NAND2_X1 U811 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U812 ( .A1(KEYINPUT101), .A2(n710), .ZN(n711) );
  NOR2_X1 U813 ( .A1(n755), .A2(n711), .ZN(n715) );
  OR2_X1 U814 ( .A1(G1996), .A2(KEYINPUT26), .ZN(n713) );
  NAND2_X1 U815 ( .A1(KEYINPUT101), .A2(n990), .ZN(n712) );
  NAND2_X1 U816 ( .A1(n713), .A2(n712), .ZN(n714) );
  OR2_X2 U817 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U818 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U819 ( .A1(n719), .A2(n718), .ZN(n729) );
  INV_X1 U820 ( .A(n720), .ZN(n721) );
  NAND2_X1 U821 ( .A1(n721), .A2(G2072), .ZN(n723) );
  NAND2_X1 U822 ( .A1(G1956), .A2(n755), .ZN(n724) );
  NAND2_X1 U823 ( .A1(n725), .A2(n724), .ZN(n730) );
  XNOR2_X1 U824 ( .A(n727), .B(n726), .ZN(n728) );
  NAND2_X1 U825 ( .A1(n729), .A2(n728), .ZN(n733) );
  NAND2_X1 U826 ( .A1(G299), .A2(n730), .ZN(n731) );
  XNOR2_X1 U827 ( .A(n731), .B(KEYINPUT28), .ZN(n732) );
  NAND2_X1 U828 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U829 ( .A(n734), .B(KEYINPUT29), .ZN(n740) );
  NAND2_X1 U830 ( .A1(G1961), .A2(n755), .ZN(n738) );
  XOR2_X1 U831 ( .A(G2078), .B(KEYINPUT25), .Z(n735) );
  XNOR2_X1 U832 ( .A(KEYINPUT100), .B(n735), .ZN(n946) );
  NAND2_X1 U833 ( .A1(n736), .A2(n946), .ZN(n737) );
  NAND2_X1 U834 ( .A1(n738), .A2(n737), .ZN(n747) );
  NOR2_X1 U835 ( .A1(G301), .A2(n747), .ZN(n739) );
  XNOR2_X1 U836 ( .A(n741), .B(KEYINPUT103), .ZN(n753) );
  NOR2_X1 U837 ( .A1(G2084), .A2(n755), .ZN(n764) );
  NOR2_X1 U838 ( .A1(n826), .A2(G1966), .ZN(n742) );
  NAND2_X1 U839 ( .A1(G8), .A2(n765), .ZN(n743) );
  XOR2_X1 U840 ( .A(KEYINPUT30), .B(KEYINPUT104), .Z(n744) );
  XNOR2_X1 U841 ( .A(n745), .B(n744), .ZN(n746) );
  NOR2_X1 U842 ( .A1(G168), .A2(n746), .ZN(n749) );
  AND2_X1 U843 ( .A1(G301), .A2(n747), .ZN(n748) );
  XNOR2_X1 U844 ( .A(n751), .B(n750), .ZN(n752) );
  NAND2_X1 U845 ( .A1(n766), .A2(G286), .ZN(n760) );
  NOR2_X1 U846 ( .A1(G1971), .A2(n826), .ZN(n757) );
  NOR2_X1 U847 ( .A1(G2090), .A2(n755), .ZN(n756) );
  NOR2_X1 U848 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U849 ( .A1(n758), .A2(G303), .ZN(n759) );
  NAND2_X1 U850 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U851 ( .A(n761), .B(KEYINPUT106), .ZN(n762) );
  NAND2_X1 U852 ( .A1(n762), .A2(G8), .ZN(n763) );
  XNOR2_X1 U853 ( .A(n763), .B(KEYINPUT32), .ZN(n770) );
  NAND2_X1 U854 ( .A1(G8), .A2(n764), .ZN(n768) );
  AND2_X1 U855 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U856 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U857 ( .A1(n770), .A2(n769), .ZN(n821) );
  NOR2_X1 U858 ( .A1(G1976), .A2(G288), .ZN(n812) );
  NOR2_X1 U859 ( .A1(G1971), .A2(G303), .ZN(n771) );
  NOR2_X1 U860 ( .A1(n812), .A2(n771), .ZN(n972) );
  NAND2_X1 U861 ( .A1(n821), .A2(n972), .ZN(n773) );
  XNOR2_X1 U862 ( .A(n773), .B(n772), .ZN(n774) );
  NAND2_X1 U863 ( .A1(G1976), .A2(G288), .ZN(n971) );
  NAND2_X1 U864 ( .A1(n774), .A2(n971), .ZN(n775) );
  NOR2_X1 U865 ( .A1(n826), .A2(n775), .ZN(n776) );
  NOR2_X1 U866 ( .A1(KEYINPUT33), .A2(n776), .ZN(n778) );
  XNOR2_X1 U867 ( .A(n778), .B(n777), .ZN(n816) );
  XOR2_X1 U868 ( .A(G1981), .B(G305), .Z(n983) );
  NOR2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n842) );
  XNOR2_X1 U870 ( .A(G2067), .B(KEYINPUT37), .ZN(n840) );
  NAND2_X1 U871 ( .A1(G140), .A2(n893), .ZN(n782) );
  NAND2_X1 U872 ( .A1(G104), .A2(n894), .ZN(n781) );
  NAND2_X1 U873 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U874 ( .A(KEYINPUT34), .B(n783), .ZN(n790) );
  XNOR2_X1 U875 ( .A(KEYINPUT35), .B(KEYINPUT94), .ZN(n788) );
  NAND2_X1 U876 ( .A1(n899), .A2(G116), .ZN(n786) );
  NAND2_X1 U877 ( .A1(n898), .A2(G128), .ZN(n784) );
  XOR2_X1 U878 ( .A(KEYINPUT93), .B(n784), .Z(n785) );
  NAND2_X1 U879 ( .A1(n786), .A2(n785), .ZN(n787) );
  XOR2_X1 U880 ( .A(n788), .B(n787), .Z(n789) );
  NOR2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U882 ( .A(n791), .B(KEYINPUT36), .Z(n792) );
  XNOR2_X1 U883 ( .A(KEYINPUT95), .B(n792), .ZN(n905) );
  NOR2_X1 U884 ( .A1(n840), .A2(n905), .ZN(n1022) );
  NAND2_X1 U885 ( .A1(n842), .A2(n1022), .ZN(n838) );
  XNOR2_X1 U886 ( .A(n842), .B(KEYINPUT96), .ZN(n808) );
  NAND2_X1 U887 ( .A1(G129), .A2(n898), .ZN(n794) );
  NAND2_X1 U888 ( .A1(G117), .A2(n899), .ZN(n793) );
  NAND2_X1 U889 ( .A1(n794), .A2(n793), .ZN(n797) );
  NAND2_X1 U890 ( .A1(n894), .A2(G105), .ZN(n795) );
  XOR2_X1 U891 ( .A(KEYINPUT38), .B(n795), .Z(n796) );
  NOR2_X1 U892 ( .A1(n797), .A2(n796), .ZN(n799) );
  NAND2_X1 U893 ( .A1(n893), .A2(G141), .ZN(n798) );
  NAND2_X1 U894 ( .A1(n799), .A2(n798), .ZN(n890) );
  NAND2_X1 U895 ( .A1(G1996), .A2(n890), .ZN(n807) );
  NAND2_X1 U896 ( .A1(G131), .A2(n893), .ZN(n801) );
  NAND2_X1 U897 ( .A1(G119), .A2(n898), .ZN(n800) );
  NAND2_X1 U898 ( .A1(n801), .A2(n800), .ZN(n805) );
  NAND2_X1 U899 ( .A1(n899), .A2(G107), .ZN(n803) );
  NAND2_X1 U900 ( .A1(G95), .A2(n894), .ZN(n802) );
  NAND2_X1 U901 ( .A1(n803), .A2(n802), .ZN(n804) );
  OR2_X1 U902 ( .A1(n805), .A2(n804), .ZN(n908) );
  NAND2_X1 U903 ( .A1(G1991), .A2(n908), .ZN(n806) );
  NAND2_X1 U904 ( .A1(n807), .A2(n806), .ZN(n1028) );
  NAND2_X1 U905 ( .A1(n808), .A2(n1028), .ZN(n809) );
  XNOR2_X1 U906 ( .A(n809), .B(KEYINPUT97), .ZN(n835) );
  INV_X1 U907 ( .A(n835), .ZN(n810) );
  AND2_X1 U908 ( .A1(n838), .A2(n810), .ZN(n818) );
  AND2_X1 U909 ( .A1(n983), .A2(n818), .ZN(n811) );
  XNOR2_X1 U910 ( .A(G1986), .B(G290), .ZN(n968) );
  NAND2_X1 U911 ( .A1(n968), .A2(n842), .ZN(n817) );
  AND2_X1 U912 ( .A1(n811), .A2(n817), .ZN(n814) );
  NAND2_X1 U913 ( .A1(n812), .A2(KEYINPUT33), .ZN(n813) );
  NAND2_X1 U914 ( .A1(n816), .A2(n815), .ZN(n847) );
  INV_X1 U915 ( .A(n817), .ZN(n832) );
  INV_X1 U916 ( .A(n818), .ZN(n830) );
  NOR2_X1 U917 ( .A1(G2090), .A2(G303), .ZN(n819) );
  NAND2_X1 U918 ( .A1(G8), .A2(n819), .ZN(n820) );
  NAND2_X1 U919 ( .A1(n821), .A2(n820), .ZN(n822) );
  AND2_X1 U920 ( .A1(n822), .A2(n826), .ZN(n828) );
  NOR2_X1 U921 ( .A1(G1981), .A2(G305), .ZN(n823) );
  XOR2_X1 U922 ( .A(n823), .B(KEYINPUT24), .Z(n824) );
  XNOR2_X1 U923 ( .A(KEYINPUT98), .B(n824), .ZN(n825) );
  NOR2_X1 U924 ( .A1(n826), .A2(n825), .ZN(n827) );
  NOR2_X1 U925 ( .A1(n828), .A2(n827), .ZN(n829) );
  OR2_X1 U926 ( .A1(n832), .A2(n831), .ZN(n845) );
  NOR2_X1 U927 ( .A1(G1996), .A2(n890), .ZN(n1019) );
  NOR2_X1 U928 ( .A1(G1991), .A2(n908), .ZN(n1024) );
  NOR2_X1 U929 ( .A1(G1986), .A2(G290), .ZN(n833) );
  NOR2_X1 U930 ( .A1(n1024), .A2(n833), .ZN(n834) );
  NOR2_X1 U931 ( .A1(n835), .A2(n834), .ZN(n836) );
  NOR2_X1 U932 ( .A1(n1019), .A2(n836), .ZN(n837) );
  XNOR2_X1 U933 ( .A(n837), .B(KEYINPUT39), .ZN(n839) );
  NAND2_X1 U934 ( .A1(n839), .A2(n838), .ZN(n841) );
  NAND2_X1 U935 ( .A1(n840), .A2(n905), .ZN(n1037) );
  NAND2_X1 U936 ( .A1(n841), .A2(n1037), .ZN(n843) );
  NAND2_X1 U937 ( .A1(n843), .A2(n842), .ZN(n844) );
  AND2_X1 U938 ( .A1(n845), .A2(n844), .ZN(n846) );
  NAND2_X1 U939 ( .A1(n847), .A2(n846), .ZN(n848) );
  XNOR2_X1 U940 ( .A(n848), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U941 ( .A1(G2106), .A2(n849), .ZN(G217) );
  AND2_X1 U942 ( .A1(G15), .A2(G2), .ZN(n850) );
  NAND2_X1 U943 ( .A1(G661), .A2(n850), .ZN(G259) );
  NAND2_X1 U944 ( .A1(G3), .A2(G1), .ZN(n851) );
  NAND2_X1 U945 ( .A1(n852), .A2(n851), .ZN(n853) );
  XNOR2_X1 U946 ( .A(KEYINPUT112), .B(n853), .ZN(G188) );
  INV_X1 U948 ( .A(G96), .ZN(G221) );
  INV_X1 U949 ( .A(G57), .ZN(G237) );
  NOR2_X1 U950 ( .A1(n855), .A2(n854), .ZN(G325) );
  INV_X1 U951 ( .A(G325), .ZN(G261) );
  INV_X1 U952 ( .A(n856), .ZN(G319) );
  XOR2_X1 U953 ( .A(KEYINPUT42), .B(G2090), .Z(n858) );
  XNOR2_X1 U954 ( .A(G2067), .B(G2084), .ZN(n857) );
  XNOR2_X1 U955 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U956 ( .A(n859), .B(G2100), .Z(n861) );
  XNOR2_X1 U957 ( .A(G2078), .B(G2072), .ZN(n860) );
  XNOR2_X1 U958 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U959 ( .A(G2096), .B(KEYINPUT43), .Z(n863) );
  XNOR2_X1 U960 ( .A(KEYINPUT113), .B(G2678), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U962 ( .A(n865), .B(n864), .Z(G227) );
  XOR2_X1 U963 ( .A(G1971), .B(G1956), .Z(n867) );
  XNOR2_X1 U964 ( .A(G1986), .B(G1961), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U966 ( .A(n868), .B(KEYINPUT41), .Z(n870) );
  XNOR2_X1 U967 ( .A(G1996), .B(G1991), .ZN(n869) );
  XNOR2_X1 U968 ( .A(n870), .B(n869), .ZN(n874) );
  XOR2_X1 U969 ( .A(G2474), .B(G1976), .Z(n872) );
  XNOR2_X1 U970 ( .A(G1966), .B(G1981), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(n873) );
  XNOR2_X1 U972 ( .A(n874), .B(n873), .ZN(G229) );
  NAND2_X1 U973 ( .A1(n898), .A2(G124), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n875), .B(KEYINPUT44), .ZN(n877) );
  NAND2_X1 U975 ( .A1(G112), .A2(n899), .ZN(n876) );
  NAND2_X1 U976 ( .A1(n877), .A2(n876), .ZN(n881) );
  NAND2_X1 U977 ( .A1(G136), .A2(n893), .ZN(n879) );
  NAND2_X1 U978 ( .A1(G100), .A2(n894), .ZN(n878) );
  NAND2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n880) );
  NOR2_X1 U980 ( .A1(n881), .A2(n880), .ZN(G162) );
  NAND2_X1 U981 ( .A1(G130), .A2(n898), .ZN(n883) );
  NAND2_X1 U982 ( .A1(G118), .A2(n899), .ZN(n882) );
  NAND2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n888) );
  NAND2_X1 U984 ( .A1(G142), .A2(n893), .ZN(n885) );
  NAND2_X1 U985 ( .A1(G106), .A2(n894), .ZN(n884) );
  NAND2_X1 U986 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U987 ( .A(KEYINPUT45), .B(n886), .Z(n887) );
  NOR2_X1 U988 ( .A1(n888), .A2(n887), .ZN(n892) );
  XOR2_X1 U989 ( .A(G160), .B(n1023), .Z(n889) );
  XNOR2_X1 U990 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U991 ( .A(n892), .B(n891), .ZN(n907) );
  NAND2_X1 U992 ( .A1(G139), .A2(n893), .ZN(n896) );
  NAND2_X1 U993 ( .A1(G103), .A2(n894), .ZN(n895) );
  NAND2_X1 U994 ( .A1(n896), .A2(n895), .ZN(n897) );
  XNOR2_X1 U995 ( .A(KEYINPUT114), .B(n897), .ZN(n904) );
  NAND2_X1 U996 ( .A1(G127), .A2(n898), .ZN(n901) );
  NAND2_X1 U997 ( .A1(G115), .A2(n899), .ZN(n900) );
  NAND2_X1 U998 ( .A1(n901), .A2(n900), .ZN(n902) );
  XOR2_X1 U999 ( .A(KEYINPUT47), .B(n902), .Z(n903) );
  NOR2_X1 U1000 ( .A1(n904), .A2(n903), .ZN(n1031) );
  XNOR2_X1 U1001 ( .A(n905), .B(n1031), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n907), .B(n906), .ZN(n913) );
  XNOR2_X1 U1003 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n910) );
  XNOR2_X1 U1004 ( .A(n908), .B(G162), .ZN(n909) );
  XNOR2_X1 U1005 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1006 ( .A(G164), .B(n911), .Z(n912) );
  XNOR2_X1 U1007 ( .A(n913), .B(n912), .ZN(n914) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n914), .ZN(n915) );
  XOR2_X1 U1009 ( .A(KEYINPUT115), .B(n915), .Z(G395) );
  XOR2_X1 U1010 ( .A(KEYINPUT116), .B(G286), .Z(n917) );
  XNOR2_X1 U1011 ( .A(G171), .B(n966), .ZN(n916) );
  XNOR2_X1 U1012 ( .A(n917), .B(n916), .ZN(n919) );
  XNOR2_X1 U1013 ( .A(n919), .B(n918), .ZN(n920) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n920), .ZN(n921) );
  XOR2_X1 U1015 ( .A(KEYINPUT117), .B(n921), .Z(G397) );
  XOR2_X1 U1016 ( .A(KEYINPUT110), .B(G2443), .Z(n923) );
  XNOR2_X1 U1017 ( .A(G2451), .B(G2427), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(n923), .B(n922), .ZN(n924) );
  XOR2_X1 U1019 ( .A(n924), .B(G2430), .Z(n926) );
  XNOR2_X1 U1020 ( .A(G1348), .B(G1341), .ZN(n925) );
  XNOR2_X1 U1021 ( .A(n926), .B(n925), .ZN(n930) );
  XOR2_X1 U1022 ( .A(G2435), .B(KEYINPUT111), .Z(n928) );
  XNOR2_X1 U1023 ( .A(G2438), .B(G2454), .ZN(n927) );
  XNOR2_X1 U1024 ( .A(n928), .B(n927), .ZN(n929) );
  XOR2_X1 U1025 ( .A(n930), .B(n929), .Z(n932) );
  XNOR2_X1 U1026 ( .A(G2446), .B(KEYINPUT109), .ZN(n931) );
  XNOR2_X1 U1027 ( .A(n932), .B(n931), .ZN(n933) );
  NAND2_X1 U1028 ( .A1(n933), .A2(G14), .ZN(n939) );
  NAND2_X1 U1029 ( .A1(G319), .A2(n939), .ZN(n936) );
  NOR2_X1 U1030 ( .A1(G227), .A2(G229), .ZN(n934) );
  XNOR2_X1 U1031 ( .A(KEYINPUT49), .B(n934), .ZN(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n938) );
  NOR2_X1 U1033 ( .A1(G395), .A2(G397), .ZN(n937) );
  NAND2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(G225) );
  INV_X1 U1035 ( .A(G225), .ZN(G308) );
  INV_X1 U1036 ( .A(n939), .ZN(G401) );
  XOR2_X1 U1037 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n1048) );
  INV_X1 U1038 ( .A(KEYINPUT55), .ZN(n1042) );
  XNOR2_X1 U1039 ( .A(G2084), .B(G34), .ZN(n940) );
  XNOR2_X1 U1040 ( .A(n940), .B(KEYINPUT54), .ZN(n942) );
  XNOR2_X1 U1041 ( .A(G35), .B(G2090), .ZN(n941) );
  NOR2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n956) );
  XOR2_X1 U1043 ( .A(G1996), .B(G32), .Z(n943) );
  NAND2_X1 U1044 ( .A1(n943), .A2(G28), .ZN(n952) );
  XNOR2_X1 U1045 ( .A(G1991), .B(G25), .ZN(n945) );
  XNOR2_X1 U1046 ( .A(G2072), .B(G33), .ZN(n944) );
  NOR2_X1 U1047 ( .A1(n945), .A2(n944), .ZN(n950) );
  XNOR2_X1 U1048 ( .A(n946), .B(G27), .ZN(n948) );
  XNOR2_X1 U1049 ( .A(G2067), .B(G26), .ZN(n947) );
  NOR2_X1 U1050 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1052 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1053 ( .A(n953), .B(KEYINPUT120), .Z(n954) );
  XNOR2_X1 U1054 ( .A(KEYINPUT53), .B(n954), .ZN(n955) );
  NAND2_X1 U1055 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1056 ( .A(n1042), .B(n957), .ZN(n959) );
  INV_X1 U1057 ( .A(G29), .ZN(n958) );
  NAND2_X1 U1058 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1059 ( .A1(G11), .A2(n960), .ZN(n1017) );
  XNOR2_X1 U1060 ( .A(G16), .B(KEYINPUT56), .ZN(n989) );
  XNOR2_X1 U1061 ( .A(G171), .B(G1961), .ZN(n961) );
  XNOR2_X1 U1062 ( .A(n961), .B(KEYINPUT121), .ZN(n962) );
  NOR2_X1 U1063 ( .A1(n963), .A2(n962), .ZN(n979) );
  XNOR2_X1 U1064 ( .A(n990), .B(n964), .ZN(n965) );
  XNOR2_X1 U1065 ( .A(n965), .B(KEYINPUT123), .ZN(n970) );
  NOR2_X1 U1066 ( .A1(G1348), .A2(n966), .ZN(n967) );
  NOR2_X1 U1067 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1068 ( .A1(n970), .A2(n969), .ZN(n977) );
  NAND2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n974) );
  AND2_X1 U1070 ( .A1(G303), .A2(G1971), .ZN(n973) );
  NOR2_X1 U1071 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1072 ( .A(KEYINPUT122), .B(n975), .Z(n976) );
  NOR2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n981) );
  XNOR2_X1 U1075 ( .A(G1956), .B(G299), .ZN(n980) );
  NOR2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1077 ( .A(KEYINPUT124), .B(n982), .ZN(n987) );
  XNOR2_X1 U1078 ( .A(G1966), .B(G168), .ZN(n984) );
  NAND2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1080 ( .A(KEYINPUT57), .B(n985), .ZN(n986) );
  NAND2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n1015) );
  INV_X1 U1083 ( .A(G16), .ZN(n1013) );
  XNOR2_X1 U1084 ( .A(G19), .B(n990), .ZN(n994) );
  XNOR2_X1 U1085 ( .A(G1956), .B(G20), .ZN(n992) );
  XNOR2_X1 U1086 ( .A(G1981), .B(G6), .ZN(n991) );
  NOR2_X1 U1087 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n997) );
  XOR2_X1 U1089 ( .A(KEYINPUT59), .B(G1348), .Z(n995) );
  XNOR2_X1 U1090 ( .A(G4), .B(n995), .ZN(n996) );
  NOR2_X1 U1091 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1092 ( .A(KEYINPUT60), .B(n998), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(G1966), .B(G21), .ZN(n1000) );
  XNOR2_X1 U1094 ( .A(G5), .B(G1961), .ZN(n999) );
  NOR2_X1 U1095 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1096 ( .A1(n1002), .A2(n1001), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(G1986), .B(G24), .ZN(n1004) );
  XNOR2_X1 U1098 ( .A(G22), .B(G1971), .ZN(n1003) );
  NOR2_X1 U1099 ( .A1(n1004), .A2(n1003), .ZN(n1007) );
  XNOR2_X1 U1100 ( .A(G1976), .B(KEYINPUT125), .ZN(n1005) );
  XNOR2_X1 U1101 ( .A(n1005), .B(G23), .ZN(n1006) );
  NAND2_X1 U1102 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1103 ( .A(KEYINPUT58), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1104 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1105 ( .A(KEYINPUT61), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1106 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1107 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1108 ( .A1(n1017), .A2(n1016), .ZN(n1046) );
  XOR2_X1 U1109 ( .A(G2090), .B(G162), .Z(n1018) );
  NOR2_X1 U1110 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1111 ( .A(n1020), .B(KEYINPUT51), .ZN(n1021) );
  NOR2_X1 U1112 ( .A1(n1022), .A2(n1021), .ZN(n1030) );
  XNOR2_X1 U1113 ( .A(G160), .B(G2084), .ZN(n1026) );
  NOR2_X1 U1114 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1115 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1116 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1040) );
  XOR2_X1 U1118 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n1036) );
  XOR2_X1 U1119 ( .A(G2072), .B(n1031), .Z(n1033) );
  XOR2_X1 U1120 ( .A(G164), .B(G2078), .Z(n1032) );
  NOR2_X1 U1121 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1122 ( .A(n1034), .B(KEYINPUT50), .ZN(n1035) );
  XNOR2_X1 U1123 ( .A(n1036), .B(n1035), .ZN(n1038) );
  NAND2_X1 U1124 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NOR2_X1 U1125 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XNOR2_X1 U1126 ( .A(KEYINPUT52), .B(n1041), .ZN(n1043) );
  NAND2_X1 U1127 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  NAND2_X1 U1128 ( .A1(n1044), .A2(G29), .ZN(n1045) );
  NAND2_X1 U1129 ( .A1(n1046), .A2(n1045), .ZN(n1047) );
  XNOR2_X1 U1130 ( .A(n1048), .B(n1047), .ZN(G311) );
  XNOR2_X1 U1131 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

