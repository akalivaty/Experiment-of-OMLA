//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT28), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(KEYINPUT1), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  OAI22_X1  g008(.A1(new_n190), .A2(new_n192), .B1(new_n194), .B2(G128), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  XNOR2_X1  g011(.A(G143), .B(G146), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(new_n190), .ZN(new_n199));
  AND4_X1   g013(.A1(new_n197), .A2(new_n190), .A3(new_n194), .A4(new_n192), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n196), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT67), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n190), .A2(new_n194), .A3(new_n192), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT64), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n198), .A2(new_n197), .A3(new_n190), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n195), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT67), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G134), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G137), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n209), .A2(G137), .ZN(new_n212));
  OAI21_X1  g026(.A(G131), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT11), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n214), .B1(new_n209), .B2(G137), .ZN(new_n215));
  INV_X1    g029(.A(G137), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(KEYINPUT11), .A3(G134), .ZN(new_n217));
  INV_X1    g031(.A(G131), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n215), .A2(new_n217), .A3(new_n218), .A4(new_n210), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n202), .A2(new_n208), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT68), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n215), .A2(new_n217), .A3(new_n210), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G131), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n225), .A2(KEYINPUT66), .A3(new_n219), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT66), .B1(new_n225), .B2(new_n219), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AND2_X1   g042(.A1(KEYINPUT0), .A2(G128), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n194), .A2(new_n192), .A3(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT0), .B(G128), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n198), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT65), .ZN(new_n234));
  INV_X1    g048(.A(G116), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n234), .B1(new_n235), .B2(G119), .ZN(new_n236));
  INV_X1    g050(.A(G119), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(KEYINPUT65), .A3(G116), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n235), .A2(G119), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n236), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G113), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT2), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT2), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G113), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n242), .A2(new_n244), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n247), .A2(new_n236), .A3(new_n238), .A4(new_n239), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n246), .A2(new_n248), .A3(KEYINPUT69), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n246), .A2(new_n248), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n228), .A2(new_n233), .B1(new_n249), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n202), .A2(new_n208), .A3(new_n254), .A4(new_n221), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n223), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n225), .A2(new_n219), .ZN(new_n257));
  OAI22_X1  g071(.A1(new_n257), .A2(new_n232), .B1(new_n206), .B2(new_n220), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n250), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n188), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT28), .B1(new_n253), .B2(new_n222), .ZN(new_n261));
  OR2_X1    g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  XOR2_X1   g076(.A(KEYINPUT26), .B(G101), .Z(new_n263));
  INV_X1    g077(.A(G237), .ZN(new_n264));
  INV_X1    g078(.A(G953), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n264), .A2(new_n265), .A3(G210), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n263), .B(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n268));
  XOR2_X1   g082(.A(new_n267), .B(new_n268), .Z(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT31), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT30), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n272), .B1(new_n228), .B2(new_n233), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n223), .A2(new_n273), .A3(new_n255), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n258), .A2(new_n272), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n275), .A2(new_n250), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n256), .A2(new_n269), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n271), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n274), .A2(new_n276), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n280), .A2(KEYINPUT31), .A3(new_n256), .A4(new_n269), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n262), .A2(new_n270), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(G472), .A2(G902), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n283), .B(KEYINPUT71), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n187), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT32), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n279), .A2(new_n281), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n270), .B1(new_n260), .B2(new_n261), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n284), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n289), .A2(KEYINPUT72), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n285), .A2(new_n286), .A3(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n284), .A2(new_n286), .ZN(new_n293));
  AOI21_X1  g107(.A(KEYINPUT73), .B1(new_n289), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT73), .ZN(new_n295));
  INV_X1    g109(.A(new_n293), .ZN(new_n296));
  AOI211_X1 g110(.A(new_n295), .B(new_n296), .C1(new_n287), .C2(new_n288), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n261), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n270), .A2(new_n300), .ZN(new_n301));
  AND2_X1   g115(.A1(new_n223), .A2(new_n255), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n228), .A2(new_n233), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n223), .A2(new_n303), .A3(new_n255), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n252), .A2(new_n249), .ZN(new_n305));
  AOI22_X1  g119(.A1(new_n302), .A2(new_n253), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n299), .B(new_n301), .C1(new_n306), .C2(new_n188), .ZN(new_n307));
  INV_X1    g121(.A(G902), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n302), .A2(new_n253), .B1(new_n274), .B2(new_n276), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n300), .B1(new_n309), .B2(new_n269), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n260), .A2(new_n261), .A3(new_n270), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n307), .B(new_n308), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G472), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n292), .A2(new_n298), .A3(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(G214), .B1(G237), .B2(G902), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT83), .ZN(new_n317));
  INV_X1    g131(.A(G104), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT3), .B1(new_n318), .B2(G107), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT3), .ZN(new_n320));
  INV_X1    g134(.A(G107), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(G104), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n318), .A2(G107), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n319), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G101), .ZN(new_n325));
  AND2_X1   g139(.A1(KEYINPUT78), .A2(G101), .ZN(new_n326));
  NOR2_X1   g140(.A1(KEYINPUT78), .A2(G101), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n328), .A2(new_n319), .A3(new_n322), .A4(new_n323), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n325), .A2(KEYINPUT4), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT4), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n324), .A2(new_n331), .A3(G101), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n330), .A2(new_n250), .A3(new_n332), .ZN(new_n333));
  NOR3_X1   g147(.A1(new_n235), .A2(KEYINPUT5), .A3(G119), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(new_n241), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT5), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n335), .B1(new_n240), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n323), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n318), .A2(G107), .ZN(new_n339));
  OAI21_X1  g153(.A(G101), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n337), .A2(new_n248), .A3(new_n329), .A4(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n333), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT6), .ZN(new_n343));
  XNOR2_X1  g157(.A(G110), .B(G122), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n344), .A2(KEYINPUT80), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n342), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n333), .A2(new_n341), .A3(new_n344), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT6), .ZN(new_n348));
  INV_X1    g162(.A(new_n345), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n349), .B1(new_n333), .B2(new_n341), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n346), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT81), .ZN(new_n352));
  AND3_X1   g166(.A1(new_n232), .A2(new_n352), .A3(G125), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n352), .B1(new_n232), .B2(G125), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G125), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n356), .B(new_n196), .C1(new_n199), .C2(new_n200), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n265), .A2(G224), .ZN(new_n359));
  XOR2_X1   g173(.A(new_n359), .B(KEYINPUT82), .Z(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n355), .A2(new_n357), .A3(new_n360), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n317), .B1(new_n351), .B2(new_n364), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n355), .A2(new_n357), .A3(new_n360), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n360), .B1(new_n355), .B2(new_n357), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n342), .A2(new_n345), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(KEYINPUT6), .A3(new_n347), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n368), .A2(new_n370), .A3(KEYINPUT83), .A4(new_n346), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n359), .A2(KEYINPUT7), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n355), .A2(KEYINPUT84), .A3(new_n357), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n232), .A2(G125), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT81), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n232), .A2(new_n352), .A3(G125), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n377), .A2(new_n357), .A3(new_n378), .A4(new_n374), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n337), .A2(new_n248), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n329), .A2(new_n340), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n341), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n344), .B(KEYINPUT8), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n375), .A2(new_n381), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n357), .A2(new_n376), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n373), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n347), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n308), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT85), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT85), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n394), .B(new_n308), .C1(new_n388), .C2(new_n391), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n372), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(G210), .B1(G237), .B2(G902), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n372), .A2(new_n397), .A3(new_n393), .A4(new_n395), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n316), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(G221), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT9), .B(G234), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n402), .B1(new_n404), .B2(new_n308), .ZN(new_n405));
  INV_X1    g219(.A(G469), .ZN(new_n406));
  XNOR2_X1  g220(.A(G110), .B(G140), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n265), .A2(G227), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n407), .B(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n329), .A2(KEYINPUT10), .A3(new_n340), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n202), .A2(new_n208), .A3(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT10), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n414), .B1(new_n206), .B2(new_n383), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n330), .A2(new_n233), .A3(new_n332), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n228), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT79), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI211_X1 g234(.A(KEYINPUT79), .B(new_n228), .C1(new_n413), .C2(new_n417), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n228), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n202), .A2(new_n208), .A3(new_n412), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n423), .A2(new_n424), .A3(new_n415), .A4(new_n416), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n410), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n201), .A2(new_n329), .A3(new_n340), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n206), .A2(new_n383), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(KEYINPUT12), .B1(new_n429), .B2(new_n228), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT12), .ZN(new_n431));
  AOI211_X1 g245(.A(new_n431), .B(new_n257), .C1(new_n427), .C2(new_n428), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n425), .A2(new_n410), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n406), .B(new_n308), .C1(new_n426), .C2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n434), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n425), .B1(new_n430), .B2(new_n432), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n422), .A2(new_n437), .B1(new_n409), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(G469), .B1(new_n439), .B2(G902), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n405), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G478), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(KEYINPUT15), .ZN(new_n443));
  INV_X1    g257(.A(G217), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n403), .A2(new_n444), .A3(G953), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G122), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G116), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n321), .B1(new_n448), .B2(KEYINPUT14), .ZN(new_n449));
  XNOR2_X1  g263(.A(G116), .B(G122), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n449), .B(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(G128), .B(G143), .ZN(new_n453));
  OR2_X1    g267(.A1(new_n453), .A2(KEYINPUT90), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(KEYINPUT90), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n209), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n454), .A2(G134), .A3(new_n455), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n452), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n453), .A2(KEYINPUT13), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n191), .A2(G128), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n460), .B(G134), .C1(KEYINPUT13), .C2(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n450), .B(new_n321), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n464), .B1(new_n209), .B2(new_n456), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n446), .B1(new_n459), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n457), .A2(new_n458), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n451), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n457), .A2(new_n462), .A3(new_n463), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n469), .A3(new_n445), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(KEYINPUT91), .B1(new_n471), .B2(new_n308), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT91), .ZN(new_n473));
  AOI211_X1 g287(.A(new_n473), .B(G902), .C1(new_n466), .C2(new_n470), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n443), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(G902), .B1(new_n466), .B2(new_n470), .ZN(new_n476));
  OAI22_X1  g290(.A1(new_n476), .A2(KEYINPUT91), .B1(KEYINPUT15), .B2(new_n442), .ZN(new_n477));
  INV_X1    g291(.A(G952), .ZN(new_n478));
  AOI211_X1 g292(.A(G953), .B(new_n478), .C1(G234), .C2(G237), .ZN(new_n479));
  AOI211_X1 g293(.A(new_n308), .B(new_n265), .C1(G234), .C2(G237), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT21), .B(G898), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n475), .A2(new_n477), .A3(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(G125), .B(G140), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT16), .ZN(new_n486));
  OR3_X1    g300(.A1(new_n356), .A2(KEYINPUT16), .A3(G140), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(G146), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n193), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT87), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n264), .A2(new_n265), .A3(G214), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n191), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n264), .A2(new_n265), .A3(G143), .A4(G214), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n493), .B1(new_n497), .B2(G131), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT17), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n495), .A2(KEYINPUT87), .A3(new_n218), .A4(new_n496), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n497), .A2(G131), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n498), .A2(new_n499), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n497), .A2(KEYINPUT17), .A3(G131), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n492), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(G113), .B(G122), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT89), .B(G104), .ZN(new_n506));
  XOR2_X1   g320(.A(new_n505), .B(new_n506), .Z(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n485), .B(G146), .ZN(new_n509));
  OR2_X1    g323(.A1(new_n509), .A2(KEYINPUT86), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(KEYINPUT86), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(KEYINPUT18), .A2(G131), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n497), .B(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n504), .A2(new_n508), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n508), .B1(new_n504), .B2(new_n515), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n308), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(G475), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT20), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT19), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n485), .B1(KEYINPUT88), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n522), .B1(new_n485), .B2(new_n523), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n524), .A2(G146), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(new_n490), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n515), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n507), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n504), .A2(new_n508), .A3(new_n515), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(G475), .A2(G902), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n520), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n532), .ZN(new_n534));
  AOI211_X1 g348(.A(KEYINPUT20), .B(new_n534), .C1(new_n529), .C2(new_n530), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n519), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n484), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n401), .A2(new_n441), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT92), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT22), .B(G137), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n265), .A2(G221), .A3(G234), .ZN(new_n542));
  XOR2_X1   g356(.A(new_n541), .B(new_n542), .Z(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  AND2_X1   g358(.A1(new_n485), .A2(new_n193), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n545), .B1(new_n489), .B2(G146), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT74), .B1(new_n189), .B2(G119), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT74), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n548), .A2(new_n237), .A3(G128), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n547), .B(new_n549), .C1(new_n237), .C2(G128), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT24), .B(G110), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n550), .A2(KEYINPUT75), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n237), .A2(G128), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n189), .A2(KEYINPUT23), .A3(G119), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n237), .A2(G128), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n553), .B(new_n554), .C1(new_n555), .C2(KEYINPUT23), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n552), .B1(G110), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT75), .B1(new_n550), .B2(new_n551), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n546), .B(KEYINPUT76), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n558), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n561), .B(new_n552), .C1(G110), .C2(new_n556), .ZN(new_n562));
  AOI21_X1  g376(.A(KEYINPUT76), .B1(new_n562), .B2(new_n546), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n556), .A2(G110), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n565), .B1(new_n551), .B2(new_n550), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n492), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n544), .B1(new_n564), .B2(new_n567), .ZN(new_n568));
  OAI221_X1 g382(.A(new_n543), .B1(new_n492), .B2(new_n566), .C1(new_n560), .C2(new_n563), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n444), .B1(G234), .B2(new_n308), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(G902), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n568), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(KEYINPUT77), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n568), .A2(new_n308), .A3(new_n569), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT25), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT25), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n568), .A2(new_n576), .A3(new_n308), .A4(new_n569), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n575), .A2(new_n577), .A3(new_n570), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n401), .A2(new_n441), .A3(KEYINPUT92), .A4(new_n537), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n314), .A2(new_n540), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  XOR2_X1   g396(.A(new_n582), .B(new_n328), .Z(G3));
  AND2_X1   g397(.A1(new_n580), .A2(new_n441), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n285), .A2(new_n291), .ZN(new_n585));
  INV_X1    g399(.A(G472), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n586), .B1(new_n289), .B2(new_n308), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n395), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n347), .A2(new_n390), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n590), .A2(new_n375), .A3(new_n387), .A4(new_n381), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n394), .B1(new_n591), .B2(new_n308), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n397), .B1(new_n593), .B2(new_n372), .ZN(new_n594));
  AND4_X1   g408(.A1(new_n397), .A2(new_n372), .A3(new_n393), .A4(new_n395), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n315), .B(new_n483), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT33), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT93), .ZN(new_n598));
  OR2_X1    g412(.A1(new_n597), .A2(KEYINPUT93), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n471), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n466), .A2(new_n470), .A3(KEYINPUT93), .A4(new_n597), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n308), .A2(G478), .ZN(new_n604));
  OAI22_X1  g418(.A1(new_n603), .A2(new_n604), .B1(G478), .B2(new_n476), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n536), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n596), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n584), .A2(new_n588), .A3(new_n607), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT34), .B(G104), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G6));
  INV_X1    g424(.A(KEYINPUT95), .ZN(new_n611));
  AOI22_X1  g425(.A1(new_n475), .A2(new_n477), .B1(G475), .B2(new_n518), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n531), .A2(new_n520), .A3(new_n532), .ZN(new_n613));
  OR2_X1    g427(.A1(new_n613), .A2(KEYINPUT94), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n508), .B1(new_n515), .B2(new_n527), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n532), .B1(new_n516), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT20), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n617), .A2(KEYINPUT94), .A3(new_n613), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n612), .A2(new_n614), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n611), .B1(new_n596), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n475), .A2(new_n477), .ZN(new_n621));
  AND4_X1   g435(.A1(new_n519), .A2(new_n614), .A3(new_n621), .A4(new_n618), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n622), .A2(new_n401), .A3(KEYINPUT95), .A4(new_n483), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n624), .A2(new_n588), .A3(new_n584), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(new_n321), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT96), .B(KEYINPUT35), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G9));
  NOR2_X1   g442(.A1(new_n564), .A2(new_n567), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n544), .A2(KEYINPUT36), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n629), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n571), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n578), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n540), .A2(new_n588), .A3(new_n581), .A4(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT37), .B(G110), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(KEYINPUT97), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n635), .B(new_n637), .ZN(G12));
  AND3_X1   g452(.A1(new_n401), .A2(new_n441), .A3(new_n634), .ZN(new_n639));
  INV_X1    g453(.A(G900), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n479), .B1(new_n480), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n612), .A2(new_n614), .A3(new_n618), .A4(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n285), .A2(new_n286), .A3(new_n291), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n295), .B1(new_n282), .B2(new_n296), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n289), .A2(KEYINPUT73), .A3(new_n293), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n646), .A2(new_n313), .A3(new_n647), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n639), .B(new_n644), .C1(new_n645), .C2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(KEYINPUT98), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT98), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n314), .A2(new_n651), .A3(new_n639), .A4(new_n644), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G128), .ZN(G30));
  NOR2_X1   g468(.A1(new_n306), .A2(new_n269), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n277), .A2(new_n278), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n308), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(G472), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n292), .A2(new_n298), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT99), .ZN(new_n660));
  INV_X1    g474(.A(new_n536), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n475), .A2(new_n477), .ZN(new_n662));
  NOR4_X1   g476(.A1(new_n634), .A2(new_n316), .A3(new_n661), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT100), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n399), .A2(new_n400), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT38), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n641), .B(KEYINPUT39), .Z(new_n667));
  NAND2_X1  g481(.A1(new_n441), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n668), .B(KEYINPUT40), .Z(new_n669));
  NAND4_X1  g483(.A1(new_n660), .A2(new_n664), .A3(new_n666), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G143), .ZN(G45));
  NOR2_X1   g485(.A1(new_n606), .A2(new_n641), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n314), .A2(new_n639), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G146), .ZN(G48));
  NAND2_X1  g488(.A1(new_n422), .A2(new_n425), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n435), .B1(new_n675), .B2(new_n409), .ZN(new_n676));
  OAI21_X1  g490(.A(G469), .B1(new_n676), .B2(G902), .ZN(new_n677));
  INV_X1    g491(.A(new_n405), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n677), .A2(new_n678), .A3(new_n436), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n314), .A2(new_n580), .A3(new_n607), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT41), .B(G113), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G15));
  NAND4_X1  g497(.A1(new_n624), .A2(new_n314), .A3(new_n580), .A4(new_n680), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G116), .ZN(G18));
  NAND2_X1  g499(.A1(new_n634), .A2(new_n537), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n315), .B1(new_n594), .B2(new_n595), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n686), .A2(new_n679), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n314), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G119), .ZN(G21));
  AOI21_X1  g504(.A(new_n316), .B1(new_n475), .B2(new_n477), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n665), .A2(new_n536), .A3(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n677), .A2(new_n678), .A3(new_n436), .A4(new_n483), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n299), .B1(new_n306), .B2(new_n188), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n270), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n284), .B1(new_n696), .B2(new_n287), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n579), .A2(new_n587), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G122), .ZN(G24));
  AND2_X1   g514(.A1(new_n578), .A2(new_n633), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n701), .A2(new_n587), .A3(new_n697), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n679), .A2(new_n687), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n702), .A2(new_n672), .A3(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(KEYINPUT101), .B(G125), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G27));
  INV_X1    g520(.A(KEYINPUT103), .ZN(new_n707));
  AOI21_X1  g521(.A(KEYINPUT32), .B1(new_n289), .B2(new_n290), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n282), .A2(new_n296), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n707), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n289), .A2(new_n293), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n711), .B(KEYINPUT103), .C1(KEYINPUT32), .C2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n710), .A2(new_n313), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n580), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n399), .A2(new_n315), .A3(new_n400), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(KEYINPUT102), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT102), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n399), .A2(new_n718), .A3(new_n315), .A4(new_n400), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n717), .A2(new_n672), .A3(new_n441), .A4(new_n719), .ZN(new_n720));
  OAI21_X1  g534(.A(KEYINPUT42), .B1(new_n715), .B2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n717), .A2(new_n441), .A3(new_n719), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n672), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(KEYINPUT42), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n723), .A2(new_n725), .A3(new_n314), .A4(new_n580), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n721), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n218), .ZN(G33));
  XNOR2_X1  g542(.A(new_n643), .B(KEYINPUT104), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n723), .A2(new_n729), .A3(new_n314), .A4(new_n580), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G134), .ZN(G36));
  OR2_X1    g545(.A1(new_n439), .A2(KEYINPUT45), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n439), .A2(KEYINPUT45), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(G469), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(G469), .A2(G902), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT105), .ZN(new_n738));
  OR3_X1    g552(.A1(new_n737), .A2(new_n738), .A3(KEYINPUT46), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n738), .B1(new_n737), .B2(KEYINPUT46), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n737), .A2(KEYINPUT46), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n739), .A2(new_n436), .A3(new_n740), .A4(new_n741), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n742), .A2(new_n678), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n667), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n661), .A2(new_n605), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(KEYINPUT43), .ZN(new_n746));
  OR3_X1    g560(.A1(new_n746), .A2(new_n588), .A3(new_n701), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT44), .ZN(new_n748));
  OR2_X1    g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n717), .A2(new_n719), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n747), .A2(new_n748), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n744), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n216), .ZN(G39));
  AND2_X1   g568(.A1(new_n743), .A2(KEYINPUT47), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n743), .A2(KEYINPUT47), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n314), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n758), .A2(new_n579), .A3(new_n672), .A4(new_n750), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(KEYINPUT106), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G140), .ZN(G42));
  INV_X1    g576(.A(new_n479), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n746), .A2(new_n763), .ZN(new_n764));
  XOR2_X1   g578(.A(new_n764), .B(KEYINPUT115), .Z(new_n765));
  INV_X1    g579(.A(new_n698), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI211_X1 g581(.A(new_n478), .B(G953), .C1(new_n767), .C2(new_n703), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n750), .A2(new_n680), .ZN(new_n769));
  NOR4_X1   g583(.A1(new_n660), .A2(new_n579), .A3(new_n763), .A4(new_n769), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n605), .A2(new_n536), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n765), .A2(new_n769), .ZN(new_n773));
  INV_X1    g587(.A(new_n715), .ZN(new_n774));
  XNOR2_X1  g588(.A(KEYINPUT117), .B(KEYINPUT48), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n775), .B1(new_n773), .B2(new_n774), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n768), .B(new_n772), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n778), .A2(KEYINPUT118), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(KEYINPUT118), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n666), .A2(new_n315), .A3(new_n679), .ZN(new_n782));
  XOR2_X1   g596(.A(new_n782), .B(KEYINPUT116), .Z(new_n783));
  NAND2_X1  g597(.A1(new_n767), .A2(new_n783), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n784), .A2(KEYINPUT50), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n773), .A2(new_n702), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n784), .A2(KEYINPUT50), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n605), .A2(new_n536), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n770), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n785), .A2(new_n786), .A3(new_n787), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n767), .A2(new_n750), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n755), .A2(new_n756), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n677), .A2(new_n405), .A3(new_n436), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n781), .B1(new_n790), .B2(new_n794), .ZN(new_n795));
  AOI22_X1  g609(.A1(new_n779), .A2(new_n780), .B1(new_n795), .B2(KEYINPUT51), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n795), .A2(KEYINPUT51), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT108), .ZN(new_n799));
  AND4_X1   g613(.A1(new_n314), .A2(new_n723), .A3(new_n729), .A4(new_n580), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n662), .A2(new_n519), .A3(new_n642), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n614), .A2(new_n618), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n701), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n803), .B1(new_n645), .B2(new_n648), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n587), .A2(new_n697), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n634), .A3(new_n672), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n722), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n799), .B1(new_n800), .B2(new_n807), .ZN(new_n808));
  AOI22_X1  g622(.A1(new_n314), .A2(new_n803), .B1(new_n672), .B2(new_n702), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n730), .B(KEYINPUT108), .C1(new_n809), .C2(new_n722), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  AOI22_X1  g625(.A1(new_n314), .A2(new_n688), .B1(new_n694), .B2(new_n698), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n684), .A2(new_n812), .A3(new_n681), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n727), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n662), .A2(new_n536), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n771), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n596), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n817), .A2(new_n588), .A3(new_n584), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n582), .A2(new_n635), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT107), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT107), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n582), .A2(new_n635), .A3(new_n818), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n811), .A2(new_n814), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(KEYINPUT109), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT109), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n811), .A2(new_n814), .A3(new_n823), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n680), .A2(new_n401), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n806), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n648), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n724), .B1(new_n830), .B2(new_n292), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n829), .B1(new_n639), .B2(new_n831), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n441), .A2(new_n665), .A3(new_n642), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n659), .A2(new_n663), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n653), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT112), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT112), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n653), .A2(new_n832), .A3(new_n838), .A4(new_n834), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n836), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n837), .B1(new_n836), .B2(new_n839), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n825), .B(new_n827), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n813), .A2(KEYINPUT113), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT113), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n684), .A2(new_n812), .A3(new_n681), .A4(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n721), .A2(KEYINPUT53), .A3(new_n726), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n849), .A2(new_n811), .A3(new_n823), .A4(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n836), .A2(new_n837), .A3(new_n839), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT111), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n853), .B1(new_n835), .B2(new_n837), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n673), .A2(new_n704), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n855), .B1(new_n652), .B2(new_n650), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n856), .A2(KEYINPUT111), .A3(KEYINPUT52), .A4(new_n834), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n851), .B1(new_n852), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n844), .A2(new_n845), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n842), .A2(KEYINPUT53), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n825), .A2(KEYINPUT110), .A3(new_n827), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n858), .A2(new_n852), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(new_n843), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT110), .B1(new_n825), .B2(new_n827), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n862), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n861), .B1(new_n867), .B2(new_n845), .ZN(new_n868));
  OAI22_X1  g682(.A1(new_n798), .A2(new_n868), .B1(G952), .B2(G953), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n677), .A2(new_n436), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n870), .A2(KEYINPUT49), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(KEYINPUT49), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n745), .A2(new_n405), .A3(new_n316), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n872), .A2(new_n580), .A3(new_n873), .ZN(new_n874));
  OR4_X1    g688(.A1(new_n660), .A2(new_n666), .A3(new_n871), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n869), .A2(new_n875), .ZN(G75));
  NAND2_X1  g690(.A1(new_n844), .A2(new_n860), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(G210), .A3(G902), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT56), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n351), .B(new_n364), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT55), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n880), .A2(new_n882), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n265), .A2(G952), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(G51));
  INV_X1    g700(.A(new_n877), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n734), .B(KEYINPUT120), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n887), .A2(new_n308), .A3(new_n888), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n735), .B(KEYINPUT57), .Z(new_n890));
  AOI21_X1  g704(.A(new_n845), .B1(new_n844), .B2(new_n860), .ZN(new_n891));
  AOI211_X1 g705(.A(KEYINPUT54), .B(new_n859), .C1(new_n842), .C2(new_n843), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n676), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT119), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n889), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n893), .A2(KEYINPUT119), .A3(new_n894), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n885), .B1(new_n897), .B2(new_n898), .ZN(G54));
  NOR2_X1   g713(.A1(new_n887), .A2(new_n308), .ZN(new_n900));
  AND2_X1   g714(.A1(KEYINPUT58), .A2(G475), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n900), .A2(new_n531), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n531), .B1(new_n900), .B2(new_n901), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n902), .A2(new_n903), .A3(new_n885), .ZN(G60));
  XOR2_X1   g718(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n905));
  NOR2_X1   g719(.A1(new_n442), .A2(new_n308), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n905), .B(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n868), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n603), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n877), .A2(KEYINPUT54), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n861), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n602), .A2(new_n907), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n885), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n909), .A2(new_n913), .A3(KEYINPUT122), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT122), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n602), .B1(new_n868), .B2(new_n907), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n912), .B1(new_n891), .B2(new_n892), .ZN(new_n917));
  INV_X1    g731(.A(new_n885), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n915), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n914), .A2(new_n920), .ZN(G63));
  NAND2_X1  g735(.A1(new_n568), .A2(new_n569), .ZN(new_n922));
  XNOR2_X1  g736(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n444), .A2(new_n308), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n922), .B1(new_n887), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n877), .A2(new_n632), .A3(new_n925), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n927), .A2(new_n918), .A3(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT61), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(G66));
  INV_X1    g745(.A(G224), .ZN(new_n932));
  OAI21_X1  g746(.A(G953), .B1(new_n481), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n813), .B1(new_n820), .B2(new_n822), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n933), .B1(new_n934), .B2(G953), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n351), .B1(G898), .B2(new_n265), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT124), .Z(new_n937));
  XNOR2_X1  g751(.A(new_n935), .B(new_n937), .ZN(G69));
  NAND2_X1  g752(.A1(new_n274), .A2(new_n275), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(new_n524), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n727), .B1(new_n757), .B2(new_n760), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n744), .A2(new_n692), .A3(new_n715), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n942), .A2(new_n753), .A3(new_n800), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n941), .A2(new_n856), .A3(new_n943), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n944), .A2(new_n265), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n265), .A2(G900), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT125), .Z(new_n947));
  OAI21_X1  g761(.A(new_n940), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n940), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n816), .A2(new_n668), .ZN(new_n950));
  AND4_X1   g764(.A1(new_n314), .A2(new_n950), .A3(new_n580), .A4(new_n750), .ZN(new_n951));
  AOI211_X1 g765(.A(new_n753), .B(new_n951), .C1(new_n757), .C2(new_n760), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n670), .A2(new_n856), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n952), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n949), .B1(new_n956), .B2(G953), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n948), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n265), .B1(G227), .B2(G900), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(G72));
  XNOR2_X1  g774(.A(new_n309), .B(KEYINPUT127), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n269), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n952), .A2(new_n934), .A3(new_n954), .A4(new_n955), .ZN(new_n963));
  NAND2_X1  g777(.A1(G472), .A2(G902), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT63), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT126), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n962), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n309), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n656), .B1(new_n270), .B2(new_n968), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n867), .A2(new_n965), .A3(new_n969), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n941), .A2(new_n934), .A3(new_n943), .A4(new_n856), .ZN(new_n971));
  AOI211_X1 g785(.A(new_n269), .B(new_n961), .C1(new_n971), .C2(new_n966), .ZN(new_n972));
  NOR4_X1   g786(.A1(new_n967), .A2(new_n970), .A3(new_n972), .A4(new_n885), .ZN(G57));
endmodule


