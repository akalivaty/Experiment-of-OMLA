//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n827, new_n828,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(G8gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT14), .ZN(new_n208));
  INV_X1    g007(.A(G29gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n211));
  AOI21_X1  g010(.A(G36gat), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G36gat), .ZN(new_n213));
  NOR3_X1   g012(.A1(new_n208), .A2(new_n213), .A3(G29gat), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT15), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n214), .ZN(new_n216));
  INV_X1    g015(.A(new_n211), .ZN(new_n217));
  NOR2_X1   g016(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n213), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT15), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n216), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G43gat), .B(G50gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n215), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n222), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n224), .B(KEYINPUT15), .C1(new_n212), .C2(new_n214), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(KEYINPUT17), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT17), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n228), .B1(new_n223), .B2(new_n225), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n207), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G229gat), .A2(G233gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n206), .A2(new_n226), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT18), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT90), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n230), .A2(KEYINPUT18), .A3(new_n231), .A4(new_n232), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n206), .B(new_n226), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n231), .B(KEYINPUT13), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G113gat), .B(G141gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G169gat), .B(G197gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(KEYINPUT12), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n233), .A2(KEYINPUT90), .A3(new_n234), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n237), .A2(new_n242), .A3(new_n248), .A4(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT89), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n233), .A2(KEYINPUT89), .A3(new_n234), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n252), .A2(new_n242), .A3(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n250), .B1(new_n254), .B2(new_n248), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n257));
  XNOR2_X1  g056(.A(G113gat), .B(G120gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n258), .A2(KEYINPUT1), .ZN(new_n259));
  XNOR2_X1  g058(.A(G127gat), .B(G134gat), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n257), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n260), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n262), .B(KEYINPUT68), .C1(KEYINPUT1), .C2(new_n258), .ZN(new_n263));
  INV_X1    g062(.A(new_n258), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(new_n260), .A3(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n261), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268));
  INV_X1    g067(.A(G155gat), .ZN(new_n269));
  INV_X1    g068(.A(G162gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n268), .B1(new_n271), .B2(KEYINPUT2), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT78), .ZN(new_n273));
  INV_X1    g072(.A(G141gat), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n273), .B1(new_n274), .B2(G148gat), .ZN(new_n275));
  INV_X1    g074(.A(G148gat), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n275), .B1(G141gat), .B2(new_n276), .ZN(new_n277));
  NOR3_X1   g076(.A1(new_n273), .A2(new_n274), .A3(G148gat), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n272), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G141gat), .B(G148gat), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n268), .B(new_n271), .C1(new_n280), .C2(KEYINPUT2), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT4), .B1(new_n267), .B2(new_n282), .ZN(new_n283));
  OR2_X1    g082(.A1(new_n283), .A2(KEYINPUT81), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n261), .A2(new_n263), .A3(new_n266), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT4), .ZN(new_n286));
  INV_X1    g085(.A(new_n282), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(KEYINPUT81), .A3(new_n283), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n267), .A2(KEYINPUT79), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT79), .ZN(new_n291));
  NAND4_X1  g090(.A1(new_n261), .A2(new_n291), .A3(new_n263), .A4(new_n266), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n282), .A2(KEYINPUT3), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT3), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n279), .A2(new_n294), .A3(new_n281), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n290), .A2(new_n292), .A3(new_n293), .A4(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n284), .A2(new_n289), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(G225gat), .A2(G233gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n299), .A2(KEYINPUT5), .ZN(new_n300));
  OR2_X1    g099(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n290), .A2(KEYINPUT80), .A3(new_n292), .A4(new_n282), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n290), .A2(new_n292), .A3(new_n282), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT80), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n298), .B1(new_n304), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n288), .A2(new_n283), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n309), .A2(new_n298), .A3(new_n296), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT5), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n301), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G1gat), .B(G29gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n313), .B(KEYINPUT0), .ZN(new_n314));
  XNOR2_X1  g113(.A(G57gat), .B(G85gat), .ZN(new_n315));
  XOR2_X1   g114(.A(new_n314), .B(new_n315), .Z(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT6), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n301), .B(new_n316), .C1(new_n308), .C2(new_n311), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n312), .A2(KEYINPUT6), .A3(new_n317), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  XOR2_X1   g122(.A(G8gat), .B(G36gat), .Z(new_n324));
  XNOR2_X1  g123(.A(new_n324), .B(KEYINPUT75), .ZN(new_n325));
  XNOR2_X1  g124(.A(G64gat), .B(G92gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT74), .ZN(new_n328));
  XNOR2_X1  g127(.A(G197gat), .B(G204gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT22), .ZN(new_n330));
  INV_X1    g129(.A(G211gat), .ZN(new_n331));
  INV_X1    g130(.A(G218gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G211gat), .B(G218gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  AND2_X1   g136(.A1(new_n329), .A2(new_n333), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT73), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n335), .B1(new_n334), .B2(KEYINPUT73), .ZN(new_n341));
  AOI211_X1 g140(.A(new_n328), .B(new_n337), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n341), .A3(new_n328), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(KEYINPUT27), .B(G183gat), .Z(new_n346));
  OAI21_X1  g145(.A(KEYINPUT66), .B1(new_n346), .B2(G190gat), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G169gat), .A2(G176gat), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT26), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(G169gat), .ZN(new_n353));
  INV_X1    g152(.A(G176gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT67), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n352), .A2(KEYINPUT67), .A3(new_n355), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n358), .B(new_n359), .C1(KEYINPUT26), .C2(new_n355), .ZN(new_n360));
  OAI211_X1 g159(.A(KEYINPUT66), .B(KEYINPUT28), .C1(new_n346), .C2(G190gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(G183gat), .A2(G190gat), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n349), .A2(new_n360), .A3(new_n361), .A4(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT23), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n355), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n353), .A2(new_n354), .A3(KEYINPUT23), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n365), .A2(new_n350), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n370));
  MUX2_X1   g169(.A(KEYINPUT65), .B(new_n369), .S(new_n370), .Z(new_n371));
  AND2_X1   g170(.A1(new_n362), .A2(KEYINPUT64), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n362), .A2(KEYINPUT64), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n372), .A2(new_n373), .A3(KEYINPUT24), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n368), .B1(new_n371), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT25), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n362), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n378), .A2(new_n370), .ZN(new_n379));
  NOR3_X1   g178(.A1(new_n379), .A2(new_n367), .A3(KEYINPUT25), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n363), .A2(new_n376), .A3(new_n381), .ZN(new_n382));
  AND2_X1   g181(.A1(G226gat), .A2(G233gat), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT29), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n383), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n345), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n345), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n382), .A2(new_n383), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n380), .B1(KEYINPUT25), .B2(new_n375), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT29), .B1(new_n390), .B2(new_n363), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n388), .B(new_n389), .C1(new_n383), .C2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n327), .B1(new_n387), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT30), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n387), .A2(new_n327), .A3(new_n392), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n387), .A2(new_n392), .ZN(new_n397));
  INV_X1    g196(.A(new_n327), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  XOR2_X1   g198(.A(KEYINPUT76), .B(KEYINPUT30), .Z(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n399), .A2(KEYINPUT77), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT77), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n403), .B1(new_n393), .B2(new_n400), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n396), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n323), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT85), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT83), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n295), .A2(new_n385), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n409), .B1(new_n342), .B2(new_n344), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n338), .A2(new_n335), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n385), .B1(new_n411), .B2(new_n337), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n294), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n282), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(G228gat), .A2(G233gat), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n408), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n338), .A2(new_n335), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n336), .B1(new_n338), .B2(new_n339), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n334), .A2(KEYINPUT73), .ZN(new_n420));
  OAI211_X1 g219(.A(KEYINPUT74), .B(new_n418), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  AOI22_X1  g220(.A1(new_n421), .A2(new_n343), .B1(new_n385), .B2(new_n295), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n287), .B1(new_n412), .B2(new_n294), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n408), .B(new_n416), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n417), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n410), .A2(G228gat), .A3(G233gat), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n421), .A2(new_n385), .A3(new_n343), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT84), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n421), .A2(KEYINPUT84), .A3(new_n385), .A4(new_n343), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(new_n294), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n427), .B1(new_n432), .B2(new_n282), .ZN(new_n433));
  NOR3_X1   g232(.A1(new_n426), .A2(new_n433), .A3(G22gat), .ZN(new_n434));
  INV_X1    g233(.A(G22gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n432), .A2(new_n282), .ZN(new_n436));
  INV_X1    g235(.A(new_n427), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n416), .B1(new_n422), .B2(new_n423), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT83), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n424), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n435), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n407), .B1(new_n434), .B2(new_n442), .ZN(new_n443));
  XOR2_X1   g242(.A(G78gat), .B(G106gat), .Z(new_n444));
  XNOR2_X1  g243(.A(new_n444), .B(G50gat), .ZN(new_n445));
  XOR2_X1   g244(.A(KEYINPUT82), .B(KEYINPUT31), .Z(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(G22gat), .B1(new_n426), .B2(new_n433), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n438), .A2(new_n435), .A3(new_n441), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(KEYINPUT85), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n443), .A2(new_n448), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT86), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n449), .A2(new_n450), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n454), .A2(new_n407), .A3(new_n447), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n452), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n453), .B1(new_n452), .B2(new_n455), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n406), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n297), .A2(new_n299), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n304), .A2(new_n298), .A3(new_n307), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(new_n460), .A3(KEYINPUT39), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT39), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n297), .A2(new_n462), .A3(new_n299), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n461), .A2(new_n316), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT40), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n461), .A2(KEYINPUT40), .A3(new_n316), .A4(new_n463), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n318), .A3(new_n467), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n452), .B(new_n455), .C1(new_n405), .C2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT37), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n387), .A2(new_n470), .A3(new_n392), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n470), .B1(new_n387), .B2(new_n392), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n327), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n393), .B1(new_n473), .B2(KEYINPUT38), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT38), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n475), .B(new_n327), .C1(new_n471), .C2(new_n472), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n474), .A2(new_n321), .A3(new_n322), .A4(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT87), .B1(new_n469), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n382), .A2(new_n285), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n390), .A2(new_n267), .A3(new_n363), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(G227gat), .A2(G233gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT71), .B1(new_n484), .B2(KEYINPUT34), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT71), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT34), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n482), .A2(new_n486), .A3(new_n487), .A4(new_n483), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n484), .A2(KEYINPUT34), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n485), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n480), .A2(G227gat), .A3(G233gat), .A4(new_n481), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT32), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT70), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n492), .A2(KEYINPUT70), .A3(KEYINPUT32), .ZN(new_n496));
  XNOR2_X1  g295(.A(G15gat), .B(G43gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(G71gat), .B(G99gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT33), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n499), .B1(new_n492), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n495), .A2(new_n496), .A3(new_n501), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n492), .B(KEYINPUT32), .C1(new_n500), .C2(new_n499), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n491), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n503), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n490), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n506), .A3(KEYINPUT72), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT36), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT72), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n505), .A2(new_n509), .A3(new_n490), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n507), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n504), .A2(new_n506), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT36), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  OR2_X1    g313(.A1(new_n405), .A2(new_n468), .ZN(new_n515));
  AOI211_X1 g314(.A(KEYINPUT85), .B(new_n448), .C1(new_n449), .C2(new_n450), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n447), .B1(new_n454), .B2(new_n407), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n516), .B1(new_n517), .B2(new_n451), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT87), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n515), .A2(new_n518), .A3(new_n519), .A4(new_n477), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n458), .A2(new_n479), .A3(new_n514), .A4(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n406), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n510), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT35), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n522), .A2(new_n523), .A3(new_n524), .A4(new_n518), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n512), .A2(new_n455), .A3(new_n452), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT35), .B1(new_n526), .B2(new_n406), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n256), .B1(new_n521), .B2(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(G99gat), .B(G106gat), .Z(new_n530));
  NAND2_X1  g329(.A1(G99gat), .A2(G106gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT8), .ZN(new_n532));
  OR2_X1    g331(.A1(G85gat), .A2(G92gat), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n532), .A2(KEYINPUT95), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT95), .B1(new_n532), .B2(new_n533), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT94), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OR2_X1    g338(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n540));
  NAND2_X1  g339(.A1(G85gat), .A2(G92gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(KEYINPUT93), .A2(KEYINPUT94), .A3(KEYINPUT7), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  AND3_X1   g342(.A1(KEYINPUT93), .A2(KEYINPUT94), .A3(KEYINPUT7), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT94), .B1(KEYINPUT93), .B2(KEYINPUT7), .ZN(new_n545));
  AND2_X1   g344(.A1(G85gat), .A2(G92gat), .ZN(new_n546));
  NOR2_X1   g345(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n547));
  OAI22_X1  g346(.A1(new_n544), .A2(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n530), .B1(new_n536), .B2(new_n549), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n543), .A2(new_n548), .ZN(new_n551));
  INV_X1    g350(.A(new_n530), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT95), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT8), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n554), .B1(G99gat), .B2(G106gat), .ZN(new_n555));
  NOR2_X1   g354(.A1(G85gat), .A2(G92gat), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n553), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n532), .A2(new_n533), .A3(KEYINPUT95), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n551), .A2(new_n552), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n550), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n561), .B1(new_n227), .B2(new_n229), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT96), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT96), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n564), .B(new_n561), .C1(new_n227), .C2(new_n229), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n226), .A2(new_n560), .A3(new_n550), .ZN(new_n567));
  NAND2_X1  g366(.A1(G232gat), .A2(G233gat), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT41), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(G190gat), .B(G218gat), .Z(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n569), .A2(KEYINPUT41), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n576), .B(KEYINPUT92), .Z(new_n577));
  XNOR2_X1  g376(.A(G134gat), .B(G162gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n574), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n566), .A2(new_n580), .A3(new_n572), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n575), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n579), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n580), .B1(new_n566), .B2(new_n572), .ZN(new_n584));
  AOI211_X1 g383(.A(new_n574), .B(new_n571), .C1(new_n563), .C2(new_n565), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G57gat), .B(G64gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(G71gat), .A2(G78gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(G71gat), .A2(G78gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT9), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n590), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n592), .B(new_n591), .C1(new_n589), .C2(new_n594), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT21), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G127gat), .B(G155gat), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n600), .B(new_n601), .Z(new_n602));
  AND2_X1   g401(.A1(new_n596), .A2(new_n597), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n206), .B1(KEYINPUT21), .B2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n602), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G231gat), .A2(G233gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT91), .ZN(new_n607));
  XOR2_X1   g406(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G183gat), .B(G211gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n605), .B(new_n611), .Z(new_n612));
  NAND2_X1  g411(.A1(new_n588), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G120gat), .B(G148gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(G176gat), .B(G204gat), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n614), .B(new_n615), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G230gat), .A2(G233gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n618), .B(KEYINPUT97), .Z(new_n619));
  NOR3_X1   g418(.A1(new_n536), .A2(new_n549), .A3(new_n530), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n552), .B1(new_n551), .B2(new_n559), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n598), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT10), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n550), .A2(new_n560), .A3(new_n603), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n550), .A2(new_n560), .A3(new_n603), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT10), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n619), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n619), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n629), .B1(new_n622), .B2(new_n624), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n617), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n631), .B(KEYINPUT99), .Z(new_n632));
  AOI21_X1  g431(.A(new_n603), .B1(new_n550), .B2(new_n560), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n626), .A2(new_n633), .A3(KEYINPUT10), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n624), .A2(new_n623), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n629), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(KEYINPUT98), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT98), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n628), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n630), .A2(new_n617), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n637), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n632), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n613), .A2(new_n642), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n529), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n323), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT100), .B(G1gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(G1324gat));
  INV_X1    g447(.A(new_n644), .ZN(new_n649));
  OAI21_X1  g448(.A(G8gat), .B1(new_n649), .B2(new_n405), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n650), .A2(KEYINPUT101), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n402), .A2(new_n404), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n652), .A2(new_n395), .A3(new_n394), .ZN(new_n653));
  XOR2_X1   g452(.A(KEYINPUT16), .B(G8gat), .Z(new_n654));
  NAND3_X1  g453(.A1(new_n644), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT42), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n650), .A2(KEYINPUT101), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n651), .A2(new_n656), .A3(new_n657), .ZN(G1325gat));
  OAI21_X1  g457(.A(G15gat), .B1(new_n649), .B2(new_n514), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n529), .A2(new_n523), .ZN(new_n660));
  INV_X1    g459(.A(G15gat), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n660), .A2(new_n661), .A3(new_n643), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(new_n662), .ZN(G1326gat));
  OR2_X1    g462(.A1(new_n456), .A2(new_n457), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n529), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n643), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n666), .A2(KEYINPUT102), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(KEYINPUT102), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT43), .B(G22gat), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n669), .B1(new_n667), .B2(new_n668), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(G1327gat));
  NAND2_X1  g471(.A1(new_n521), .A2(new_n528), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n642), .A2(new_n612), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(new_n256), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n673), .A2(new_n587), .A3(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n677), .A2(new_n209), .A3(new_n645), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT45), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n680), .B1(new_n673), .B2(new_n587), .ZN(new_n681));
  AND3_X1   g480(.A1(new_n582), .A2(new_n586), .A3(KEYINPUT104), .ZN(new_n682));
  AOI21_X1  g481(.A(KEYINPUT104), .B1(new_n582), .B2(new_n586), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  AOI211_X1 g484(.A(KEYINPUT44), .B(new_n685), .C1(new_n521), .C2(new_n528), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n676), .B(KEYINPUT103), .Z(new_n688));
  AND2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n645), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n679), .B1(new_n691), .B2(new_n209), .ZN(G1328gat));
  NAND3_X1  g491(.A1(new_n677), .A2(new_n213), .A3(new_n653), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n693), .B(KEYINPUT46), .Z(new_n694));
  NAND2_X1  g493(.A1(new_n689), .A2(new_n653), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n694), .B1(new_n696), .B2(new_n213), .ZN(G1329gat));
  INV_X1    g496(.A(G43gat), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n675), .A2(new_n588), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n660), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n514), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n701), .B(new_n688), .C1(new_n681), .C2(new_n686), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n700), .B1(new_n703), .B2(new_n698), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT47), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1330gat));
  INV_X1    g505(.A(new_n518), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n707), .B(new_n688), .C1(new_n681), .C2(new_n686), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(G50gat), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT105), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT48), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n675), .A2(G50gat), .A3(new_n588), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n711), .B1(new_n665), .B2(new_n712), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n709), .A2(new_n710), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n710), .B1(new_n709), .B2(new_n713), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n687), .A2(new_n664), .A3(new_n688), .ZN(new_n716));
  AOI22_X1  g515(.A1(new_n716), .A2(G50gat), .B1(new_n665), .B2(new_n712), .ZN(new_n717));
  OAI22_X1  g516(.A1(new_n714), .A2(new_n715), .B1(new_n717), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g517(.A(new_n642), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n613), .A2(new_n719), .A3(new_n255), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n673), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n645), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT106), .B(G57gat), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1332gat));
  AOI21_X1  g523(.A(new_n405), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT107), .ZN(new_n727));
  NOR2_X1   g526(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1333gat));
  NAND2_X1  g528(.A1(new_n721), .A2(new_n701), .ZN(new_n730));
  AOI21_X1  g529(.A(G71gat), .B1(new_n507), .B2(new_n510), .ZN(new_n731));
  AOI22_X1  g530(.A1(new_n730), .A2(G71gat), .B1(new_n721), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g532(.A1(new_n721), .A2(new_n664), .ZN(new_n734));
  XNOR2_X1  g533(.A(KEYINPUT108), .B(G78gat), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1335gat));
  NOR2_X1   g535(.A1(new_n255), .A2(new_n612), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n673), .A2(new_n587), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT51), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(G85gat), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n740), .A2(new_n741), .A3(new_n645), .A4(new_n642), .ZN(new_n742));
  INV_X1    g541(.A(new_n737), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n719), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n687), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n645), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n742), .B1(new_n747), .B2(new_n741), .ZN(G1336gat));
  AOI211_X1 g547(.A(new_n588), .B(new_n743), .C1(new_n521), .C2(new_n528), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n739), .B1(new_n749), .B2(KEYINPUT109), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n738), .A2(new_n751), .A3(KEYINPUT51), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n719), .A2(new_n405), .A3(G92gat), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n750), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n750), .A2(KEYINPUT110), .A3(new_n752), .A4(new_n753), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n653), .B(new_n744), .C1(new_n681), .C2(new_n686), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(G92gat), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n756), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT52), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT52), .B1(new_n740), .B2(new_n753), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n759), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(G1337gat));
  INV_X1    g563(.A(G99gat), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n740), .A2(new_n765), .A3(new_n523), .A4(new_n642), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n745), .A2(new_n701), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n766), .B1(new_n768), .B2(new_n765), .ZN(G1338gat));
  NOR3_X1   g568(.A1(new_n518), .A2(G106gat), .A3(new_n719), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT53), .B1(new_n740), .B2(new_n770), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n707), .B(new_n744), .C1(new_n681), .C2(new_n686), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT111), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(G106gat), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n772), .A2(KEYINPUT111), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n771), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n664), .B(new_n744), .C1(new_n681), .C2(new_n686), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n777), .A2(G106gat), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n750), .A2(new_n752), .A3(new_n770), .ZN(new_n779));
  OAI21_X1  g578(.A(KEYINPUT53), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n776), .A2(new_n780), .ZN(G1339gat));
  INV_X1    g580(.A(new_n612), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n625), .A2(new_n619), .A3(new_n627), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n783), .A2(KEYINPUT54), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n637), .A2(new_n784), .A3(new_n639), .ZN(new_n785));
  AOI211_X1 g584(.A(KEYINPUT54), .B(new_n619), .C1(new_n625), .C2(new_n627), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n786), .A2(KEYINPUT112), .A3(new_n616), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n789), .B(new_n629), .C1(new_n634), .C2(new_n635), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n788), .B1(new_n790), .B2(new_n617), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n785), .B(KEYINPUT55), .C1(new_n787), .C2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n641), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT113), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n792), .A2(KEYINPUT113), .A3(new_n641), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT112), .B1(new_n786), .B2(new_n616), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n790), .A2(new_n788), .A3(new_n617), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT55), .B1(new_n799), .B2(new_n785), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n795), .A2(new_n255), .A3(new_n796), .A4(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n239), .A2(new_n240), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n231), .B1(new_n230), .B2(new_n232), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n247), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n642), .A2(new_n250), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n684), .B1(new_n802), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n800), .B1(new_n793), .B2(new_n794), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n809));
  AND3_X1   g608(.A1(new_n250), .A2(new_n809), .A3(new_n805), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n809), .B1(new_n250), .B2(new_n805), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AND4_X1   g611(.A1(new_n684), .A2(new_n808), .A3(new_n812), .A4(new_n796), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n782), .B1(new_n807), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n643), .A2(new_n256), .ZN(new_n815));
  AOI211_X1 g614(.A(new_n323), .B(new_n526), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n816), .A2(new_n405), .ZN(new_n817));
  AOI21_X1  g616(.A(G113gat), .B1(new_n817), .B2(new_n255), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n664), .B1(new_n814), .B2(new_n815), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n819), .A2(new_n645), .A3(new_n405), .A4(new_n523), .ZN(new_n820));
  XOR2_X1   g619(.A(new_n820), .B(KEYINPUT115), .Z(new_n821));
  AND2_X1   g620(.A1(new_n255), .A2(G113gat), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n818), .B1(new_n821), .B2(new_n822), .ZN(G1340gat));
  AOI21_X1  g622(.A(G120gat), .B1(new_n817), .B2(new_n642), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n642), .A2(G120gat), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n824), .B1(new_n821), .B2(new_n825), .ZN(G1341gat));
  INV_X1    g625(.A(new_n821), .ZN(new_n827));
  OAI21_X1  g626(.A(G127gat), .B1(new_n827), .B2(new_n782), .ZN(new_n828));
  INV_X1    g627(.A(G127gat), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n817), .A2(new_n829), .A3(new_n612), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(G1342gat));
  OAI21_X1  g630(.A(G134gat), .B1(new_n827), .B2(new_n588), .ZN(new_n832));
  INV_X1    g631(.A(G134gat), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n653), .A2(new_n588), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n816), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  XOR2_X1   g634(.A(new_n835), .B(KEYINPUT56), .Z(new_n836));
  NAND2_X1  g635(.A1(new_n832), .A2(new_n836), .ZN(G1343gat));
  NOR3_X1   g636(.A1(new_n701), .A2(new_n323), .A3(new_n653), .ZN(new_n838));
  INV_X1    g637(.A(new_n813), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n801), .A2(new_n255), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n806), .B1(new_n840), .B2(new_n793), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n588), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n612), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n815), .ZN(new_n844));
  OAI211_X1 g643(.A(KEYINPUT57), .B(new_n664), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n814), .A2(new_n815), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT57), .B1(new_n846), .B2(new_n707), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n845), .B1(new_n847), .B2(KEYINPUT116), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n849));
  AOI211_X1 g648(.A(new_n849), .B(KEYINPUT57), .C1(new_n846), .C2(new_n707), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n255), .B(new_n838), .C1(new_n848), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(G141gat), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n846), .A2(new_n645), .A3(new_n707), .A4(new_n514), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n853), .A2(new_n653), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n274), .A3(new_n255), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT58), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT58), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n852), .A2(new_n858), .A3(new_n855), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(G1344gat));
  NOR2_X1   g659(.A1(new_n276), .A2(KEYINPUT59), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n838), .B1(new_n848), .B2(new_n850), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n861), .B1(new_n862), .B2(new_n719), .ZN(new_n863));
  XOR2_X1   g662(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n864));
  NAND2_X1  g663(.A1(new_n846), .A2(new_n707), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(KEYINPUT57), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n808), .A2(new_n587), .A3(new_n812), .A4(new_n796), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n612), .B1(new_n842), .B2(new_n868), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n867), .B(new_n664), .C1(new_n869), .C2(new_n844), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n838), .A2(new_n642), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n276), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n863), .B1(new_n864), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n854), .A2(new_n276), .A3(new_n642), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(G1345gat));
  OAI211_X1 g675(.A(new_n612), .B(new_n838), .C1(new_n848), .C2(new_n850), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(G155gat), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n854), .A2(new_n269), .A3(new_n612), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n878), .A2(KEYINPUT118), .A3(new_n879), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1346gat));
  OAI21_X1  g683(.A(G162gat), .B1(new_n862), .B2(new_n685), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n834), .A2(new_n270), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n885), .B1(new_n853), .B2(new_n886), .ZN(G1347gat));
  AOI21_X1  g686(.A(new_n645), .B1(new_n814), .B2(new_n815), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n526), .A2(new_n405), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(G169gat), .B1(new_n890), .B2(new_n255), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n645), .A2(new_n405), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n523), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT119), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n819), .A2(new_n894), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n895), .A2(new_n353), .A3(new_n256), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n891), .A2(new_n896), .ZN(G1348gat));
  NAND3_X1  g696(.A1(new_n890), .A2(new_n354), .A3(new_n642), .ZN(new_n898));
  OAI21_X1  g697(.A(G176gat), .B1(new_n895), .B2(new_n719), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1349gat));
  NOR2_X1   g699(.A1(new_n782), .A2(new_n346), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n819), .A2(new_n612), .A3(new_n894), .ZN(new_n902));
  AOI22_X1  g701(.A1(new_n890), .A2(new_n901), .B1(new_n902), .B2(G183gat), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT60), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n905), .A2(KEYINPUT120), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n905), .A2(KEYINPUT120), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT121), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n908), .B1(new_n903), .B2(new_n904), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n903), .A2(new_n908), .A3(new_n904), .ZN(new_n910));
  OAI22_X1  g709(.A1(new_n906), .A2(new_n907), .B1(new_n909), .B2(new_n910), .ZN(G1350gat));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912));
  OAI21_X1  g711(.A(G190gat), .B1(new_n895), .B2(new_n588), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n914), .A2(KEYINPUT123), .A3(new_n915), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n913), .A2(KEYINPUT122), .A3(KEYINPUT61), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n919), .B1(new_n913), .B2(KEYINPUT61), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n916), .A2(new_n917), .A3(new_n918), .A4(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(G190gat), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n890), .A2(new_n922), .A3(new_n684), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(G1351gat));
  NAND2_X1  g723(.A1(new_n871), .A2(KEYINPUT126), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n514), .A2(new_n892), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n866), .A2(new_n870), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n925), .A2(new_n926), .A3(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(G197gat), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n930), .A2(new_n931), .A3(new_n256), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n514), .A2(new_n653), .A3(new_n707), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT124), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(new_n888), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT125), .ZN(new_n936));
  AOI21_X1  g735(.A(G197gat), .B1(new_n936), .B2(new_n255), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n932), .A2(new_n937), .ZN(G1352gat));
  OAI21_X1  g737(.A(G204gat), .B1(new_n930), .B2(new_n719), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n935), .A2(G204gat), .A3(new_n719), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT62), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(G1353gat));
  NAND3_X1  g741(.A1(new_n936), .A2(new_n331), .A3(new_n612), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n871), .A2(new_n612), .A3(new_n926), .ZN(new_n944));
  AND4_X1   g743(.A1(KEYINPUT127), .A2(new_n944), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n945));
  OAI21_X1  g744(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  AOI22_X1  g746(.A1(new_n944), .A2(new_n947), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n943), .B1(new_n945), .B2(new_n948), .ZN(G1354gat));
  NOR3_X1   g748(.A1(new_n930), .A2(new_n332), .A3(new_n588), .ZN(new_n950));
  AOI21_X1  g749(.A(G218gat), .B1(new_n936), .B2(new_n684), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n950), .A2(new_n951), .ZN(G1355gat));
endmodule


