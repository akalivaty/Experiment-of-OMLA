

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U554 ( .A(KEYINPUT72), .B(n586), .ZN(n1007) );
  NOR2_X1 U555 ( .A1(n730), .A2(n729), .ZN(n732) );
  INV_X1 U556 ( .A(KEYINPUT29), .ZN(n714) );
  INV_X1 U557 ( .A(KEYINPUT106), .ZN(n782) );
  NAND2_X1 U558 ( .A1(n901), .A2(G137), .ZN(n535) );
  AND2_X1 U559 ( .A1(n1019), .A2(n830), .ZN(n518) );
  NOR2_X1 U560 ( .A1(n699), .A2(n698), .ZN(n701) );
  INV_X1 U561 ( .A(KEYINPUT100), .ZN(n731) );
  XNOR2_X1 U562 ( .A(n732), .B(n731), .ZN(n733) );
  XNOR2_X1 U563 ( .A(n744), .B(KEYINPUT32), .ZN(n753) );
  INV_X1 U564 ( .A(KEYINPUT17), .ZN(n533) );
  NOR2_X1 U565 ( .A1(n644), .A2(G651), .ZN(n654) );
  NOR2_X1 U566 ( .A1(G651), .A2(G543), .ZN(n519) );
  XNOR2_X1 U567 ( .A(n519), .B(KEYINPUT64), .ZN(n649) );
  NAND2_X1 U568 ( .A1(G89), .A2(n649), .ZN(n520) );
  XNOR2_X1 U569 ( .A(n520), .B(KEYINPUT4), .ZN(n522) );
  XOR2_X1 U570 ( .A(KEYINPUT0), .B(G543), .Z(n644) );
  INV_X1 U571 ( .A(G651), .ZN(n524) );
  NOR2_X1 U572 ( .A1(n644), .A2(n524), .ZN(n647) );
  NAND2_X1 U573 ( .A1(G76), .A2(n647), .ZN(n521) );
  NAND2_X1 U574 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U575 ( .A(KEYINPUT5), .B(n523), .ZN(n531) );
  NOR2_X1 U576 ( .A1(G543), .A2(n524), .ZN(n525) );
  XOR2_X2 U577 ( .A(KEYINPUT1), .B(n525), .Z(n653) );
  NAND2_X1 U578 ( .A1(G63), .A2(n653), .ZN(n527) );
  NAND2_X1 U579 ( .A1(G51), .A2(n654), .ZN(n526) );
  NAND2_X1 U580 ( .A1(n527), .A2(n526), .ZN(n529) );
  XOR2_X1 U581 ( .A(KEYINPUT74), .B(KEYINPUT6), .Z(n528) );
  XNOR2_X1 U582 ( .A(n529), .B(n528), .ZN(n530) );
  NAND2_X1 U583 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U584 ( .A(KEYINPUT7), .B(n532), .ZN(G168) );
  XOR2_X1 U585 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  AND2_X1 U586 ( .A1(G2104), .A2(G2105), .ZN(n897) );
  NAND2_X1 U587 ( .A1(n897), .A2(G113), .ZN(n536) );
  NOR2_X1 U588 ( .A1(G2104), .A2(G2105), .ZN(n534) );
  XNOR2_X2 U589 ( .A(n534), .B(n533), .ZN(n901) );
  NAND2_X1 U590 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U591 ( .A(n537), .B(KEYINPUT65), .ZN(n690) );
  INV_X1 U592 ( .A(G2104), .ZN(n554) );
  AND2_X1 U593 ( .A1(n554), .A2(G2105), .ZN(n895) );
  NAND2_X1 U594 ( .A1(G125), .A2(n895), .ZN(n688) );
  AND2_X1 U595 ( .A1(n690), .A2(n688), .ZN(n540) );
  NAND2_X1 U596 ( .A1(G2104), .A2(G101), .ZN(n538) );
  OR2_X1 U597 ( .A1(G2105), .A2(n538), .ZN(n539) );
  XOR2_X1 U598 ( .A(KEYINPUT23), .B(n539), .Z(n686) );
  AND2_X1 U599 ( .A1(n540), .A2(n686), .ZN(G160) );
  XOR2_X1 U600 ( .A(G2443), .B(G2446), .Z(n542) );
  XNOR2_X1 U601 ( .A(G2427), .B(G2451), .ZN(n541) );
  XNOR2_X1 U602 ( .A(n542), .B(n541), .ZN(n548) );
  XOR2_X1 U603 ( .A(G2430), .B(G2454), .Z(n544) );
  XNOR2_X1 U604 ( .A(G1348), .B(G1341), .ZN(n543) );
  XNOR2_X1 U605 ( .A(n544), .B(n543), .ZN(n546) );
  XOR2_X1 U606 ( .A(G2435), .B(G2438), .Z(n545) );
  XNOR2_X1 U607 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U608 ( .A(n548), .B(n547), .Z(n549) );
  AND2_X1 U609 ( .A1(G14), .A2(n549), .ZN(G401) );
  AND2_X1 U610 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U611 ( .A(G132), .ZN(G219) );
  INV_X1 U612 ( .A(G82), .ZN(G220) );
  INV_X1 U613 ( .A(G69), .ZN(G235) );
  NAND2_X1 U614 ( .A1(n897), .A2(G114), .ZN(n553) );
  INV_X1 U615 ( .A(KEYINPUT85), .ZN(n551) );
  NAND2_X1 U616 ( .A1(G138), .A2(n901), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(n552) );
  NAND2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n558) );
  NOR2_X1 U619 ( .A1(G2105), .A2(n554), .ZN(n903) );
  NAND2_X1 U620 ( .A1(G102), .A2(n903), .ZN(n556) );
  NAND2_X1 U621 ( .A1(G126), .A2(n895), .ZN(n555) );
  NAND2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U623 ( .A1(n558), .A2(n557), .ZN(G164) );
  NAND2_X1 U624 ( .A1(G77), .A2(n647), .ZN(n560) );
  NAND2_X1 U625 ( .A1(G90), .A2(n649), .ZN(n559) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(KEYINPUT9), .B(n561), .ZN(n565) );
  NAND2_X1 U628 ( .A1(G64), .A2(n653), .ZN(n563) );
  NAND2_X1 U629 ( .A1(G52), .A2(n654), .ZN(n562) );
  AND2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(G301) );
  INV_X1 U632 ( .A(G301), .ZN(G171) );
  NAND2_X1 U633 ( .A1(G7), .A2(G661), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n566), .B(KEYINPUT10), .ZN(n567) );
  XOR2_X1 U635 ( .A(KEYINPUT70), .B(n567), .Z(n835) );
  NAND2_X1 U636 ( .A1(n835), .A2(G567), .ZN(n568) );
  XNOR2_X1 U637 ( .A(n568), .B(KEYINPUT71), .ZN(n569) );
  XNOR2_X1 U638 ( .A(KEYINPUT11), .B(n569), .ZN(G234) );
  NAND2_X1 U639 ( .A1(G56), .A2(n653), .ZN(n570) );
  XOR2_X1 U640 ( .A(KEYINPUT14), .B(n570), .Z(n576) );
  NAND2_X1 U641 ( .A1(G81), .A2(n649), .ZN(n571) );
  XNOR2_X1 U642 ( .A(n571), .B(KEYINPUT12), .ZN(n573) );
  NAND2_X1 U643 ( .A1(G68), .A2(n647), .ZN(n572) );
  NAND2_X1 U644 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U645 ( .A(KEYINPUT13), .B(n574), .Z(n575) );
  NOR2_X1 U646 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U647 ( .A1(n654), .A2(G43), .ZN(n577) );
  NAND2_X1 U648 ( .A1(n578), .A2(n577), .ZN(n1001) );
  INV_X1 U649 ( .A(G860), .ZN(n614) );
  OR2_X1 U650 ( .A1(n1001), .A2(n614), .ZN(G153) );
  NAND2_X1 U651 ( .A1(n653), .A2(G66), .ZN(n580) );
  NAND2_X1 U652 ( .A1(G92), .A2(n649), .ZN(n579) );
  NAND2_X1 U653 ( .A1(n580), .A2(n579), .ZN(n584) );
  NAND2_X1 U654 ( .A1(G79), .A2(n647), .ZN(n582) );
  NAND2_X1 U655 ( .A1(G54), .A2(n654), .ZN(n581) );
  NAND2_X1 U656 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U657 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U658 ( .A(KEYINPUT15), .B(n585), .Z(n586) );
  NOR2_X1 U659 ( .A1(G868), .A2(n1007), .ZN(n587) );
  XNOR2_X1 U660 ( .A(n587), .B(KEYINPUT73), .ZN(n589) );
  NAND2_X1 U661 ( .A1(G868), .A2(G301), .ZN(n588) );
  NAND2_X1 U662 ( .A1(n589), .A2(n588), .ZN(G284) );
  NAND2_X1 U663 ( .A1(G78), .A2(n647), .ZN(n591) );
  NAND2_X1 U664 ( .A1(G91), .A2(n649), .ZN(n590) );
  NAND2_X1 U665 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n654), .A2(G53), .ZN(n592) );
  XOR2_X1 U667 ( .A(KEYINPUT68), .B(n592), .Z(n593) );
  NOR2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U669 ( .A1(n653), .A2(G65), .ZN(n595) );
  NAND2_X1 U670 ( .A1(n596), .A2(n595), .ZN(G299) );
  INV_X1 U671 ( .A(G868), .ZN(n668) );
  NOR2_X1 U672 ( .A1(G286), .A2(n668), .ZN(n598) );
  NOR2_X1 U673 ( .A1(G868), .A2(G299), .ZN(n597) );
  NOR2_X1 U674 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U675 ( .A1(n614), .A2(G559), .ZN(n599) );
  NAND2_X1 U676 ( .A1(n599), .A2(n1007), .ZN(n600) );
  XNOR2_X1 U677 ( .A(n600), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U678 ( .A1(G868), .A2(n1001), .ZN(n603) );
  NAND2_X1 U679 ( .A1(n1007), .A2(G868), .ZN(n601) );
  NOR2_X1 U680 ( .A1(G559), .A2(n601), .ZN(n602) );
  NOR2_X1 U681 ( .A1(n603), .A2(n602), .ZN(G282) );
  NAND2_X1 U682 ( .A1(G123), .A2(n895), .ZN(n604) );
  XOR2_X1 U683 ( .A(KEYINPUT75), .B(n604), .Z(n605) );
  XNOR2_X1 U684 ( .A(n605), .B(KEYINPUT18), .ZN(n607) );
  NAND2_X1 U685 ( .A1(G111), .A2(n897), .ZN(n606) );
  NAND2_X1 U686 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U687 ( .A1(G135), .A2(n901), .ZN(n609) );
  NAND2_X1 U688 ( .A1(G99), .A2(n903), .ZN(n608) );
  NAND2_X1 U689 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U690 ( .A1(n611), .A2(n610), .ZN(n975) );
  XNOR2_X1 U691 ( .A(n975), .B(G2096), .ZN(n612) );
  INV_X1 U692 ( .A(G2100), .ZN(n849) );
  NAND2_X1 U693 ( .A1(n612), .A2(n849), .ZN(G156) );
  NAND2_X1 U694 ( .A1(n1007), .A2(G559), .ZN(n613) );
  XOR2_X1 U695 ( .A(n1001), .B(n613), .Z(n665) );
  NAND2_X1 U696 ( .A1(n614), .A2(n665), .ZN(n621) );
  NAND2_X1 U697 ( .A1(n653), .A2(G67), .ZN(n616) );
  NAND2_X1 U698 ( .A1(G93), .A2(n649), .ZN(n615) );
  NAND2_X1 U699 ( .A1(n616), .A2(n615), .ZN(n620) );
  NAND2_X1 U700 ( .A1(G80), .A2(n647), .ZN(n618) );
  NAND2_X1 U701 ( .A1(G55), .A2(n654), .ZN(n617) );
  NAND2_X1 U702 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U703 ( .A1(n620), .A2(n619), .ZN(n667) );
  XOR2_X1 U704 ( .A(n621), .B(n667), .Z(G145) );
  NAND2_X1 U705 ( .A1(G62), .A2(n653), .ZN(n622) );
  XOR2_X1 U706 ( .A(KEYINPUT80), .B(n622), .Z(n627) );
  NAND2_X1 U707 ( .A1(G75), .A2(n647), .ZN(n624) );
  NAND2_X1 U708 ( .A1(G88), .A2(n649), .ZN(n623) );
  NAND2_X1 U709 ( .A1(n624), .A2(n623), .ZN(n625) );
  XOR2_X1 U710 ( .A(KEYINPUT81), .B(n625), .Z(n626) );
  NOR2_X1 U711 ( .A1(n627), .A2(n626), .ZN(n629) );
  NAND2_X1 U712 ( .A1(n654), .A2(G50), .ZN(n628) );
  NAND2_X1 U713 ( .A1(n629), .A2(n628), .ZN(G303) );
  NAND2_X1 U714 ( .A1(G73), .A2(n647), .ZN(n630) );
  XNOR2_X1 U715 ( .A(n630), .B(KEYINPUT2), .ZN(n637) );
  NAND2_X1 U716 ( .A1(n654), .A2(G48), .ZN(n632) );
  NAND2_X1 U717 ( .A1(G86), .A2(n649), .ZN(n631) );
  NAND2_X1 U718 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U719 ( .A1(G61), .A2(n653), .ZN(n633) );
  XNOR2_X1 U720 ( .A(KEYINPUT79), .B(n633), .ZN(n634) );
  NOR2_X1 U721 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U722 ( .A1(n637), .A2(n636), .ZN(G305) );
  NAND2_X1 U723 ( .A1(G651), .A2(G74), .ZN(n638) );
  XNOR2_X1 U724 ( .A(n638), .B(KEYINPUT76), .ZN(n640) );
  NAND2_X1 U725 ( .A1(G49), .A2(n654), .ZN(n639) );
  NAND2_X1 U726 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U727 ( .A(KEYINPUT77), .B(n641), .Z(n642) );
  NOR2_X1 U728 ( .A1(n653), .A2(n642), .ZN(n643) );
  XNOR2_X1 U729 ( .A(n643), .B(KEYINPUT78), .ZN(n646) );
  NAND2_X1 U730 ( .A1(G87), .A2(n644), .ZN(n645) );
  NAND2_X1 U731 ( .A1(n646), .A2(n645), .ZN(G288) );
  NAND2_X1 U732 ( .A1(n647), .A2(G72), .ZN(n648) );
  XNOR2_X1 U733 ( .A(n648), .B(KEYINPUT66), .ZN(n651) );
  NAND2_X1 U734 ( .A1(G85), .A2(n649), .ZN(n650) );
  NAND2_X1 U735 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U736 ( .A(KEYINPUT67), .B(n652), .ZN(n658) );
  NAND2_X1 U737 ( .A1(G60), .A2(n653), .ZN(n656) );
  NAND2_X1 U738 ( .A1(G47), .A2(n654), .ZN(n655) );
  AND2_X1 U739 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U740 ( .A1(n658), .A2(n657), .ZN(G290) );
  XNOR2_X1 U741 ( .A(KEYINPUT19), .B(KEYINPUT82), .ZN(n659) );
  XNOR2_X1 U742 ( .A(n659), .B(n667), .ZN(n660) );
  XOR2_X1 U743 ( .A(G303), .B(n660), .Z(n663) );
  XOR2_X1 U744 ( .A(G299), .B(G305), .Z(n661) );
  XNOR2_X1 U745 ( .A(n661), .B(G288), .ZN(n662) );
  XNOR2_X1 U746 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U747 ( .A(n664), .B(G290), .ZN(n843) );
  XOR2_X1 U748 ( .A(n843), .B(n665), .Z(n666) );
  NOR2_X1 U749 ( .A1(n668), .A2(n666), .ZN(n670) );
  AND2_X1 U750 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U751 ( .A1(n670), .A2(n669), .ZN(G295) );
  NAND2_X1 U752 ( .A1(G2084), .A2(G2078), .ZN(n671) );
  XOR2_X1 U753 ( .A(KEYINPUT20), .B(n671), .Z(n672) );
  NAND2_X1 U754 ( .A1(G2090), .A2(n672), .ZN(n673) );
  XNOR2_X1 U755 ( .A(KEYINPUT21), .B(n673), .ZN(n674) );
  NAND2_X1 U756 ( .A1(n674), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U757 ( .A(KEYINPUT69), .B(G57), .ZN(G237) );
  XNOR2_X1 U758 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U759 ( .A1(G235), .A2(G237), .ZN(n675) );
  NAND2_X1 U760 ( .A1(G120), .A2(n675), .ZN(n676) );
  XNOR2_X1 U761 ( .A(KEYINPUT83), .B(n676), .ZN(n677) );
  NAND2_X1 U762 ( .A1(n677), .A2(G108), .ZN(n841) );
  NAND2_X1 U763 ( .A1(G567), .A2(n841), .ZN(n682) );
  NOR2_X1 U764 ( .A1(G220), .A2(G219), .ZN(n678) );
  XOR2_X1 U765 ( .A(KEYINPUT22), .B(n678), .Z(n679) );
  NOR2_X1 U766 ( .A1(G218), .A2(n679), .ZN(n680) );
  NAND2_X1 U767 ( .A1(G96), .A2(n680), .ZN(n842) );
  NAND2_X1 U768 ( .A1(G2106), .A2(n842), .ZN(n681) );
  NAND2_X1 U769 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U770 ( .A(KEYINPUT84), .B(n683), .ZN(n918) );
  NAND2_X1 U771 ( .A1(G661), .A2(G483), .ZN(n684) );
  NOR2_X1 U772 ( .A1(n918), .A2(n684), .ZN(n840) );
  NAND2_X1 U773 ( .A1(n840), .A2(G36), .ZN(G176) );
  INV_X1 U774 ( .A(G299), .ZN(n709) );
  OR2_X1 U775 ( .A1(G164), .A2(G1384), .ZN(n784) );
  AND2_X1 U776 ( .A1(G40), .A2(n686), .ZN(n687) );
  AND2_X1 U777 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U778 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U779 ( .A(n691), .B(KEYINPUT86), .ZN(n786) );
  OR2_X2 U780 ( .A1(n784), .A2(n786), .ZN(n736) );
  INV_X1 U781 ( .A(n736), .ZN(n717) );
  NAND2_X1 U782 ( .A1(n717), .A2(G2072), .ZN(n692) );
  XNOR2_X1 U783 ( .A(n692), .B(KEYINPUT27), .ZN(n694) );
  AND2_X1 U784 ( .A1(G1956), .A2(n736), .ZN(n693) );
  NOR2_X1 U785 ( .A1(n694), .A2(n693), .ZN(n708) );
  NOR2_X1 U786 ( .A1(n709), .A2(n708), .ZN(n695) );
  XOR2_X1 U787 ( .A(n695), .B(KEYINPUT28), .Z(n713) );
  INV_X1 U788 ( .A(G1996), .ZN(n860) );
  NOR2_X1 U789 ( .A1(n736), .A2(n860), .ZN(n696) );
  XNOR2_X1 U790 ( .A(n696), .B(KEYINPUT26), .ZN(n699) );
  AND2_X1 U791 ( .A1(n736), .A2(G1341), .ZN(n697) );
  OR2_X1 U792 ( .A1(n697), .A2(n1001), .ZN(n698) );
  NOR2_X1 U793 ( .A1(n701), .A2(n1007), .ZN(n700) );
  XOR2_X1 U794 ( .A(n700), .B(KEYINPUT98), .Z(n707) );
  NAND2_X1 U795 ( .A1(n701), .A2(n1007), .ZN(n705) );
  NOR2_X1 U796 ( .A1(G2067), .A2(n736), .ZN(n703) );
  NOR2_X1 U797 ( .A1(n717), .A2(G1348), .ZN(n702) );
  NOR2_X1 U798 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U799 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U800 ( .A1(n707), .A2(n706), .ZN(n711) );
  NAND2_X1 U801 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U802 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U803 ( .A1(n713), .A2(n712), .ZN(n715) );
  XNOR2_X1 U804 ( .A(n715), .B(n714), .ZN(n721) );
  INV_X1 U805 ( .A(G1961), .ZN(n1006) );
  NAND2_X1 U806 ( .A1(n736), .A2(n1006), .ZN(n719) );
  XOR2_X1 U807 ( .A(G2078), .B(KEYINPUT25), .Z(n716) );
  XNOR2_X1 U808 ( .A(KEYINPUT97), .B(n716), .ZN(n920) );
  NAND2_X1 U809 ( .A1(n717), .A2(n920), .ZN(n718) );
  NAND2_X1 U810 ( .A1(n719), .A2(n718), .ZN(n728) );
  NAND2_X1 U811 ( .A1(n728), .A2(G171), .ZN(n720) );
  NAND2_X1 U812 ( .A1(n721), .A2(n720), .ZN(n735) );
  NAND2_X1 U813 ( .A1(G8), .A2(n736), .ZN(n773) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n773), .ZN(n748) );
  NOR2_X1 U815 ( .A1(G2084), .A2(n736), .ZN(n722) );
  XNOR2_X1 U816 ( .A(n722), .B(KEYINPUT96), .ZN(n745) );
  INV_X1 U817 ( .A(n745), .ZN(n723) );
  NAND2_X1 U818 ( .A1(n723), .A2(G8), .ZN(n724) );
  NOR2_X1 U819 ( .A1(n748), .A2(n724), .ZN(n726) );
  XNOR2_X1 U820 ( .A(KEYINPUT99), .B(KEYINPUT30), .ZN(n725) );
  XNOR2_X1 U821 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U822 ( .A1(n727), .A2(G168), .ZN(n730) );
  NOR2_X1 U823 ( .A1(G171), .A2(n728), .ZN(n729) );
  XNOR2_X1 U824 ( .A(KEYINPUT31), .B(n733), .ZN(n734) );
  NAND2_X1 U825 ( .A1(n735), .A2(n734), .ZN(n746) );
  NAND2_X1 U826 ( .A1(n746), .A2(G286), .ZN(n741) );
  NOR2_X1 U827 ( .A1(G1971), .A2(n773), .ZN(n738) );
  NOR2_X1 U828 ( .A1(G2090), .A2(n736), .ZN(n737) );
  NOR2_X1 U829 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U830 ( .A1(n739), .A2(G303), .ZN(n740) );
  NAND2_X1 U831 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U832 ( .A(n742), .B(KEYINPUT102), .ZN(n743) );
  NAND2_X1 U833 ( .A1(n743), .A2(G8), .ZN(n744) );
  NAND2_X1 U834 ( .A1(n745), .A2(G8), .ZN(n751) );
  INV_X1 U835 ( .A(n746), .ZN(n747) );
  NOR2_X1 U836 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U837 ( .A(KEYINPUT101), .B(n749), .Z(n750) );
  NAND2_X1 U838 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U839 ( .A1(n753), .A2(n752), .ZN(n771) );
  NOR2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n1011) );
  NOR2_X1 U841 ( .A1(G1971), .A2(G303), .ZN(n754) );
  XOR2_X1 U842 ( .A(n754), .B(KEYINPUT103), .Z(n755) );
  NOR2_X1 U843 ( .A1(n1011), .A2(n755), .ZN(n756) );
  NAND2_X1 U844 ( .A1(n771), .A2(n756), .ZN(n757) );
  NAND2_X1 U845 ( .A1(G1976), .A2(G288), .ZN(n1012) );
  NAND2_X1 U846 ( .A1(n757), .A2(n1012), .ZN(n758) );
  XNOR2_X1 U847 ( .A(n758), .B(KEYINPUT104), .ZN(n764) );
  NAND2_X1 U848 ( .A1(n1011), .A2(KEYINPUT33), .ZN(n759) );
  NOR2_X1 U849 ( .A1(n773), .A2(n759), .ZN(n762) );
  XNOR2_X1 U850 ( .A(KEYINPUT105), .B(G1981), .ZN(n760) );
  XNOR2_X1 U851 ( .A(n760), .B(G305), .ZN(n1021) );
  INV_X1 U852 ( .A(n1021), .ZN(n761) );
  OR2_X1 U853 ( .A1(n762), .A2(n761), .ZN(n776) );
  OR2_X1 U854 ( .A1(n773), .A2(n776), .ZN(n763) );
  NOR2_X1 U855 ( .A1(n764), .A2(n763), .ZN(n781) );
  NOR2_X1 U856 ( .A1(G1981), .A2(G305), .ZN(n765) );
  XOR2_X1 U857 ( .A(n765), .B(KEYINPUT94), .Z(n766) );
  XNOR2_X1 U858 ( .A(KEYINPUT24), .B(n766), .ZN(n767) );
  NOR2_X1 U859 ( .A1(n773), .A2(n767), .ZN(n768) );
  XNOR2_X1 U860 ( .A(KEYINPUT95), .B(n768), .ZN(n775) );
  NOR2_X1 U861 ( .A1(G2090), .A2(G303), .ZN(n769) );
  NAND2_X1 U862 ( .A1(G8), .A2(n769), .ZN(n770) );
  NAND2_X1 U863 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U864 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U865 ( .A1(n775), .A2(n774), .ZN(n779) );
  INV_X1 U866 ( .A(n776), .ZN(n777) );
  NAND2_X1 U867 ( .A1(n777), .A2(KEYINPUT33), .ZN(n778) );
  NAND2_X1 U868 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n783) );
  XNOR2_X1 U870 ( .A(n783), .B(n782), .ZN(n820) );
  INV_X1 U871 ( .A(n784), .ZN(n785) );
  NOR2_X1 U872 ( .A1(n786), .A2(n785), .ZN(n830) );
  XNOR2_X1 U873 ( .A(G2067), .B(KEYINPUT37), .ZN(n828) );
  NAND2_X1 U874 ( .A1(G140), .A2(n901), .ZN(n788) );
  NAND2_X1 U875 ( .A1(G104), .A2(n903), .ZN(n787) );
  NAND2_X1 U876 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U877 ( .A(KEYINPUT34), .B(n789), .ZN(n794) );
  NAND2_X1 U878 ( .A1(G116), .A2(n897), .ZN(n791) );
  NAND2_X1 U879 ( .A1(G128), .A2(n895), .ZN(n790) );
  NAND2_X1 U880 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U881 ( .A(KEYINPUT35), .B(n792), .Z(n793) );
  NOR2_X1 U882 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U883 ( .A(KEYINPUT36), .B(n795), .ZN(n876) );
  NOR2_X1 U884 ( .A1(n828), .A2(n876), .ZN(n971) );
  NAND2_X1 U885 ( .A1(n830), .A2(n971), .ZN(n826) );
  XOR2_X1 U886 ( .A(KEYINPUT88), .B(G1991), .Z(n924) );
  NAND2_X1 U887 ( .A1(G131), .A2(n901), .ZN(n797) );
  NAND2_X1 U888 ( .A1(G119), .A2(n895), .ZN(n796) );
  NAND2_X1 U889 ( .A1(n797), .A2(n796), .ZN(n800) );
  NAND2_X1 U890 ( .A1(G107), .A2(n897), .ZN(n798) );
  XNOR2_X1 U891 ( .A(KEYINPUT87), .B(n798), .ZN(n799) );
  NOR2_X1 U892 ( .A1(n800), .A2(n799), .ZN(n802) );
  NAND2_X1 U893 ( .A1(n903), .A2(G95), .ZN(n801) );
  AND2_X1 U894 ( .A1(n802), .A2(n801), .ZN(n892) );
  NOR2_X1 U895 ( .A1(n924), .A2(n892), .ZN(n814) );
  XOR2_X1 U896 ( .A(KEYINPUT38), .B(KEYINPUT90), .Z(n804) );
  NAND2_X1 U897 ( .A1(G105), .A2(n903), .ZN(n803) );
  XNOR2_X1 U898 ( .A(n804), .B(n803), .ZN(n807) );
  NAND2_X1 U899 ( .A1(n897), .A2(G117), .ZN(n805) );
  XNOR2_X1 U900 ( .A(KEYINPUT89), .B(n805), .ZN(n806) );
  NOR2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n809) );
  NAND2_X1 U902 ( .A1(n895), .A2(G129), .ZN(n808) );
  NAND2_X1 U903 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U904 ( .A(n810), .B(KEYINPUT91), .ZN(n812) );
  NAND2_X1 U905 ( .A1(G141), .A2(n901), .ZN(n811) );
  NAND2_X1 U906 ( .A1(n812), .A2(n811), .ZN(n888) );
  AND2_X1 U907 ( .A1(n888), .A2(G1996), .ZN(n813) );
  NOR2_X1 U908 ( .A1(n814), .A2(n813), .ZN(n977) );
  XOR2_X1 U909 ( .A(n830), .B(KEYINPUT92), .Z(n815) );
  NOR2_X1 U910 ( .A1(n977), .A2(n815), .ZN(n823) );
  INV_X1 U911 ( .A(n823), .ZN(n816) );
  NAND2_X1 U912 ( .A1(n826), .A2(n816), .ZN(n817) );
  XOR2_X1 U913 ( .A(KEYINPUT93), .B(n817), .Z(n818) );
  XNOR2_X1 U914 ( .A(G1986), .B(G290), .ZN(n1019) );
  NOR2_X1 U915 ( .A1(n818), .A2(n518), .ZN(n819) );
  NAND2_X1 U916 ( .A1(n820), .A2(n819), .ZN(n833) );
  NOR2_X1 U917 ( .A1(G1996), .A2(n888), .ZN(n981) );
  AND2_X1 U918 ( .A1(n924), .A2(n892), .ZN(n970) );
  NOR2_X1 U919 ( .A1(G1986), .A2(G290), .ZN(n821) );
  NOR2_X1 U920 ( .A1(n970), .A2(n821), .ZN(n822) );
  NOR2_X1 U921 ( .A1(n823), .A2(n822), .ZN(n824) );
  NOR2_X1 U922 ( .A1(n981), .A2(n824), .ZN(n825) );
  XNOR2_X1 U923 ( .A(n825), .B(KEYINPUT39), .ZN(n827) );
  NAND2_X1 U924 ( .A1(n827), .A2(n826), .ZN(n829) );
  NAND2_X1 U925 ( .A1(n828), .A2(n876), .ZN(n986) );
  NAND2_X1 U926 ( .A1(n829), .A2(n986), .ZN(n831) );
  NAND2_X1 U927 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U928 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U929 ( .A(KEYINPUT40), .B(n834), .ZN(G329) );
  NAND2_X1 U930 ( .A1(G2106), .A2(n835), .ZN(G217) );
  INV_X1 U931 ( .A(n835), .ZN(G223) );
  NAND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n837) );
  INV_X1 U933 ( .A(G661), .ZN(n836) );
  NOR2_X1 U934 ( .A1(n837), .A2(n836), .ZN(n838) );
  XNOR2_X1 U935 ( .A(n838), .B(KEYINPUT107), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U937 ( .A1(n840), .A2(n839), .ZN(G188) );
  XOR2_X1 U938 ( .A(G120), .B(KEYINPUT108), .Z(G236) );
  INV_X1 U940 ( .A(G108), .ZN(G238) );
  INV_X1 U941 ( .A(G96), .ZN(G221) );
  NOR2_X1 U942 ( .A1(n842), .A2(n841), .ZN(G325) );
  INV_X1 U943 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U944 ( .A(G286), .B(n843), .ZN(n846) );
  XOR2_X1 U945 ( .A(KEYINPUT114), .B(G171), .Z(n844) );
  XNOR2_X1 U946 ( .A(n844), .B(n1007), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n847), .B(n1001), .ZN(n848) );
  NOR2_X1 U949 ( .A1(G37), .A2(n848), .ZN(G397) );
  XNOR2_X1 U950 ( .A(n849), .B(G2096), .ZN(n851) );
  XNOR2_X1 U951 ( .A(KEYINPUT42), .B(G2678), .ZN(n850) );
  XNOR2_X1 U952 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U953 ( .A(KEYINPUT43), .B(G2090), .Z(n853) );
  XNOR2_X1 U954 ( .A(G2067), .B(G2072), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U956 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U957 ( .A(G2084), .B(G2078), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n857), .B(n856), .ZN(G227) );
  XNOR2_X1 U959 ( .A(G1956), .B(n1006), .ZN(n859) );
  XNOR2_X1 U960 ( .A(G1986), .B(G1981), .ZN(n858) );
  XNOR2_X1 U961 ( .A(n859), .B(n858), .ZN(n864) );
  XOR2_X1 U962 ( .A(G1971), .B(G1976), .Z(n862) );
  XOR2_X1 U963 ( .A(n860), .B(G1991), .Z(n861) );
  XNOR2_X1 U964 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U965 ( .A(n864), .B(n863), .Z(n866) );
  XNOR2_X1 U966 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n865) );
  XNOR2_X1 U967 ( .A(n866), .B(n865), .ZN(n868) );
  XOR2_X1 U968 ( .A(G1966), .B(G2474), .Z(n867) );
  XNOR2_X1 U969 ( .A(n868), .B(n867), .ZN(G229) );
  NAND2_X1 U970 ( .A1(G124), .A2(n895), .ZN(n869) );
  XNOR2_X1 U971 ( .A(n869), .B(KEYINPUT44), .ZN(n871) );
  NAND2_X1 U972 ( .A1(n897), .A2(G112), .ZN(n870) );
  NAND2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n875) );
  NAND2_X1 U974 ( .A1(G136), .A2(n901), .ZN(n873) );
  NAND2_X1 U975 ( .A1(G100), .A2(n903), .ZN(n872) );
  NAND2_X1 U976 ( .A1(n873), .A2(n872), .ZN(n874) );
  NOR2_X1 U977 ( .A1(n875), .A2(n874), .ZN(G162) );
  XNOR2_X1 U978 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n878) );
  XNOR2_X1 U979 ( .A(n876), .B(G162), .ZN(n877) );
  XNOR2_X1 U980 ( .A(n878), .B(n877), .ZN(n887) );
  NAND2_X1 U981 ( .A1(G139), .A2(n901), .ZN(n880) );
  NAND2_X1 U982 ( .A1(G103), .A2(n903), .ZN(n879) );
  NAND2_X1 U983 ( .A1(n880), .A2(n879), .ZN(n886) );
  NAND2_X1 U984 ( .A1(n897), .A2(G115), .ZN(n881) );
  XOR2_X1 U985 ( .A(KEYINPUT113), .B(n881), .Z(n883) );
  NAND2_X1 U986 ( .A1(n895), .A2(G127), .ZN(n882) );
  NAND2_X1 U987 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U988 ( .A(KEYINPUT47), .B(n884), .Z(n885) );
  NOR2_X1 U989 ( .A1(n886), .A2(n885), .ZN(n988) );
  XOR2_X1 U990 ( .A(n887), .B(n988), .Z(n890) );
  XOR2_X1 U991 ( .A(G164), .B(n888), .Z(n889) );
  XNOR2_X1 U992 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U993 ( .A(n891), .B(n975), .Z(n894) );
  XNOR2_X1 U994 ( .A(G160), .B(n892), .ZN(n893) );
  XNOR2_X1 U995 ( .A(n894), .B(n893), .ZN(n910) );
  NAND2_X1 U996 ( .A1(G130), .A2(n895), .ZN(n896) );
  XNOR2_X1 U997 ( .A(n896), .B(KEYINPUT110), .ZN(n900) );
  NAND2_X1 U998 ( .A1(G118), .A2(n897), .ZN(n898) );
  XOR2_X1 U999 ( .A(KEYINPUT111), .B(n898), .Z(n899) );
  NAND2_X1 U1000 ( .A1(n900), .A2(n899), .ZN(n908) );
  NAND2_X1 U1001 ( .A1(n901), .A2(G142), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n902), .B(KEYINPUT112), .ZN(n905) );
  NAND2_X1 U1003 ( .A1(G106), .A2(n903), .ZN(n904) );
  NAND2_X1 U1004 ( .A1(n905), .A2(n904), .ZN(n906) );
  XOR2_X1 U1005 ( .A(KEYINPUT45), .B(n906), .Z(n907) );
  NOR2_X1 U1006 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(n910), .B(n909), .ZN(n911) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n911), .ZN(G395) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n912) );
  XNOR2_X1 U1010 ( .A(KEYINPUT49), .B(n912), .ZN(n913) );
  NOR2_X1 U1011 ( .A1(G397), .A2(n913), .ZN(n917) );
  NOR2_X1 U1012 ( .A1(n918), .A2(G401), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(KEYINPUT115), .B(n914), .ZN(n915) );
  NOR2_X1 U1014 ( .A1(G395), .A2(n915), .ZN(n916) );
  NAND2_X1 U1015 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(n918), .ZN(G319) );
  INV_X1 U1018 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U1019 ( .A(G2090), .B(G35), .ZN(n933) );
  XOR2_X1 U1020 ( .A(G2072), .B(G33), .Z(n919) );
  NAND2_X1 U1021 ( .A1(G28), .A2(n919), .ZN(n930) );
  XNOR2_X1 U1022 ( .A(n920), .B(G27), .ZN(n922) );
  XOR2_X1 U1023 ( .A(G1996), .B(G32), .Z(n921) );
  NAND2_X1 U1024 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1025 ( .A(KEYINPUT119), .B(n923), .ZN(n928) );
  XOR2_X1 U1026 ( .A(n924), .B(G25), .Z(n926) );
  XNOR2_X1 U1027 ( .A(G2067), .B(G26), .ZN(n925) );
  NOR2_X1 U1028 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1031 ( .A(KEYINPUT53), .B(n931), .ZN(n932) );
  NOR2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n936) );
  XOR2_X1 U1033 ( .A(G2084), .B(G34), .Z(n934) );
  XNOR2_X1 U1034 ( .A(KEYINPUT54), .B(n934), .ZN(n935) );
  NAND2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n939) );
  NOR2_X1 U1036 ( .A1(G29), .A2(KEYINPUT55), .ZN(n937) );
  NAND2_X1 U1037 ( .A1(n939), .A2(n937), .ZN(n938) );
  NAND2_X1 U1038 ( .A1(G11), .A2(n938), .ZN(n969) );
  INV_X1 U1039 ( .A(KEYINPUT55), .ZN(n995) );
  OR2_X1 U1040 ( .A1(n995), .A2(n939), .ZN(n967) );
  XNOR2_X1 U1041 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n964) );
  XNOR2_X1 U1042 ( .A(G1348), .B(KEYINPUT59), .ZN(n940) );
  XNOR2_X1 U1043 ( .A(n940), .B(G4), .ZN(n944) );
  XNOR2_X1 U1044 ( .A(G1981), .B(G6), .ZN(n942) );
  XNOR2_X1 U1045 ( .A(G1341), .B(G19), .ZN(n941) );
  NOR2_X1 U1046 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1047 ( .A1(n944), .A2(n943), .ZN(n947) );
  XOR2_X1 U1048 ( .A(G20), .B(G1956), .Z(n945) );
  XNOR2_X1 U1049 ( .A(KEYINPUT123), .B(n945), .ZN(n946) );
  NOR2_X1 U1050 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1051 ( .A(KEYINPUT60), .B(n948), .ZN(n950) );
  XOR2_X1 U1052 ( .A(G1961), .B(G5), .Z(n949) );
  NAND2_X1 U1053 ( .A1(n950), .A2(n949), .ZN(n953) );
  XNOR2_X1 U1054 ( .A(G21), .B(G1966), .ZN(n951) );
  XNOR2_X1 U1055 ( .A(KEYINPUT124), .B(n951), .ZN(n952) );
  NOR2_X1 U1056 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1057 ( .A(KEYINPUT125), .B(n954), .Z(n962) );
  XNOR2_X1 U1058 ( .A(G1976), .B(G23), .ZN(n956) );
  XNOR2_X1 U1059 ( .A(G22), .B(G1971), .ZN(n955) );
  NOR2_X1 U1060 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1061 ( .A(KEYINPUT126), .B(n957), .Z(n959) );
  XNOR2_X1 U1062 ( .A(G1986), .B(G24), .ZN(n958) );
  NOR2_X1 U1063 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1064 ( .A(KEYINPUT58), .B(n960), .ZN(n961) );
  NAND2_X1 U1065 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1066 ( .A(n964), .B(n963), .ZN(n965) );
  INV_X1 U1067 ( .A(G16), .ZN(n1000) );
  NAND2_X1 U1068 ( .A1(n965), .A2(n1000), .ZN(n966) );
  NAND2_X1 U1069 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1070 ( .A1(n969), .A2(n968), .ZN(n999) );
  XNOR2_X1 U1071 ( .A(G160), .B(G2084), .ZN(n973) );
  NOR2_X1 U1072 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1073 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1074 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1075 ( .A(KEYINPUT116), .B(n976), .ZN(n978) );
  NAND2_X1 U1076 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1077 ( .A(KEYINPUT117), .B(n979), .Z(n984) );
  XOR2_X1 U1078 ( .A(G2090), .B(G162), .Z(n980) );
  NOR2_X1 U1079 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1080 ( .A(n982), .B(KEYINPUT51), .ZN(n983) );
  NOR2_X1 U1081 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1082 ( .A(n985), .B(KEYINPUT118), .ZN(n987) );
  NAND2_X1 U1083 ( .A1(n987), .A2(n986), .ZN(n993) );
  XOR2_X1 U1084 ( .A(G2072), .B(n988), .Z(n990) );
  XOR2_X1 U1085 ( .A(G164), .B(G2078), .Z(n989) );
  NOR2_X1 U1086 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1087 ( .A(KEYINPUT50), .B(n991), .Z(n992) );
  NOR2_X1 U1088 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1089 ( .A(KEYINPUT52), .B(n994), .ZN(n996) );
  NAND2_X1 U1090 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1091 ( .A1(n997), .A2(G29), .ZN(n998) );
  NAND2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1030) );
  XNOR2_X1 U1093 ( .A(n1000), .B(KEYINPUT56), .ZN(n1028) );
  XOR2_X1 U1094 ( .A(n1001), .B(G1341), .Z(n1003) );
  XOR2_X1 U1095 ( .A(G299), .B(G1956), .Z(n1002) );
  NAND2_X1 U1096 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  XOR2_X1 U1097 ( .A(G1971), .B(G166), .Z(n1004) );
  NOR2_X1 U1098 ( .A1(n1005), .A2(n1004), .ZN(n1017) );
  XOR2_X1 U1099 ( .A(G171), .B(n1006), .Z(n1009) );
  XNOR2_X1 U1100 ( .A(G1348), .B(n1007), .ZN(n1008) );
  NAND2_X1 U1101 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1102 ( .A(n1010), .B(KEYINPUT120), .ZN(n1015) );
  INV_X1 U1103 ( .A(n1011), .ZN(n1013) );
  NAND2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1108 ( .A(KEYINPUT121), .B(n1020), .ZN(n1025) );
  XNOR2_X1 U1109 ( .A(G1966), .B(G168), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1111 ( .A(KEYINPUT57), .B(n1023), .Z(n1024) );
  NOR2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1113 ( .A(KEYINPUT122), .B(n1026), .ZN(n1027) );
  NOR2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1116 ( .A(n1031), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1117 ( .A(G150), .ZN(G311) );
endmodule

