//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938;
  INV_X1    g000(.A(G475), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NOR3_X1   g003(.A1(new_n189), .A2(KEYINPUT16), .A3(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT77), .A2(G125), .ZN(new_n191));
  INV_X1    g005(.A(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  NAND3_X1  g007(.A1(KEYINPUT77), .A2(G125), .A3(G140), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n190), .B1(new_n195), .B2(KEYINPUT16), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  XNOR2_X1  g011(.A(new_n196), .B(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n199), .A2(KEYINPUT92), .ZN(new_n200));
  INV_X1    g014(.A(G237), .ZN(new_n201));
  INV_X1    g015(.A(G953), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G214), .ZN(new_n203));
  XNOR2_X1  g017(.A(new_n200), .B(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT17), .A3(G131), .ZN(new_n205));
  XNOR2_X1  g019(.A(new_n204), .B(G131), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n198), .B(new_n205), .C1(new_n206), .C2(KEYINPUT17), .ZN(new_n207));
  XOR2_X1   g021(.A(G113), .B(G122), .Z(new_n208));
  XNOR2_X1  g022(.A(new_n208), .B(KEYINPUT94), .ZN(new_n209));
  INV_X1    g023(.A(G104), .ZN(new_n210));
  XNOR2_X1  g024(.A(new_n209), .B(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(G125), .B(G140), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(new_n197), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT78), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n213), .B(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT93), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n195), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n193), .A2(KEYINPUT93), .A3(new_n194), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n215), .B1(new_n219), .B2(new_n197), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT18), .A2(G131), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n204), .B(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n207), .A2(new_n211), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n212), .A2(KEYINPUT19), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n225), .B1(new_n219), .B2(KEYINPUT19), .ZN(new_n226));
  OR2_X1    g040(.A1(new_n226), .A2(G146), .ZN(new_n227));
  OR2_X1    g041(.A1(new_n204), .A2(G131), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n204), .A2(G131), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n228), .A2(new_n229), .B1(G146), .B2(new_n196), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n211), .B1(new_n231), .B2(new_n223), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n187), .B(new_n188), .C1(new_n224), .C2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT20), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n207), .A2(new_n211), .A3(new_n223), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n227), .A2(new_n230), .B1(new_n220), .B2(new_n222), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n236), .B1(new_n211), .B2(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n238), .A2(KEYINPUT20), .A3(new_n187), .A4(new_n188), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT95), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n207), .A2(new_n223), .ZN(new_n242));
  INV_X1    g056(.A(new_n211), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(G902), .B1(new_n244), .B2(new_n236), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n241), .A3(new_n243), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n187), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n240), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n202), .A2(G952), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n250), .B1(G234), .B2(G237), .ZN(new_n251));
  INV_X1    g065(.A(G234), .ZN(new_n252));
  OAI211_X1 g066(.A(G902), .B(G953), .C1(new_n252), .C2(new_n201), .ZN(new_n253));
  XOR2_X1   g067(.A(new_n253), .B(KEYINPUT97), .Z(new_n254));
  XOR2_X1   g068(.A(KEYINPUT21), .B(G898), .Z(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n251), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G134), .ZN(new_n258));
  XNOR2_X1  g072(.A(G128), .B(G143), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT96), .B(KEYINPUT13), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n199), .A2(G128), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n261), .B1(new_n262), .B2(new_n260), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n259), .A2(new_n258), .ZN(new_n264));
  XNOR2_X1  g078(.A(G116), .B(G122), .ZN(new_n265));
  INV_X1    g079(.A(G107), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n265), .B(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n263), .A2(new_n264), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n259), .B(new_n258), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n265), .A2(new_n266), .ZN(new_n270));
  INV_X1    g084(.A(G116), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT14), .B1(new_n271), .B2(G122), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n265), .B1(KEYINPUT14), .B2(new_n266), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n269), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n268), .A2(new_n275), .ZN(new_n276));
  XOR2_X1   g090(.A(KEYINPUT9), .B(G234), .Z(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(G217), .A3(new_n202), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n276), .B(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n188), .ZN(new_n280));
  INV_X1    g094(.A(G478), .ZN(new_n281));
  OR2_X1    g095(.A1(new_n281), .A2(KEYINPUT15), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n280), .B(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n249), .A2(new_n257), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G221), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n286), .B1(new_n277), .B2(new_n188), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT85), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT11), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n289), .B1(new_n258), .B2(G137), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n258), .A2(G137), .ZN(new_n291));
  INV_X1    g105(.A(G137), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n292), .A2(KEYINPUT11), .A3(G134), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n290), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G131), .ZN(new_n295));
  INV_X1    g109(.A(G131), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n290), .A2(new_n293), .A3(new_n296), .A4(new_n291), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(KEYINPUT67), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(KEYINPUT67), .B1(new_n295), .B2(new_n297), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G101), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n210), .A2(G107), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n266), .A2(G104), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT3), .B1(new_n210), .B2(G107), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT3), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(new_n266), .A3(G104), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n307), .A2(new_n309), .A3(new_n302), .A4(new_n303), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n310), .A2(KEYINPUT81), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(KEYINPUT81), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n306), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G128), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(KEYINPUT1), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n197), .A2(G143), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n199), .A2(G146), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n199), .B(G146), .C1(new_n314), .C2(KEYINPUT1), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n314), .A2(new_n197), .A3(G143), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n313), .A2(new_n322), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n307), .A2(new_n309), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT81), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n324), .A2(new_n325), .A3(new_n302), .A4(new_n303), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n310), .A2(KEYINPUT81), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n305), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n318), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n321), .A2(KEYINPUT83), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT83), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n319), .A2(new_n331), .A3(new_n320), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n329), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n301), .B1(new_n323), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n288), .B1(new_n335), .B2(KEYINPUT12), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n295), .A2(new_n297), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT67), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n298), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n326), .A2(new_n327), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n341), .A2(new_n306), .A3(new_n333), .ZN(new_n342));
  INV_X1    g156(.A(new_n322), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n343), .B1(new_n341), .B2(new_n306), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n340), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT12), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(KEYINPUT85), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n336), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n323), .A2(new_n334), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n349), .A2(KEYINPUT12), .A3(new_n337), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT84), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n328), .A2(new_n353), .ZN(new_n354));
  AOI211_X1 g168(.A(KEYINPUT84), .B(new_n305), .C1(new_n326), .C2(new_n327), .ZN(new_n355));
  OAI211_X1 g169(.A(KEYINPUT10), .B(new_n343), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n334), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(G143), .B(G146), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT0), .B(G128), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT64), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AND2_X1   g175(.A1(KEYINPUT0), .A2(G128), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n316), .A2(new_n317), .ZN(new_n364));
  NOR2_X1   g178(.A1(KEYINPUT0), .A2(G128), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT64), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n364), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n361), .A2(new_n363), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT66), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT66), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n361), .A2(new_n368), .A3(new_n371), .A4(new_n363), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT82), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n307), .A2(new_n309), .A3(new_n303), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G101), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n374), .B1(new_n376), .B2(KEYINPUT4), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT4), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n375), .A2(KEYINPUT82), .A3(new_n378), .A4(G101), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  OAI211_X1 g194(.A(KEYINPUT4), .B(new_n376), .C1(new_n311), .C2(new_n312), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n373), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n356), .A2(new_n301), .A3(new_n358), .A4(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(G110), .B(G140), .ZN(new_n384));
  INV_X1    g198(.A(G227), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(G953), .ZN(new_n386));
  XOR2_X1   g200(.A(new_n384), .B(new_n386), .Z(new_n387));
  AND2_X1   g201(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n352), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n387), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n382), .A2(new_n358), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n301), .B1(new_n391), .B2(new_n356), .ZN(new_n392));
  INV_X1    g206(.A(new_n383), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n390), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(G902), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT86), .ZN(new_n396));
  INV_X1    g210(.A(G469), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n350), .B1(new_n336), .B2(new_n347), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n383), .A2(new_n387), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n356), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n382), .A2(new_n358), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n340), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n387), .B1(new_n404), .B2(new_n383), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n397), .B(new_n188), .C1(new_n401), .C2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT86), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n398), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n387), .B1(new_n352), .B2(new_n383), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n400), .A2(new_n392), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n188), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G469), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n287), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(G214), .B1(G237), .B2(G902), .ZN(new_n414));
  XOR2_X1   g228(.A(G116), .B(G119), .Z(new_n415));
  XNOR2_X1  g229(.A(KEYINPUT2), .B(G113), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NOR3_X1   g231(.A1(new_n271), .A2(KEYINPUT5), .A3(G119), .ZN(new_n418));
  XNOR2_X1  g232(.A(G116), .B(G119), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n418), .B1(new_n419), .B2(KEYINPUT5), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n417), .B1(G113), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n421), .B1(new_n354), .B2(new_n355), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n419), .B(new_n416), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n381), .A2(new_n380), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT87), .ZN(new_n426));
  XOR2_X1   g240(.A(G110), .B(G122), .Z(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT87), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n381), .A2(new_n380), .A3(new_n429), .A4(new_n424), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n422), .A2(new_n426), .A3(new_n428), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n343), .A2(new_n189), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n432), .B1(new_n369), .B2(new_n189), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n202), .A2(G224), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT7), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n433), .B(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n431), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n427), .B(KEYINPUT8), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT89), .ZN(new_n439));
  AOI211_X1 g253(.A(new_n439), .B(new_n421), .C1(new_n328), .C2(KEYINPUT88), .ZN(new_n440));
  INV_X1    g254(.A(new_n421), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n341), .A2(KEYINPUT88), .A3(new_n306), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n441), .B1(new_n442), .B2(KEYINPUT89), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n328), .A2(new_n439), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n438), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n188), .B1(new_n437), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT90), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n422), .A2(new_n426), .A3(new_n430), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n427), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(KEYINPUT6), .A3(new_n431), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT6), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n449), .A2(new_n452), .A3(new_n427), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n433), .B(new_n434), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT90), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n456), .B(new_n188), .C1(new_n437), .C2(new_n446), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n448), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(G210), .B1(G237), .B2(G902), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT91), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n448), .A2(new_n455), .A3(new_n461), .A4(new_n457), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AND4_X1   g279(.A1(new_n285), .A2(new_n413), .A3(new_n414), .A4(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT32), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT71), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n201), .A2(new_n202), .A3(G210), .ZN(new_n469));
  XOR2_X1   g283(.A(new_n469), .B(KEYINPUT27), .Z(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT26), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(new_n302), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n373), .A2(new_n340), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n292), .A2(G134), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n258), .A2(G137), .ZN(new_n475));
  OAI21_X1  g289(.A(G131), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n297), .A2(new_n476), .A3(KEYINPUT68), .ZN(new_n477));
  AOI21_X1  g291(.A(KEYINPUT68), .B1(new_n297), .B2(new_n476), .ZN(new_n478));
  NOR3_X1   g292(.A1(new_n477), .A2(new_n478), .A3(new_n322), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n473), .A2(new_n423), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT69), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n479), .B1(new_n373), .B2(new_n340), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT69), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n484), .A3(new_n423), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n482), .A2(KEYINPUT28), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT28), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n369), .A2(KEYINPUT65), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT65), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n361), .A2(new_n368), .A3(new_n489), .A4(new_n363), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n488), .A2(new_n337), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n343), .A2(new_n297), .A3(new_n476), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI22_X1  g307(.A1(new_n481), .A2(new_n487), .B1(new_n424), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n472), .B1(new_n486), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(KEYINPUT30), .B1(new_n491), .B2(new_n492), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n497), .B1(KEYINPUT30), .B2(new_n483), .ZN(new_n498));
  AOI22_X1  g312(.A1(new_n498), .A2(new_n424), .B1(new_n482), .B2(new_n485), .ZN(new_n499));
  AOI21_X1  g313(.A(KEYINPUT31), .B1(new_n499), .B2(new_n472), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n482), .A2(new_n485), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT30), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n493), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n473), .A2(KEYINPUT30), .A3(new_n480), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(new_n504), .A3(new_n424), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n501), .A2(KEYINPUT31), .A3(new_n472), .A4(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n496), .B1(new_n500), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(G472), .A2(G902), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(KEYINPUT70), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n468), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n484), .B1(new_n483), .B2(new_n423), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n370), .A2(new_n372), .B1(new_n339), .B2(new_n298), .ZN(new_n514));
  NOR4_X1   g328(.A1(new_n514), .A2(KEYINPUT69), .A3(new_n424), .A4(new_n479), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n505), .B(new_n472), .C1(new_n513), .C2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT31), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n495), .B1(new_n518), .B2(new_n506), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n519), .A2(KEYINPUT71), .A3(new_n510), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n467), .B1(new_n512), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n486), .A2(new_n494), .A3(new_n472), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT29), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT72), .ZN(new_n525));
  AOI211_X1 g339(.A(new_n525), .B(new_n472), .C1(new_n501), .C2(new_n505), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n505), .B1(new_n513), .B2(new_n515), .ZN(new_n527));
  INV_X1    g341(.A(new_n472), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT72), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n524), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n528), .A2(new_n523), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n481), .A2(new_n487), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT74), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT74), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n481), .A2(new_n534), .A3(new_n487), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT73), .B1(new_n483), .B2(new_n423), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT73), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n538), .B(new_n424), .C1(new_n514), .C2(new_n479), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n537), .B(new_n539), .C1(new_n513), .C2(new_n515), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n531), .B(new_n536), .C1(new_n541), .C2(new_n487), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n188), .ZN(new_n543));
  OAI21_X1  g357(.A(G472), .B1(new_n530), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT75), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n519), .A2(new_n467), .A3(new_n510), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(G472), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n525), .B1(new_n499), .B2(new_n472), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n527), .A2(KEYINPUT72), .A3(new_n528), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n550), .A2(new_n523), .A3(new_n551), .A4(new_n522), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n540), .A2(KEYINPUT28), .B1(new_n533), .B2(new_n535), .ZN(new_n553));
  AOI21_X1  g367(.A(G902), .B1(new_n553), .B2(new_n531), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n549), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT75), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n521), .A2(new_n546), .A3(new_n548), .A4(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(G217), .B1(new_n252), .B2(G902), .ZN(new_n558));
  XNOR2_X1  g372(.A(G119), .B(G128), .ZN(new_n559));
  XOR2_X1   g373(.A(KEYINPUT24), .B(G110), .Z(new_n560));
  AOI21_X1  g374(.A(new_n198), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT76), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n559), .A2(new_n562), .A3(KEYINPUT23), .ZN(new_n563));
  OR2_X1    g377(.A1(new_n562), .A2(KEYINPUT23), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(KEYINPUT23), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n564), .A2(G119), .A3(new_n314), .A4(new_n565), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G110), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n561), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n196), .A2(G146), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n567), .A2(G110), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n560), .A2(new_n559), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n570), .B(new_n215), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n202), .A2(G221), .A3(G234), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT79), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(KEYINPUT22), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(G137), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n574), .B(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n188), .ZN(new_n580));
  AND2_X1   g394(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n558), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n579), .A2(new_n188), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(G902), .B1(new_n252), .B2(G217), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n579), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n466), .A2(new_n557), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(G101), .ZN(G3));
  NAND2_X1  g406(.A1(new_n508), .A2(new_n188), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(G472), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n594), .B1(new_n512), .B2(new_n520), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n596), .A2(new_n590), .A3(new_n413), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT33), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n276), .A2(new_n278), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT99), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n278), .B(KEYINPUT98), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n601), .B1(new_n268), .B2(new_n275), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n599), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  OR2_X1    g417(.A1(new_n602), .A2(new_n600), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n598), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n279), .A2(KEYINPUT33), .ZN(new_n606));
  OAI211_X1 g420(.A(G478), .B(new_n188), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n280), .A2(new_n281), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n249), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n458), .A2(new_n459), .ZN(new_n611));
  INV_X1    g425(.A(new_n257), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n448), .A2(new_n455), .A3(new_n460), .A4(new_n457), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n611), .A2(new_n612), .A3(new_n414), .A4(new_n613), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n597), .A2(new_n610), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT34), .B(G104), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G6));
  NAND2_X1  g431(.A1(new_n248), .A2(new_n284), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n597), .A2(new_n614), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT35), .B(G107), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G9));
  INV_X1    g435(.A(KEYINPUT36), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n578), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(new_n574), .B(new_n623), .Z(new_n624));
  AOI22_X1  g438(.A1(new_n582), .A2(new_n585), .B1(new_n587), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n466), .A2(new_n596), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(new_n627), .B(KEYINPUT37), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G110), .ZN(G12));
  AND2_X1   g443(.A1(new_n611), .A2(new_n613), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n630), .A2(new_n626), .A3(new_n414), .ZN(new_n631));
  INV_X1    g445(.A(G900), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n254), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n251), .B(KEYINPUT100), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n618), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n557), .A2(new_n631), .A3(new_n413), .A4(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G128), .ZN(G30));
  OAI21_X1  g452(.A(new_n516), .B1(new_n541), .B2(new_n472), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n639), .A2(new_n188), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n521), .B(new_n548), .C1(new_n549), .C2(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n465), .B(KEYINPUT38), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n248), .A2(new_n283), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n641), .A2(new_n642), .A3(new_n414), .A4(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n635), .B(KEYINPUT39), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n413), .A2(new_n646), .ZN(new_n647));
  OR2_X1    g461(.A1(new_n647), .A2(KEYINPUT40), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n625), .ZN(new_n649));
  AOI211_X1 g463(.A(new_n644), .B(new_n649), .C1(KEYINPUT40), .C2(new_n647), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(new_n199), .ZN(G45));
  INV_X1    g465(.A(new_n635), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n609), .B(new_n652), .C1(new_n240), .C2(new_n247), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n557), .A2(new_n631), .A3(new_n413), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G146), .ZN(G48));
  NOR2_X1   g470(.A1(new_n555), .A2(KEYINPUT75), .ZN(new_n657));
  AOI211_X1 g471(.A(new_n545), .B(new_n549), .C1(new_n552), .C2(new_n554), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n657), .A2(new_n658), .A3(new_n547), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n589), .B1(new_n659), .B2(new_n521), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT102), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n614), .A2(new_n610), .ZN(new_n662));
  INV_X1    g476(.A(new_n287), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n389), .A2(new_n394), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n188), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(G469), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n396), .B1(new_n395), .B2(new_n397), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n406), .A2(KEYINPUT86), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n663), .B(new_n666), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT101), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n408), .A2(new_n671), .A3(new_n663), .A4(new_n666), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n660), .A2(new_n661), .A3(new_n662), .A4(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n673), .A2(new_n557), .A3(new_n590), .A4(new_n662), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(KEYINPUT102), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT41), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G113), .ZN(G15));
  NOR2_X1   g493(.A1(new_n614), .A2(new_n618), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n673), .A2(new_n557), .A3(new_n590), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G116), .ZN(G18));
  INV_X1    g496(.A(new_n669), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n557), .A2(new_n631), .A3(new_n285), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G119), .ZN(G21));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n630), .A2(new_n686), .A3(new_n414), .A4(new_n643), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n643), .A2(new_n611), .A3(new_n414), .A4(new_n613), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(KEYINPUT104), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT103), .B(G472), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n593), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n500), .A2(new_n507), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n553), .A2(new_n472), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n511), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n696), .A2(new_n589), .A3(new_n257), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n690), .A2(new_n673), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G122), .ZN(G24));
  XOR2_X1   g513(.A(new_n653), .B(KEYINPUT105), .Z(new_n700));
  INV_X1    g514(.A(new_n696), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n631), .A2(new_n700), .A3(new_n683), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G125), .ZN(G27));
  OAI21_X1  g517(.A(new_n467), .B1(new_n519), .B2(new_n510), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n546), .A2(new_n548), .A3(new_n556), .A4(new_n704), .ZN(new_n705));
  AOI22_X1  g519(.A1(new_n398), .A2(new_n407), .B1(G469), .B2(new_n411), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n463), .A2(new_n414), .A3(new_n464), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n706), .A2(new_n707), .A3(new_n287), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n705), .A2(new_n708), .A3(new_n700), .A4(new_n590), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT42), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n653), .B(KEYINPUT105), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n711), .A2(KEYINPUT42), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n712), .A2(new_n557), .A3(new_n590), .A4(new_n708), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(new_n296), .ZN(G33));
  NAND4_X1  g529(.A1(new_n557), .A2(new_n590), .A3(new_n636), .A4(new_n708), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G134), .ZN(G36));
  NAND2_X1  g531(.A1(new_n248), .A2(new_n609), .ZN(new_n718));
  XOR2_X1   g532(.A(new_n718), .B(KEYINPUT43), .Z(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n595), .A3(new_n626), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n707), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n720), .A2(new_n721), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(KEYINPUT107), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n409), .A2(new_n410), .ZN(new_n728));
  XOR2_X1   g542(.A(new_n728), .B(KEYINPUT45), .Z(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(G469), .ZN(new_n730));
  NAND2_X1  g544(.A1(G469), .A2(G902), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n730), .A2(KEYINPUT46), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT46), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n733), .B(G469), .C1(new_n729), .C2(G902), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n732), .A2(new_n408), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n663), .A3(new_n646), .ZN(new_n736));
  XOR2_X1   g550(.A(new_n736), .B(KEYINPUT106), .Z(new_n737));
  NAND2_X1  g551(.A1(new_n727), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G137), .ZN(G39));
  NAND2_X1  g553(.A1(new_n735), .A2(new_n663), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT47), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n741), .A2(new_n653), .A3(new_n707), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n557), .A2(new_n590), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G140), .ZN(G42));
  NAND2_X1  g559(.A1(new_n408), .A2(new_n666), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(KEYINPUT49), .ZN(new_n747));
  XOR2_X1   g561(.A(new_n747), .B(KEYINPUT108), .Z(new_n748));
  INV_X1    g562(.A(new_n414), .ZN(new_n749));
  NOR4_X1   g563(.A1(new_n641), .A2(new_n589), .A3(new_n749), .A4(new_n287), .ZN(new_n750));
  INV_X1    g564(.A(new_n642), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n718), .B1(new_n746), .B2(KEYINPUT49), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n748), .A2(new_n750), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT54), .ZN(new_n754));
  INV_X1    g568(.A(new_n708), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n557), .A2(new_n283), .A3(new_n248), .A4(new_n652), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n700), .A2(new_n701), .ZN(new_n757));
  AOI211_X1 g571(.A(new_n625), .B(new_n755), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n710), .A2(new_n713), .A3(new_n716), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n610), .A2(new_n618), .ZN(new_n760));
  AND4_X1   g574(.A1(new_n612), .A2(new_n760), .A3(new_n414), .A4(new_n465), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n761), .A2(new_n596), .A3(new_n590), .A4(new_n413), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n591), .A2(new_n627), .A3(new_n762), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n758), .A2(new_n759), .A3(new_n763), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n681), .A2(new_n698), .A3(new_n684), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n764), .A2(new_n677), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n630), .A2(new_n626), .A3(new_n414), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n767), .B1(new_n659), .B2(new_n521), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n768), .B(new_n413), .C1(new_n636), .C2(new_n654), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n412), .B1(new_n667), .B2(new_n668), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n770), .A2(new_n663), .A3(new_n625), .A4(new_n652), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT110), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT110), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n413), .A2(new_n773), .A3(new_n625), .A4(new_n652), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(new_n641), .A3(new_n690), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n769), .A2(new_n702), .A3(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT113), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n775), .A2(new_n641), .A3(new_n690), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n637), .A2(new_n655), .A3(new_n702), .ZN(new_n781));
  OAI211_X1 g595(.A(KEYINPUT113), .B(new_n778), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n769), .A2(KEYINPUT52), .A3(new_n776), .A4(new_n702), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT111), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n766), .B(KEYINPUT53), .C1(new_n784), .C2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n788), .B1(new_n780), .B2(new_n781), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n785), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT109), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n677), .A2(new_n791), .A3(new_n765), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n791), .B1(new_n677), .B2(new_n765), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n764), .B(new_n790), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n794), .A2(KEYINPUT114), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT114), .B1(new_n794), .B2(new_n795), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n754), .B(new_n787), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n784), .A2(new_n786), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n792), .A2(new_n793), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n799), .A2(new_n795), .A3(new_n800), .A4(new_n764), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n794), .A2(KEYINPUT53), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n798), .B1(new_n803), .B2(new_n754), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  AND4_X1   g619(.A1(new_n590), .A2(new_n719), .A3(new_n634), .A4(new_n701), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n806), .A2(new_n683), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n807), .A2(new_n749), .A3(new_n751), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT50), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n683), .A2(new_n723), .A3(new_n590), .ZN(new_n810));
  INV_X1    g624(.A(new_n251), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n810), .A2(new_n641), .A3(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(new_n248), .A3(new_n608), .A4(new_n607), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n741), .B1(new_n663), .B2(new_n746), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n806), .A2(new_n723), .ZN(new_n816));
  XOR2_X1   g630(.A(new_n816), .B(KEYINPUT115), .Z(new_n817));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  AND4_X1   g632(.A1(new_n634), .A2(new_n719), .A3(new_n683), .A4(new_n723), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n626), .A3(new_n701), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n814), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n814), .A2(KEYINPUT51), .A3(new_n818), .A4(new_n820), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n589), .B1(new_n659), .B2(new_n704), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n819), .A2(new_n825), .ZN(new_n826));
  XOR2_X1   g640(.A(new_n826), .B(KEYINPUT48), .Z(new_n827));
  INV_X1    g641(.A(new_n610), .ZN(new_n828));
  AOI211_X1 g642(.A(new_n250), .B(new_n827), .C1(new_n828), .C2(new_n812), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n823), .A2(new_n824), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n807), .A2(new_n414), .A3(new_n630), .ZN(new_n831));
  XOR2_X1   g645(.A(new_n831), .B(KEYINPUT116), .Z(new_n832));
  AND3_X1   g646(.A1(new_n805), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(G952), .A2(G953), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n753), .B1(new_n833), .B2(new_n834), .ZN(G75));
  XNOR2_X1  g649(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n787), .B1(new_n796), .B2(new_n797), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(G210), .A3(G902), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT56), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n451), .A2(new_n453), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(new_n454), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n839), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n842), .B1(new_n839), .B2(new_n840), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n837), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n839), .A2(new_n840), .ZN(new_n846));
  INV_X1    g660(.A(new_n842), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n839), .A2(new_n840), .A3(new_n842), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n836), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n202), .A2(G952), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n845), .A2(new_n850), .A3(new_n852), .ZN(G51));
  XOR2_X1   g667(.A(new_n731), .B(KEYINPUT118), .Z(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT57), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n854), .A2(KEYINPUT57), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n838), .A2(KEYINPUT54), .ZN(new_n857));
  INV_X1    g671(.A(new_n798), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n855), .B(new_n856), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n664), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n730), .B(KEYINPUT119), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n838), .A2(G902), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n851), .B1(new_n860), .B2(new_n862), .ZN(G54));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT120), .B1(new_n864), .B2(new_n187), .ZN(new_n865));
  OR3_X1    g679(.A1(new_n864), .A2(new_n187), .A3(KEYINPUT120), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n838), .A2(G902), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n238), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n867), .A2(new_n868), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n869), .A2(new_n870), .A3(new_n851), .ZN(G60));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n857), .A2(new_n858), .ZN(new_n873));
  NAND2_X1  g687(.A1(G478), .A2(G902), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT59), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n875), .B1(new_n605), .B2(new_n606), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n872), .B(new_n852), .C1(new_n873), .C2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n804), .A2(new_n875), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n605), .A2(new_n606), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n838), .A2(KEYINPUT54), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n876), .B1(new_n881), .B2(new_n798), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT121), .B1(new_n882), .B2(new_n851), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n877), .A2(new_n880), .A3(new_n883), .ZN(G63));
  NAND2_X1  g698(.A1(G217), .A2(G902), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT60), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n838), .A2(new_n624), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n852), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n579), .B(KEYINPUT122), .Z(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(new_n838), .B2(new_n887), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT61), .ZN(G66));
  AOI21_X1  g708(.A(new_n202), .B1(new_n255), .B2(G224), .ZN(new_n895));
  INV_X1    g709(.A(new_n763), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n800), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n895), .B1(new_n897), .B2(new_n202), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n841), .B1(G898), .B2(new_n202), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n898), .B(new_n899), .Z(G69));
  NAND2_X1  g714(.A1(new_n825), .A2(new_n690), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n726), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n781), .B1(new_n902), .B2(new_n737), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n759), .B1(new_n742), .B2(new_n743), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n903), .A2(new_n202), .A3(new_n904), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n498), .B(new_n226), .Z(new_n906));
  OAI211_X1 g720(.A(new_n905), .B(new_n906), .C1(new_n632), .C2(new_n202), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n650), .A2(new_n781), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT62), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n647), .A2(new_n707), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n660), .A2(new_n760), .A3(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n910), .A2(new_n738), .A3(new_n744), .A4(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n906), .B1(new_n913), .B2(new_n202), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n908), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(G953), .B1(new_n385), .B2(new_n632), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n915), .B(new_n916), .ZN(G72));
  NAND3_X1  g731(.A1(new_n550), .A2(new_n516), .A3(new_n551), .ZN(new_n918));
  NAND2_X1  g732(.A1(G472), .A2(G902), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT63), .Z(new_n920));
  NAND2_X1  g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT125), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n801), .A2(new_n802), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(KEYINPUT126), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n801), .A2(new_n925), .A3(new_n802), .A4(new_n922), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n527), .B(KEYINPUT124), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n903), .A2(new_n800), .A3(new_n896), .A4(new_n904), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n920), .B(KEYINPUT123), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n851), .B1(new_n931), .B2(new_n528), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n930), .B1(new_n913), .B2(new_n897), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n933), .A2(new_n472), .A3(new_n928), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n927), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(KEYINPUT127), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n927), .A2(new_n932), .A3(new_n934), .A4(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n936), .A2(new_n938), .ZN(G57));
endmodule


