//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 0 1 1 1 1 1 0 1 0 0 1 0 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n878, new_n879, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014;
  XNOR2_X1  g000(.A(G71gat), .B(G78gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(KEYINPUT100), .ZN(new_n203));
  AND2_X1   g002(.A1(G71gat), .A2(G78gat), .ZN(new_n204));
  OR2_X1    g003(.A1(new_n204), .A2(KEYINPUT9), .ZN(new_n205));
  XOR2_X1   g004(.A(G57gat), .B(G64gat), .Z(new_n206));
  NAND2_X1  g005(.A1(new_n202), .A2(KEYINPUT100), .ZN(new_n207));
  NAND4_X1  g006(.A1(new_n203), .A2(new_n205), .A3(new_n206), .A4(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT98), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n202), .B(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n205), .A2(new_n206), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AND2_X1   g011(.A1(new_n212), .A2(KEYINPUT99), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(KEYINPUT99), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n208), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT21), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G127gat), .ZN(new_n218));
  INV_X1    g017(.A(G127gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n215), .A2(new_n216), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G15gat), .B(G22gat), .ZN(new_n222));
  OR2_X1    g021(.A1(new_n222), .A2(G1gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n222), .B1(new_n224), .B2(G1gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n225), .A3(KEYINPUT93), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n226), .B(G8gat), .C1(KEYINPUT93), .C2(new_n223), .ZN(new_n227));
  XOR2_X1   g026(.A(KEYINPUT94), .B(G8gat), .Z(new_n228));
  NAND3_X1  g027(.A1(new_n223), .A2(new_n225), .A3(new_n228), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n227), .B(new_n229), .C1(new_n215), .C2(new_n216), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n221), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n234));
  XNOR2_X1  g033(.A(G155gat), .B(G183gat), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n234), .B(new_n235), .Z(new_n236));
  NOR2_X1   g035(.A1(new_n221), .A2(new_n231), .ZN(new_n237));
  OR3_X1    g036(.A1(new_n233), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(G231gat), .A2(G233gat), .ZN(new_n239));
  INV_X1    g038(.A(G211gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n236), .B1(new_n233), .B2(new_n237), .ZN(new_n242));
  AND3_X1   g041(.A1(new_n238), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n241), .B1(new_n238), .B2(new_n242), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G232gat), .A2(G233gat), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n247), .A2(KEYINPUT41), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(G162gat), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G43gat), .B(G50gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(KEYINPUT15), .ZN(new_n252));
  NAND2_X1  g051(.A1(G29gat), .A2(G36gat), .ZN(new_n253));
  OR3_X1    g052(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n252), .B1(new_n253), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT89), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT91), .ZN(new_n260));
  OAI22_X1  g059(.A1(new_n256), .A2(new_n260), .B1(new_n251), .B2(KEYINPUT15), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n254), .A2(KEYINPUT91), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT90), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n252), .B(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n263), .A2(new_n265), .A3(new_n253), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT17), .ZN(new_n268));
  OR2_X1    g067(.A1(new_n268), .A2(KEYINPUT92), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(KEYINPUT92), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n267), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n259), .A2(KEYINPUT92), .A3(new_n266), .A4(new_n268), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G99gat), .ZN(new_n274));
  INV_X1    g073(.A(G106gat), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT101), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT101), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n277), .A2(G99gat), .A3(G106gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n276), .A2(KEYINPUT8), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G85gat), .A2(G92gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT7), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n279), .B(new_n281), .C1(G85gat), .C2(G92gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(G99gat), .B(G106gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n273), .A2(new_n285), .B1(KEYINPUT41), .B2(new_n247), .ZN(new_n286));
  INV_X1    g085(.A(G134gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n267), .A2(new_n284), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n287), .B1(new_n286), .B2(new_n288), .ZN(new_n291));
  XNOR2_X1  g090(.A(G190gat), .B(G218gat), .ZN(new_n292));
  XOR2_X1   g091(.A(new_n292), .B(KEYINPUT102), .Z(new_n293));
  NOR3_X1   g092(.A1(new_n290), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n293), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n286), .A2(new_n288), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G134gat), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n295), .B1(new_n297), .B2(new_n289), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n250), .B1(new_n294), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n293), .B1(new_n290), .B2(new_n291), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n297), .A2(new_n289), .A3(new_n295), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(new_n301), .A3(new_n249), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G230gat), .A2(G233gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n215), .A2(new_n285), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT10), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n284), .B(new_n208), .C1(new_n213), .C2(new_n214), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  OR2_X1    g108(.A1(new_n308), .A2(new_n307), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n305), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G120gat), .B(G148gat), .ZN(new_n312));
  INV_X1    g111(.A(G176gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n312), .B(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G204gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n314), .B(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n304), .B1(new_n306), .B2(new_n308), .ZN(new_n317));
  NOR3_X1   g116(.A1(new_n311), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n318), .B(KEYINPUT103), .ZN(new_n319));
  XOR2_X1   g118(.A(new_n316), .B(KEYINPUT104), .Z(new_n320));
  XNOR2_X1  g119(.A(new_n304), .B(KEYINPUT105), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n321), .B1(new_n309), .B2(new_n310), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n320), .B1(new_n322), .B2(new_n317), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n245), .A2(new_n303), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT68), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n219), .A2(KEYINPUT67), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT67), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G127gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(new_n330), .A3(G134gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n219), .A2(new_n287), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G113gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(G120gat), .ZN(new_n335));
  INV_X1    g134(.A(G120gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G113gat), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT1), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n327), .B1(new_n333), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n335), .A2(new_n337), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT1), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n342), .A2(KEYINPUT68), .A3(new_n332), .A4(new_n331), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(G148gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G141gat), .ZN(new_n346));
  INV_X1    g145(.A(G141gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(G148gat), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT2), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G155gat), .B(G162gat), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT75), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  AND2_X1   g150(.A1(G155gat), .A2(G162gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(G155gat), .A2(G162gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT75), .ZN(new_n355));
  XNOR2_X1  g154(.A(G141gat), .B(G148gat), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n354), .B(new_n355), .C1(new_n356), .C2(KEYINPUT2), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT2), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(G155gat), .ZN(new_n360));
  INV_X1    g159(.A(G162gat), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT76), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n347), .A2(KEYINPUT76), .A3(G148gat), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(new_n346), .A3(new_n365), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n351), .A2(new_n357), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT69), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n335), .A2(new_n337), .A3(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n334), .A2(KEYINPUT69), .A3(G120gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(G127gat), .B(G134gat), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n369), .A2(new_n370), .A3(new_n341), .A4(new_n371), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n344), .A2(new_n367), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n372), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n374), .B1(new_n339), .B2(new_n343), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n375), .A2(new_n367), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(G225gat), .A2(G233gat), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT5), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n366), .A2(new_n362), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n346), .A2(new_n348), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n358), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n355), .B1(new_n382), .B2(new_n354), .ZN(new_n383));
  NOR3_X1   g182(.A1(new_n349), .A2(KEYINPUT75), .A3(new_n350), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n380), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT3), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n344), .A2(new_n372), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n367), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n386), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n344), .A2(new_n367), .A3(new_n372), .ZN(new_n391));
  XNOR2_X1  g190(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n375), .A2(KEYINPUT4), .A3(new_n367), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n390), .A2(new_n393), .A3(new_n378), .A4(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT78), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n378), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n398), .B1(new_n391), .B2(new_n392), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n399), .A2(KEYINPUT78), .A3(new_n390), .A4(new_n394), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n379), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n390), .A2(KEYINPUT4), .A3(new_n391), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n373), .A2(new_n392), .ZN(new_n403));
  AOI211_X1 g202(.A(KEYINPUT5), .B(new_n398), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n405));
  XNOR2_X1  g204(.A(G1gat), .B(G29gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G57gat), .B(G85gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n407), .B(new_n408), .Z(new_n409));
  NOR3_X1   g208(.A1(new_n401), .A2(new_n404), .A3(new_n409), .ZN(new_n410));
  XOR2_X1   g209(.A(KEYINPUT80), .B(KEYINPUT6), .Z(new_n411));
  OAI21_X1  g210(.A(KEYINPUT81), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n379), .ZN(new_n413));
  AOI22_X1  g212(.A1(KEYINPUT3), .A2(new_n385), .B1(new_n344), .B2(new_n372), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n389), .A2(new_n414), .B1(new_n373), .B2(KEYINPUT4), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT78), .B1(new_n415), .B2(new_n399), .ZN(new_n416));
  INV_X1    g215(.A(new_n400), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n413), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n409), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n403), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT5), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(new_n421), .A3(new_n378), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n418), .A2(new_n419), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT81), .ZN(new_n424));
  INV_X1    g223(.A(new_n411), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n409), .B1(new_n401), .B2(new_n404), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n412), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n427), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n411), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(G8gat), .B(G36gat), .ZN(new_n432));
  INV_X1    g231(.A(G64gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  XOR2_X1   g233(.A(new_n434), .B(G92gat), .Z(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(G183gat), .A2(G190gat), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT24), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n440));
  INV_X1    g239(.A(G183gat), .ZN(new_n441));
  INV_X1    g240(.A(G190gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n439), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT64), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n446), .A2(KEYINPUT25), .ZN(new_n447));
  INV_X1    g246(.A(G169gat), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n448), .A2(new_n313), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT23), .ZN(new_n450));
  NOR3_X1   g249(.A1(new_n450), .A2(G169gat), .A3(G176gat), .ZN(new_n451));
  NOR2_X1   g250(.A1(G169gat), .A2(G176gat), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT65), .B1(new_n452), .B2(KEYINPUT23), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT65), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n454), .B(new_n450), .C1(G169gat), .C2(G176gat), .ZN(new_n455));
  AOI211_X1 g254(.A(new_n449), .B(new_n451), .C1(new_n453), .C2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n444), .A2(new_n445), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n447), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n441), .A2(KEYINPUT66), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT66), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(G183gat), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n461), .A3(KEYINPUT27), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n462), .B1(KEYINPUT27), .B2(G183gat), .ZN(new_n463));
  NOR2_X1   g262(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n437), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n452), .B(KEYINPUT26), .ZN(new_n467));
  INV_X1    g266(.A(new_n449), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  XOR2_X1   g268(.A(KEYINPUT27), .B(G183gat), .Z(new_n470));
  OAI21_X1  g269(.A(KEYINPUT28), .B1(new_n470), .B2(G190gat), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n465), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n453), .A2(new_n455), .ZN(new_n473));
  INV_X1    g272(.A(new_n451), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(new_n474), .A3(new_n468), .ZN(new_n475));
  AOI21_X1  g274(.A(G190gat), .B1(new_n459), .B2(new_n461), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n439), .A2(new_n440), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT25), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n458), .A2(new_n472), .A3(new_n479), .ZN(new_n480));
  AND2_X1   g279(.A1(G226gat), .A2(G233gat), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT29), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n458), .A2(new_n472), .A3(new_n479), .A4(new_n482), .ZN(new_n486));
  XNOR2_X1  g285(.A(KEYINPUT73), .B(G211gat), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT22), .B1(new_n487), .B2(G218gat), .ZN(new_n488));
  XOR2_X1   g287(.A(G197gat), .B(G204gat), .Z(new_n489));
  XNOR2_X1  g288(.A(G211gat), .B(G218gat), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT74), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(G218gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(G211gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n240), .A2(G218gat), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n494), .A2(new_n495), .A3(new_n491), .ZN(new_n496));
  OAI22_X1  g295(.A1(new_n488), .A2(new_n489), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n240), .A2(KEYINPUT73), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT73), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(G211gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(new_n500), .A3(G218gat), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT22), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n489), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n494), .A2(new_n495), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT74), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n503), .A2(new_n504), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n497), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n485), .A2(new_n486), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n509), .B1(new_n485), .B2(new_n486), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n436), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n485), .A2(new_n486), .ZN(new_n514));
  INV_X1    g313(.A(new_n509), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n516), .A2(new_n510), .A3(new_n435), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n513), .A2(new_n517), .A3(KEYINPUT30), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT30), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n519), .B(new_n436), .C1(new_n511), .C2(new_n512), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n431), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(G228gat), .A2(G233gat), .ZN(new_n523));
  XOR2_X1   g322(.A(new_n523), .B(KEYINPUT83), .Z(new_n524));
  AOI22_X1  g323(.A1(new_n389), .A2(new_n483), .B1(new_n508), .B2(new_n497), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n497), .A2(new_n508), .A3(new_n483), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n367), .B1(new_n526), .B2(new_n388), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n524), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT84), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OR3_X1    g329(.A1(new_n525), .A2(new_n527), .A3(new_n523), .ZN(new_n531));
  OAI211_X1 g330(.A(KEYINPUT84), .B(new_n524), .C1(new_n525), .C2(new_n527), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G78gat), .B(G106gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(G22gat), .B(G50gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n538));
  INV_X1    g337(.A(new_n536), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n530), .A2(new_n531), .A3(new_n539), .A4(new_n532), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n537), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n538), .B1(new_n537), .B2(new_n540), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n522), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT34), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n480), .A2(new_n375), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n387), .A2(new_n479), .A3(new_n458), .A4(new_n472), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(G227gat), .ZN(new_n549));
  INV_X1    g348(.A(G233gat), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n545), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  AOI211_X1 g352(.A(KEYINPUT34), .B(new_n551), .C1(new_n546), .C2(new_n547), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n546), .A2(new_n547), .A3(new_n551), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT32), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT33), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(KEYINPUT70), .B(G71gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(G99gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(G15gat), .B(G43gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n557), .A2(new_n559), .A3(new_n564), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n556), .B(KEYINPUT32), .C1(new_n558), .C2(new_n563), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n555), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT72), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n565), .A2(new_n566), .ZN(new_n570));
  INV_X1    g369(.A(new_n555), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n555), .A2(new_n565), .A3(KEYINPUT72), .A4(new_n566), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n569), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT36), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n570), .A2(KEYINPUT71), .A3(new_n555), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n555), .B1(new_n570), .B2(KEYINPUT71), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT36), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n410), .A2(new_n411), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT86), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n418), .A2(new_n422), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n582), .B1(new_n583), .B2(new_n409), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n582), .B(new_n409), .C1(new_n401), .C2(new_n404), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n581), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NOR3_X1   g386(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT37), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT37), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n589), .B1(new_n516), .B2(new_n510), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n435), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT38), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT37), .B1(new_n511), .B2(new_n512), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n516), .A2(new_n510), .A3(new_n589), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT38), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n595), .A2(new_n596), .A3(new_n435), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n592), .A2(new_n513), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n587), .A2(new_n598), .A3(new_n430), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n427), .A2(KEYINPUT86), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n402), .A2(new_n398), .A3(new_n403), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n377), .A2(new_n378), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n601), .A2(KEYINPUT39), .A3(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(KEYINPUT85), .B(KEYINPUT39), .Z(new_n604));
  NAND4_X1  g403(.A1(new_n402), .A2(new_n398), .A3(new_n403), .A4(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n603), .A2(new_n419), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT40), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT40), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n603), .A2(new_n608), .A3(new_n419), .A4(new_n605), .ZN(new_n609));
  AOI22_X1  g408(.A1(new_n600), .A2(new_n585), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n521), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n543), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT87), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n599), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n613), .B1(new_n599), .B2(new_n612), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n544), .B(new_n580), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n577), .A2(new_n578), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n617), .A2(new_n543), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n431), .A2(new_n618), .A3(new_n521), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(KEYINPUT35), .ZN(new_n620));
  AOI21_X1  g419(.A(KEYINPUT35), .B1(new_n587), .B2(new_n430), .ZN(new_n621));
  NOR3_X1   g420(.A1(new_n543), .A2(new_n574), .A3(new_n611), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n616), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G113gat), .B(G141gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(G197gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT11), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(new_n448), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT95), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n631), .A2(KEYINPUT18), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n227), .A2(new_n229), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n634), .B1(new_n271), .B2(new_n272), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n267), .A2(new_n634), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G229gat), .A2(G233gat), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n633), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OR3_X1    g439(.A1(new_n267), .A2(KEYINPUT96), .A3(new_n634), .ZN(new_n641));
  OAI21_X1  g440(.A(KEYINPUT96), .B1(new_n267), .B2(new_n634), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n641), .A2(new_n636), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n639), .B(KEYINPUT13), .Z(new_n644));
  AND2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n639), .ZN(new_n646));
  NOR4_X1   g445(.A1(new_n635), .A2(new_n646), .A3(new_n637), .A4(new_n632), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n640), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT88), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n630), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n638), .A2(new_n639), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(new_n632), .ZN(new_n652));
  INV_X1    g451(.A(new_n645), .ZN(new_n653));
  INV_X1    g452(.A(new_n647), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n630), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n655), .A2(KEYINPUT88), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n650), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n625), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(KEYINPUT97), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT97), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n625), .A2(new_n661), .A3(new_n658), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n326), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n431), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g465(.A1(new_n663), .A2(new_n611), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(G8gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT106), .ZN(new_n669));
  NOR2_X1   g468(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n670));
  AND2_X1   g469(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT42), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n672), .A2(new_n673), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n669), .B1(new_n674), .B2(new_n675), .ZN(G1325gat));
  INV_X1    g475(.A(new_n574), .ZN(new_n677));
  AOI21_X1  g476(.A(G15gat), .B1(new_n663), .B2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT107), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n576), .A2(new_n679), .A3(new_n579), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n679), .B1(new_n576), .B2(new_n579), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n683), .A2(G15gat), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n678), .B1(new_n663), .B2(new_n684), .ZN(G1326gat));
  INV_X1    g484(.A(G22gat), .ZN(new_n686));
  INV_X1    g485(.A(new_n326), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n661), .B1(new_n625), .B2(new_n658), .ZN(new_n688));
  INV_X1    g487(.A(new_n658), .ZN(new_n689));
  AOI211_X1 g488(.A(KEYINPUT97), .B(new_n689), .C1(new_n616), .C2(new_n624), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n543), .B(new_n687), .C1(new_n688), .C2(new_n690), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n691), .A2(KEYINPUT108), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(KEYINPUT108), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n693), .B1(new_n692), .B2(new_n694), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n686), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n692), .A2(new_n694), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(KEYINPUT43), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n692), .A2(new_n694), .A3(new_n693), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n699), .A2(G22gat), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n697), .A2(new_n701), .ZN(G1327gat));
  OAI211_X1 g501(.A(new_n682), .B(new_n544), .C1(new_n614), .C2(new_n615), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n624), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n299), .A2(new_n302), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT44), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707));
  AOI211_X1 g506(.A(new_n707), .B(new_n303), .C1(new_n616), .C2(new_n624), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n245), .A2(new_n324), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n689), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(G29gat), .B1(new_n713), .B2(new_n431), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n660), .A2(new_n662), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n711), .A2(new_n303), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n718));
  INV_X1    g517(.A(G29gat), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n717), .A2(new_n718), .A3(new_n719), .A4(new_n664), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT45), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n715), .A2(new_n719), .A3(new_n716), .ZN(new_n722));
  OAI21_X1  g521(.A(KEYINPUT109), .B1(new_n722), .B2(new_n431), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n720), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n721), .B1(new_n720), .B2(new_n723), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n714), .B1(new_n724), .B2(new_n725), .ZN(G1328gat));
  INV_X1    g525(.A(G36gat), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n717), .A2(new_n727), .ZN(new_n728));
  OR3_X1    g527(.A1(new_n728), .A2(KEYINPUT46), .A3(new_n521), .ZN(new_n729));
  OAI21_X1  g528(.A(G36gat), .B1(new_n713), .B2(new_n521), .ZN(new_n730));
  OAI21_X1  g529(.A(KEYINPUT46), .B1(new_n728), .B2(new_n521), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(G1329gat));
  AOI22_X1  g531(.A1(new_n619), .A2(KEYINPUT35), .B1(new_n622), .B2(new_n621), .ZN(new_n733));
  INV_X1    g532(.A(new_n543), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n734), .B1(new_n431), .B2(new_n521), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n423), .A2(new_n425), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n736), .B1(new_n600), .B2(new_n585), .ZN(new_n737));
  INV_X1    g536(.A(new_n430), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n592), .A2(new_n513), .A3(new_n597), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n607), .A2(new_n609), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n741), .B(new_n611), .C1(new_n584), .C2(new_n586), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n734), .ZN(new_n743));
  OAI21_X1  g542(.A(KEYINPUT87), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n599), .A2(new_n612), .A3(new_n613), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n735), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n733), .B1(new_n746), .B2(new_n682), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n707), .B1(new_n747), .B2(new_n303), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n625), .A2(KEYINPUT44), .A3(new_n705), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n748), .A2(new_n683), .A3(new_n712), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G43gat), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n574), .A2(G43gat), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n716), .B(new_n752), .C1(new_n688), .C2(new_n690), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n751), .A2(KEYINPUT47), .A3(new_n753), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n715), .A2(KEYINPUT110), .A3(new_n716), .A4(new_n752), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n755), .A2(new_n757), .A3(new_n751), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT47), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n759), .B1(new_n758), .B2(new_n760), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n754), .B1(new_n761), .B2(new_n762), .ZN(G1330gat));
  NOR2_X1   g562(.A1(new_n734), .A2(G50gat), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n748), .A2(new_n543), .A3(new_n712), .A4(new_n749), .ZN(new_n765));
  AOI22_X1  g564(.A1(new_n717), .A2(new_n764), .B1(G50gat), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(KEYINPUT112), .B1(new_n765), .B2(G50gat), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT48), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n766), .B(new_n769), .ZN(G1331gat));
  INV_X1    g569(.A(new_n245), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n747), .A2(new_n771), .A3(new_n705), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n325), .A2(new_n658), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n664), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G57gat), .ZN(G1332gat));
  AND2_X1   g575(.A1(new_n774), .A2(new_n611), .ZN(new_n777));
  NOR2_X1   g576(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n778));
  AND2_X1   g577(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n780), .B1(new_n777), .B2(new_n778), .ZN(G1333gat));
  AOI21_X1  g580(.A(G71gat), .B1(new_n774), .B2(new_n677), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n683), .A2(G71gat), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n774), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n784), .B(new_n785), .ZN(G1334gat));
  NAND2_X1  g585(.A1(new_n774), .A2(new_n543), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g587(.A(new_n303), .B1(new_n703), .B2(new_n624), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n245), .A2(new_n658), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n789), .A2(KEYINPUT51), .A3(new_n790), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(G85gat), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n325), .A2(new_n431), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n709), .A2(new_n797), .A3(new_n790), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n799), .B2(new_n796), .ZN(G1336gat));
  NAND4_X1  g599(.A1(new_n748), .A2(new_n324), .A3(new_n749), .A4(new_n790), .ZN(new_n801));
  OAI21_X1  g600(.A(G92gat), .B1(new_n801), .B2(new_n521), .ZN(new_n802));
  INV_X1    g601(.A(new_n795), .ZN(new_n803));
  OR3_X1    g602(.A1(new_n325), .A2(new_n521), .A3(G92gat), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n805), .A2(KEYINPUT113), .A3(new_n806), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n806), .A2(KEYINPUT113), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n806), .A2(KEYINPUT113), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n805), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n807), .A2(new_n810), .ZN(G1337gat));
  OAI21_X1  g610(.A(G99gat), .B1(new_n801), .B2(new_n682), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n324), .A2(new_n677), .A3(new_n274), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n812), .B1(new_n803), .B2(new_n813), .ZN(G1338gat));
  OAI21_X1  g613(.A(G106gat), .B1(new_n801), .B2(new_n734), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n325), .A2(G106gat), .A3(new_n734), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n795), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(KEYINPUT115), .A3(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n816), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n822), .B1(new_n793), .B2(new_n794), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n709), .A2(new_n543), .A3(new_n324), .A4(new_n790), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n823), .B1(new_n824), .B2(G106gat), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT114), .B1(new_n825), .B2(KEYINPUT115), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n815), .A2(KEYINPUT114), .A3(new_n817), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT53), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n821), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(G1339gat));
  NAND3_X1  g629(.A1(new_n309), .A2(new_n310), .A3(new_n321), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n309), .A2(new_n310), .ZN(new_n832));
  OAI211_X1 g631(.A(KEYINPUT54), .B(new_n831), .C1(new_n832), .C2(new_n305), .ZN(new_n833));
  INV_X1    g632(.A(new_n316), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n834), .B1(new_n322), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT55), .ZN(new_n838));
  OAI21_X1  g637(.A(KEYINPUT116), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n833), .A2(new_n836), .A3(new_n840), .A4(KEYINPUT55), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n839), .A2(new_n319), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n648), .A2(new_n630), .ZN(new_n843));
  OAI21_X1  g642(.A(KEYINPUT117), .B1(new_n638), .B2(new_n639), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n845), .B(new_n646), .C1(new_n635), .C2(new_n637), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n844), .B(new_n846), .C1(new_n644), .C2(new_n643), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n629), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n837), .A2(new_n838), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n843), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n303), .A2(new_n842), .A3(new_n850), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n843), .A2(new_n848), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n324), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n658), .A2(new_n849), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n853), .B1(new_n854), .B2(new_n842), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n851), .B1(new_n855), .B2(new_n303), .ZN(new_n856));
  OAI22_X1  g655(.A1(new_n856), .A2(new_n245), .B1(new_n658), .B2(new_n326), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(new_n664), .A3(new_n622), .ZN(new_n858));
  OAI21_X1  g657(.A(G113gat), .B1(new_n858), .B2(new_n689), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n326), .A2(new_n658), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n839), .A2(new_n319), .A3(new_n841), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n705), .A2(new_n861), .A3(new_n852), .A4(new_n849), .ZN(new_n862));
  AOI22_X1  g661(.A1(new_n650), .A2(new_n657), .B1(new_n838), .B2(new_n837), .ZN(new_n863));
  AOI22_X1  g662(.A1(new_n863), .A2(new_n861), .B1(new_n324), .B2(new_n852), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n862), .B1(new_n864), .B2(new_n705), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n860), .B1(new_n865), .B2(new_n771), .ZN(new_n866));
  INV_X1    g665(.A(new_n618), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n866), .A2(new_n431), .A3(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n869), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(new_n521), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n658), .A2(new_n334), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n859), .B1(new_n872), .B2(new_n873), .ZN(G1340gat));
  OAI21_X1  g673(.A(G120gat), .B1(new_n858), .B2(new_n325), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n324), .A2(new_n336), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n872), .B2(new_n876), .ZN(G1341gat));
  NAND2_X1  g676(.A1(new_n328), .A2(new_n330), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n858), .A2(new_n878), .A3(new_n771), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n872), .A2(new_n771), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(new_n880), .B2(new_n878), .ZN(G1342gat));
  NAND4_X1  g680(.A1(new_n870), .A2(new_n521), .A3(new_n705), .A4(new_n871), .ZN(new_n882));
  OR3_X1    g681(.A1(new_n882), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n883));
  OAI21_X1  g682(.A(G134gat), .B1(new_n858), .B2(new_n303), .ZN(new_n884));
  OAI21_X1  g683(.A(KEYINPUT56), .B1(new_n882), .B2(G134gat), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(G1343gat));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n648), .A2(new_n649), .A3(new_n630), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n656), .B1(new_n655), .B2(KEYINPUT88), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n890), .B1(new_n833), .B2(new_n836), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n838), .B1(new_n837), .B2(KEYINPUT119), .ZN(new_n892));
  OAI22_X1  g691(.A1(new_n888), .A2(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n853), .B(new_n887), .C1(new_n893), .C2(new_n842), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n303), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n892), .A2(new_n891), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n861), .A2(new_n896), .A3(new_n658), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n887), .B1(new_n897), .B2(new_n853), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n862), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n860), .B1(new_n899), .B2(new_n771), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT57), .B1(new_n900), .B2(new_n734), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n866), .A2(new_n734), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT57), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n683), .A2(new_n431), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n906), .A2(new_n611), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n901), .A2(new_n904), .A3(new_n658), .A4(new_n907), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n908), .A2(G141gat), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n902), .A2(new_n905), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT121), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n689), .A2(G141gat), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n902), .A2(KEYINPUT121), .A3(new_n905), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n912), .A2(new_n521), .A3(new_n913), .A4(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT58), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n902), .A2(new_n907), .A3(new_n913), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n918), .B1(new_n908), .B2(G141gat), .ZN(new_n919));
  OAI22_X1  g718(.A1(new_n909), .A2(new_n917), .B1(new_n919), .B2(new_n916), .ZN(G1344gat));
  NAND4_X1  g719(.A1(new_n912), .A2(new_n521), .A3(new_n324), .A4(new_n914), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n921), .A2(KEYINPUT59), .A3(new_n345), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n903), .B1(new_n900), .B2(new_n734), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n902), .A2(KEYINPUT57), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n325), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(KEYINPUT59), .A3(new_n907), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n901), .A2(new_n904), .A3(new_n907), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n927), .A2(new_n325), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n926), .B1(new_n928), .B2(KEYINPUT59), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n922), .B1(new_n929), .B2(G148gat), .ZN(G1345gat));
  AND2_X1   g729(.A1(new_n912), .A2(new_n914), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n931), .A2(new_n521), .A3(new_n245), .ZN(new_n932));
  INV_X1    g731(.A(new_n927), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n245), .A2(G155gat), .ZN(new_n934));
  XOR2_X1   g733(.A(new_n934), .B(KEYINPUT122), .Z(new_n935));
  AOI22_X1  g734(.A1(new_n932), .A2(new_n360), .B1(new_n933), .B2(new_n935), .ZN(G1346gat));
  OAI21_X1  g735(.A(G162gat), .B1(new_n927), .B2(new_n303), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n931), .A2(new_n361), .A3(new_n521), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n938), .B2(new_n303), .ZN(G1347gat));
  NOR3_X1   g738(.A1(new_n867), .A2(KEYINPUT123), .A3(new_n521), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n866), .A2(new_n664), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(KEYINPUT123), .B1(new_n867), .B2(new_n521), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n944), .A2(new_n448), .A3(new_n658), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n866), .A2(new_n664), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n543), .A2(new_n574), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n946), .A2(KEYINPUT124), .A3(new_n611), .A4(new_n947), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n857), .A2(new_n431), .A3(new_n611), .A4(new_n947), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT124), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n952), .A2(new_n658), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n945), .B1(new_n953), .B2(new_n448), .ZN(G1348gat));
  AOI21_X1  g753(.A(G176gat), .B1(new_n944), .B2(new_n324), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n325), .A2(new_n313), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n955), .B1(new_n952), .B2(new_n956), .ZN(G1349gat));
  NAND3_X1  g756(.A1(new_n948), .A2(new_n951), .A3(new_n245), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n958), .A2(new_n459), .A3(new_n461), .ZN(new_n959));
  OR3_X1    g758(.A1(new_n943), .A2(new_n470), .A3(new_n771), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(KEYINPUT60), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT60), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n959), .A2(new_n963), .A3(new_n960), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n962), .A2(new_n964), .ZN(G1350gat));
  NAND3_X1  g764(.A1(new_n948), .A2(new_n951), .A3(new_n705), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(G190gat), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(KEYINPUT125), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT125), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n966), .A2(new_n969), .A3(G190gat), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n968), .A2(KEYINPUT61), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n944), .A2(new_n442), .A3(new_n705), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT61), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n967), .A2(KEYINPUT125), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n971), .A2(new_n972), .A3(new_n974), .ZN(G1351gat));
  NAND3_X1  g774(.A1(new_n682), .A2(new_n431), .A3(new_n611), .ZN(new_n976));
  NOR3_X1   g775(.A1(new_n866), .A2(new_n734), .A3(new_n976), .ZN(new_n977));
  INV_X1    g776(.A(G197gat), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n977), .A2(new_n978), .A3(new_n658), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n976), .B1(new_n923), .B2(new_n924), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n980), .A2(new_n658), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n979), .B1(new_n981), .B2(new_n978), .ZN(G1352gat));
  INV_X1    g781(.A(KEYINPUT127), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT62), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT126), .ZN(new_n985));
  NOR4_X1   g784(.A1(new_n866), .A2(G204gat), .A3(new_n734), .A4(new_n976), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n985), .B1(new_n986), .B2(new_n324), .ZN(new_n987));
  INV_X1    g786(.A(new_n976), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n857), .A2(new_n315), .A3(new_n543), .A4(new_n988), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n989), .A2(KEYINPUT126), .A3(new_n325), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n984), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g790(.A(KEYINPUT126), .B1(new_n989), .B2(new_n325), .ZN(new_n992));
  NAND4_X1  g791(.A1(new_n977), .A2(new_n985), .A3(new_n315), .A4(new_n324), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n992), .A2(new_n993), .A3(KEYINPUT62), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n315), .B1(new_n925), .B2(new_n988), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n983), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AND3_X1   g796(.A1(new_n992), .A2(new_n993), .A3(KEYINPUT62), .ZN(new_n998));
  AOI21_X1  g797(.A(KEYINPUT62), .B1(new_n992), .B2(new_n993), .ZN(new_n999));
  NOR2_X1   g798(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n923), .A2(new_n924), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n1001), .A2(new_n324), .A3(new_n988), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1002), .A2(G204gat), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n1000), .A2(new_n1003), .A3(KEYINPUT127), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n997), .A2(new_n1004), .ZN(G1353gat));
  NOR2_X1   g804(.A1(new_n771), .A2(new_n487), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n977), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n980), .A2(new_n245), .ZN(new_n1008));
  AOI21_X1  g807(.A(KEYINPUT63), .B1(new_n1008), .B2(G211gat), .ZN(new_n1009));
  INV_X1    g808(.A(KEYINPUT63), .ZN(new_n1010));
  AOI211_X1 g809(.A(new_n1010), .B(new_n240), .C1(new_n980), .C2(new_n245), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n1007), .B1(new_n1009), .B2(new_n1011), .ZN(G1354gat));
  AOI21_X1  g811(.A(G218gat), .B1(new_n977), .B2(new_n705), .ZN(new_n1013));
  NOR2_X1   g812(.A1(new_n303), .A2(new_n493), .ZN(new_n1014));
  AOI21_X1  g813(.A(new_n1013), .B1(new_n980), .B2(new_n1014), .ZN(G1355gat));
endmodule


