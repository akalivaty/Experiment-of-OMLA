

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594;

  XNOR2_X1 U322 ( .A(n324), .B(n323), .ZN(n430) );
  XNOR2_X1 U323 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U324 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U325 ( .A(n380), .B(n379), .Z(n530) );
  XNOR2_X1 U326 ( .A(n375), .B(n374), .ZN(n377) );
  XOR2_X1 U327 ( .A(n374), .B(n365), .Z(n526) );
  XOR2_X1 U328 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n290) );
  XOR2_X1 U329 ( .A(n290), .B(n318), .Z(n291) );
  AND2_X1 U330 ( .A1(G230GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U331 ( .A(n434), .B(n433), .ZN(n470) );
  NOR2_X1 U332 ( .A1(n544), .A2(n467), .ZN(n468) );
  XNOR2_X1 U333 ( .A(n423), .B(n292), .ZN(n424) );
  XNOR2_X1 U334 ( .A(n484), .B(KEYINPUT55), .ZN(n485) );
  XNOR2_X1 U335 ( .A(n425), .B(n424), .ZN(n427) );
  INV_X1 U336 ( .A(KEYINPUT54), .ZN(n480) );
  XNOR2_X1 U337 ( .A(n291), .B(n430), .ZN(n327) );
  NOR2_X1 U338 ( .A1(n412), .A2(n411), .ZN(n496) );
  XNOR2_X1 U339 ( .A(n373), .B(n372), .ZN(n375) );
  INV_X1 U340 ( .A(KEYINPUT36), .ZN(n333) );
  INV_X1 U341 ( .A(KEYINPUT101), .ZN(n453) );
  XNOR2_X1 U342 ( .A(n464), .B(n333), .ZN(n334) );
  NOR2_X1 U343 ( .A1(n543), .A2(n488), .ZN(n489) );
  XNOR2_X1 U344 ( .A(n453), .B(KEYINPUT38), .ZN(n454) );
  XNOR2_X1 U345 ( .A(n566), .B(n334), .ZN(n592) );
  XOR2_X1 U346 ( .A(KEYINPUT120), .B(n489), .Z(n574) );
  INV_X1 U347 ( .A(G43GAT), .ZN(n460) );
  XNOR2_X1 U348 ( .A(n455), .B(n454), .ZN(n510) );
  XNOR2_X1 U349 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U350 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U351 ( .A(n494), .B(n493), .ZN(G1351GAT) );
  XNOR2_X1 U352 ( .A(n463), .B(n462), .ZN(G1330GAT) );
  XOR2_X1 U353 ( .A(KEYINPUT81), .B(KEYINPUT0), .Z(n294) );
  XNOR2_X1 U354 ( .A(G113GAT), .B(G134GAT), .ZN(n293) );
  XNOR2_X1 U355 ( .A(n294), .B(n293), .ZN(n378) );
  XOR2_X1 U356 ( .A(n378), .B(G1GAT), .Z(n296) );
  NAND2_X1 U357 ( .A1(G225GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U358 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U359 ( .A(KEYINPUT92), .B(KEYINPUT5), .Z(n298) );
  XNOR2_X1 U360 ( .A(KEYINPUT1), .B(G57GAT), .ZN(n297) );
  XNOR2_X1 U361 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U362 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U363 ( .A(KEYINPUT6), .B(G155GAT), .Z(n302) );
  XNOR2_X1 U364 ( .A(G127GAT), .B(G148GAT), .ZN(n301) );
  XNOR2_X1 U365 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U366 ( .A(n304), .B(n303), .ZN(n309) );
  XNOR2_X1 U367 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n305) );
  XNOR2_X1 U368 ( .A(n305), .B(KEYINPUT2), .ZN(n389) );
  XOR2_X1 U369 ( .A(G85GAT), .B(n389), .Z(n307) );
  XNOR2_X1 U370 ( .A(G120GAT), .B(G162GAT), .ZN(n306) );
  XNOR2_X1 U371 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U372 ( .A(n309), .B(n308), .Z(n314) );
  XOR2_X1 U373 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n311) );
  XNOR2_X1 U374 ( .A(KEYINPUT89), .B(KEYINPUT4), .ZN(n310) );
  XNOR2_X1 U375 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U376 ( .A(G29GAT), .B(n312), .ZN(n313) );
  XNOR2_X1 U377 ( .A(n314), .B(n313), .ZN(n524) );
  XOR2_X1 U378 ( .A(KEYINPUT69), .B(KEYINPUT7), .Z(n316) );
  XNOR2_X1 U379 ( .A(G43GAT), .B(G29GAT), .ZN(n315) );
  XNOR2_X1 U380 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U381 ( .A(KEYINPUT8), .B(n317), .Z(n447) );
  NAND2_X1 U382 ( .A1(G232GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U383 ( .A(G99GAT), .B(G106GAT), .ZN(n324) );
  INV_X1 U384 ( .A(G85GAT), .ZN(n319) );
  NAND2_X1 U385 ( .A1(G92GAT), .A2(n319), .ZN(n322) );
  INV_X1 U386 ( .A(G92GAT), .ZN(n320) );
  NAND2_X1 U387 ( .A1(n320), .A2(G85GAT), .ZN(n321) );
  NAND2_X1 U388 ( .A1(n322), .A2(n321), .ZN(n323) );
  XNOR2_X1 U389 ( .A(G36GAT), .B(G190GAT), .ZN(n325) );
  XNOR2_X1 U390 ( .A(n325), .B(G218GAT), .ZN(n355) );
  XNOR2_X1 U391 ( .A(G134GAT), .B(n355), .ZN(n326) );
  XNOR2_X1 U392 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U393 ( .A(G50GAT), .B(G162GAT), .Z(n390) );
  XNOR2_X1 U394 ( .A(n390), .B(KEYINPUT11), .ZN(n329) );
  INV_X1 U395 ( .A(KEYINPUT65), .ZN(n328) );
  XNOR2_X1 U396 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U397 ( .A(n447), .B(n332), .ZN(n566) );
  INV_X1 U398 ( .A(KEYINPUT78), .ZN(n464) );
  XOR2_X1 U399 ( .A(G211GAT), .B(G78GAT), .Z(n336) );
  XNOR2_X1 U400 ( .A(G183GAT), .B(G71GAT), .ZN(n335) );
  XNOR2_X1 U401 ( .A(n336), .B(n335), .ZN(n349) );
  XOR2_X1 U402 ( .A(G22GAT), .B(G155GAT), .Z(n386) );
  XOR2_X1 U403 ( .A(G15GAT), .B(G127GAT), .Z(n376) );
  XOR2_X1 U404 ( .A(n386), .B(n376), .Z(n338) );
  NAND2_X1 U405 ( .A1(G231GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U406 ( .A(n338), .B(n337), .ZN(n342) );
  XNOR2_X1 U407 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n339) );
  XNOR2_X1 U408 ( .A(n339), .B(KEYINPUT70), .ZN(n428) );
  XNOR2_X1 U409 ( .A(n428), .B(KEYINPUT14), .ZN(n340) );
  XNOR2_X1 U410 ( .A(n340), .B(KEYINPUT12), .ZN(n341) );
  XOR2_X1 U411 ( .A(n342), .B(n341), .Z(n347) );
  XOR2_X1 U412 ( .A(G1GAT), .B(G8GAT), .Z(n440) );
  XOR2_X1 U413 ( .A(KEYINPUT79), .B(KEYINPUT15), .Z(n344) );
  XNOR2_X1 U414 ( .A(G64GAT), .B(KEYINPUT80), .ZN(n343) );
  XNOR2_X1 U415 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U416 ( .A(n440), .B(n345), .ZN(n346) );
  XNOR2_X1 U417 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U418 ( .A(n349), .B(n348), .Z(n549) );
  XNOR2_X1 U419 ( .A(KEYINPUT27), .B(KEYINPUT95), .ZN(n366) );
  XNOR2_X1 U420 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n350) );
  XNOR2_X1 U421 ( .A(n350), .B(KEYINPUT18), .ZN(n351) );
  XOR2_X1 U422 ( .A(n351), .B(KEYINPUT83), .Z(n353) );
  XNOR2_X1 U423 ( .A(G169GAT), .B(G183GAT), .ZN(n352) );
  XNOR2_X1 U424 ( .A(n353), .B(n352), .ZN(n374) );
  XNOR2_X1 U425 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n354) );
  XNOR2_X1 U426 ( .A(n354), .B(G211GAT), .ZN(n397) );
  XNOR2_X1 U427 ( .A(G8GAT), .B(n397), .ZN(n361) );
  INV_X1 U428 ( .A(n355), .ZN(n359) );
  XOR2_X1 U429 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n357) );
  NAND2_X1 U430 ( .A1(G226GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U431 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U432 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U433 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U434 ( .A(G176GAT), .B(G64GAT), .Z(n417) );
  XOR2_X1 U435 ( .A(n362), .B(n417), .Z(n364) );
  XNOR2_X1 U436 ( .A(G204GAT), .B(G92GAT), .ZN(n363) );
  XNOR2_X1 U437 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U438 ( .A(n366), .B(n526), .Z(n407) );
  NAND2_X1 U439 ( .A1(n524), .A2(n407), .ZN(n539) );
  XOR2_X1 U440 ( .A(G176GAT), .B(KEYINPUT20), .Z(n368) );
  NAND2_X1 U441 ( .A1(G227GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U442 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U443 ( .A(n369), .B(KEYINPUT82), .Z(n373) );
  XOR2_X1 U444 ( .A(KEYINPUT64), .B(G99GAT), .Z(n371) );
  XNOR2_X1 U445 ( .A(G43GAT), .B(G190GAT), .ZN(n370) );
  XNOR2_X1 U446 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U447 ( .A(n377), .B(n376), .Z(n380) );
  XOR2_X1 U448 ( .A(G120GAT), .B(G71GAT), .Z(n418) );
  XNOR2_X1 U449 ( .A(n378), .B(n418), .ZN(n379) );
  INV_X1 U450 ( .A(n530), .ZN(n543) );
  XOR2_X1 U451 ( .A(KEYINPUT88), .B(KEYINPUT22), .Z(n382) );
  XNOR2_X1 U452 ( .A(KEYINPUT85), .B(KEYINPUT87), .ZN(n381) );
  XNOR2_X1 U453 ( .A(n382), .B(n381), .ZN(n401) );
  XOR2_X1 U454 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n384) );
  XNOR2_X1 U455 ( .A(KEYINPUT84), .B(KEYINPUT86), .ZN(n383) );
  XNOR2_X1 U456 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U457 ( .A(n385), .B(G106GAT), .Z(n388) );
  XNOR2_X1 U458 ( .A(n386), .B(G218GAT), .ZN(n387) );
  XNOR2_X1 U459 ( .A(n388), .B(n387), .ZN(n394) );
  XOR2_X1 U460 ( .A(n390), .B(n389), .Z(n392) );
  NAND2_X1 U461 ( .A1(G228GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U462 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U463 ( .A(n394), .B(n393), .Z(n399) );
  XOR2_X1 U464 ( .A(G78GAT), .B(G148GAT), .Z(n396) );
  XNOR2_X1 U465 ( .A(KEYINPUT73), .B(G204GAT), .ZN(n395) );
  XNOR2_X1 U466 ( .A(n396), .B(n395), .ZN(n429) );
  XNOR2_X1 U467 ( .A(n429), .B(n397), .ZN(n398) );
  XNOR2_X1 U468 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U469 ( .A(n401), .B(n400), .ZN(n483) );
  XOR2_X1 U470 ( .A(KEYINPUT28), .B(n483), .Z(n532) );
  INV_X1 U471 ( .A(n532), .ZN(n541) );
  NAND2_X1 U472 ( .A1(n543), .A2(n541), .ZN(n402) );
  NOR2_X1 U473 ( .A1(n539), .A2(n402), .ZN(n412) );
  INV_X1 U474 ( .A(n526), .ZN(n479) );
  NOR2_X1 U475 ( .A1(n543), .A2(n479), .ZN(n403) );
  XOR2_X1 U476 ( .A(KEYINPUT96), .B(n403), .Z(n404) );
  NAND2_X1 U477 ( .A1(n404), .A2(n483), .ZN(n405) );
  XNOR2_X1 U478 ( .A(n405), .B(KEYINPUT25), .ZN(n409) );
  NOR2_X1 U479 ( .A1(n530), .A2(n483), .ZN(n406) );
  XNOR2_X1 U480 ( .A(KEYINPUT26), .B(n406), .ZN(n577) );
  AND2_X1 U481 ( .A1(n407), .A2(n577), .ZN(n408) );
  NOR2_X1 U482 ( .A1(n409), .A2(n408), .ZN(n410) );
  NOR2_X1 U483 ( .A1(n524), .A2(n410), .ZN(n411) );
  NOR2_X1 U484 ( .A1(n549), .A2(n496), .ZN(n413) );
  XNOR2_X1 U485 ( .A(KEYINPUT99), .B(n413), .ZN(n414) );
  NOR2_X1 U486 ( .A1(n592), .A2(n414), .ZN(n416) );
  XNOR2_X1 U487 ( .A(KEYINPUT37), .B(KEYINPUT100), .ZN(n415) );
  XNOR2_X1 U488 ( .A(n416), .B(n415), .ZN(n523) );
  XOR2_X1 U489 ( .A(KEYINPUT31), .B(KEYINPUT72), .Z(n420) );
  XNOR2_X1 U490 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U491 ( .A(n420), .B(n419), .ZN(n425) );
  XOR2_X1 U492 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n422) );
  XNOR2_X1 U493 ( .A(KEYINPUT32), .B(KEYINPUT33), .ZN(n421) );
  XNOR2_X1 U494 ( .A(n422), .B(n421), .ZN(n423) );
  INV_X1 U495 ( .A(KEYINPUT74), .ZN(n426) );
  XNOR2_X1 U496 ( .A(n427), .B(n426), .ZN(n434) );
  XNOR2_X1 U497 ( .A(n429), .B(n428), .ZN(n432) );
  XNOR2_X1 U498 ( .A(n430), .B(KEYINPUT71), .ZN(n431) );
  XOR2_X1 U499 ( .A(KEYINPUT66), .B(KEYINPUT68), .Z(n436) );
  XNOR2_X1 U500 ( .A(G197GAT), .B(G141GAT), .ZN(n435) );
  XNOR2_X1 U501 ( .A(n436), .B(n435), .ZN(n451) );
  XOR2_X1 U502 ( .A(G22GAT), .B(G15GAT), .Z(n438) );
  XNOR2_X1 U503 ( .A(G36GAT), .B(G50GAT), .ZN(n437) );
  XNOR2_X1 U504 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U505 ( .A(n439), .B(G113GAT), .Z(n442) );
  XNOR2_X1 U506 ( .A(G169GAT), .B(n440), .ZN(n441) );
  XNOR2_X1 U507 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U508 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n444) );
  NAND2_X1 U509 ( .A1(G229GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U510 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U511 ( .A(n446), .B(n445), .Z(n449) );
  XNOR2_X1 U512 ( .A(n447), .B(KEYINPUT29), .ZN(n448) );
  XNOR2_X1 U513 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U514 ( .A(n451), .B(n450), .ZN(n579) );
  INV_X1 U515 ( .A(n579), .ZN(n544) );
  NAND2_X1 U516 ( .A1(n470), .A2(n544), .ZN(n452) );
  XOR2_X1 U517 ( .A(KEYINPUT77), .B(n452), .Z(n499) );
  NOR2_X1 U518 ( .A1(n523), .A2(n499), .ZN(n455) );
  NAND2_X1 U519 ( .A1(n524), .A2(n510), .ZN(n459) );
  XOR2_X1 U520 ( .A(G29GAT), .B(KEYINPUT98), .Z(n457) );
  XNOR2_X1 U521 ( .A(KEYINPUT102), .B(KEYINPUT39), .ZN(n456) );
  XNOR2_X1 U522 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U523 ( .A(n459), .B(n458), .ZN(G1328GAT) );
  NAND2_X1 U524 ( .A1(n510), .A2(n530), .ZN(n463) );
  XOR2_X1 U525 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n461) );
  XNOR2_X1 U526 ( .A(n464), .B(n566), .ZN(n553) );
  INV_X1 U527 ( .A(n553), .ZN(n490) );
  INV_X1 U528 ( .A(KEYINPUT111), .ZN(n469) );
  INV_X1 U529 ( .A(n549), .ZN(n586) );
  NOR2_X1 U530 ( .A1(n586), .A2(n592), .ZN(n465) );
  XNOR2_X1 U531 ( .A(n465), .B(KEYINPUT45), .ZN(n466) );
  NAND2_X1 U532 ( .A1(n466), .A2(n470), .ZN(n467) );
  XNOR2_X1 U533 ( .A(n469), .B(n468), .ZN(n477) );
  XOR2_X1 U534 ( .A(KEYINPUT41), .B(n470), .Z(n570) );
  INV_X1 U535 ( .A(n570), .ZN(n512) );
  NAND2_X1 U536 ( .A1(n512), .A2(n544), .ZN(n472) );
  XNOR2_X1 U537 ( .A(KEYINPUT110), .B(KEYINPUT46), .ZN(n471) );
  XNOR2_X1 U538 ( .A(n472), .B(n471), .ZN(n474) );
  AND2_X1 U539 ( .A1(n566), .A2(n586), .ZN(n473) );
  AND2_X1 U540 ( .A1(n474), .A2(n473), .ZN(n475) );
  XOR2_X1 U541 ( .A(n475), .B(KEYINPUT47), .Z(n476) );
  NOR2_X1 U542 ( .A1(n477), .A2(n476), .ZN(n478) );
  XNOR2_X1 U543 ( .A(n478), .B(KEYINPUT48), .ZN(n538) );
  NOR2_X1 U544 ( .A1(n538), .A2(n479), .ZN(n481) );
  XNOR2_X1 U545 ( .A(n481), .B(n480), .ZN(n482) );
  NOR2_X1 U546 ( .A1(n524), .A2(n482), .ZN(n578) );
  NAND2_X1 U547 ( .A1(n578), .A2(n483), .ZN(n486) );
  XOR2_X1 U548 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n484) );
  XNOR2_X1 U549 ( .A(n486), .B(n485), .ZN(n487) );
  INV_X1 U550 ( .A(n487), .ZN(n488) );
  NOR2_X1 U551 ( .A1(n490), .A2(n574), .ZN(n494) );
  XNOR2_X1 U552 ( .A(KEYINPUT122), .B(KEYINPUT58), .ZN(n492) );
  INV_X1 U553 ( .A(G190GAT), .ZN(n491) );
  XNOR2_X1 U554 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n502) );
  NOR2_X1 U555 ( .A1(n586), .A2(n553), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n495), .B(KEYINPUT16), .ZN(n498) );
  INV_X1 U557 ( .A(n496), .ZN(n497) );
  NAND2_X1 U558 ( .A1(n498), .A2(n497), .ZN(n513) );
  NOR2_X1 U559 ( .A1(n499), .A2(n513), .ZN(n500) );
  XOR2_X1 U560 ( .A(KEYINPUT97), .B(n500), .Z(n506) );
  NAND2_X1 U561 ( .A1(n524), .A2(n506), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n502), .B(n501), .ZN(G1324GAT) );
  NAND2_X1 U563 ( .A1(n506), .A2(n526), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n503), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U565 ( .A(G15GAT), .B(KEYINPUT35), .Z(n505) );
  NAND2_X1 U566 ( .A1(n506), .A2(n530), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n505), .B(n504), .ZN(G1326GAT) );
  NAND2_X1 U568 ( .A1(n532), .A2(n506), .ZN(n507) );
  XNOR2_X1 U569 ( .A(n507), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U570 ( .A(G36GAT), .B(KEYINPUT103), .Z(n509) );
  NAND2_X1 U571 ( .A1(n526), .A2(n510), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(G1329GAT) );
  NAND2_X1 U573 ( .A1(n532), .A2(n510), .ZN(n511) );
  XNOR2_X1 U574 ( .A(G50GAT), .B(n511), .ZN(G1331GAT) );
  XNOR2_X1 U575 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n515) );
  NAND2_X1 U576 ( .A1(n579), .A2(n512), .ZN(n522) );
  NOR2_X1 U577 ( .A1(n522), .A2(n513), .ZN(n518) );
  NAND2_X1 U578 ( .A1(n524), .A2(n518), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n515), .B(n514), .ZN(G1332GAT) );
  NAND2_X1 U580 ( .A1(n518), .A2(n526), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n516), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U582 ( .A1(n530), .A2(n518), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n517), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT105), .B(KEYINPUT43), .Z(n520) );
  NAND2_X1 U585 ( .A1(n518), .A2(n532), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U587 ( .A(G78GAT), .B(n521), .Z(G1335GAT) );
  NOR2_X1 U588 ( .A1(n523), .A2(n522), .ZN(n533) );
  NAND2_X1 U589 ( .A1(n524), .A2(n533), .ZN(n525) );
  XNOR2_X1 U590 ( .A(G85GAT), .B(n525), .ZN(G1336GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n528) );
  NAND2_X1 U592 ( .A1(n533), .A2(n526), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U594 ( .A(G92GAT), .B(n529), .ZN(G1337GAT) );
  NAND2_X1 U595 ( .A1(n530), .A2(n533), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n531), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n537) );
  XOR2_X1 U598 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n535) );
  NAND2_X1 U599 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n537), .B(n536), .ZN(G1339GAT) );
  NOR2_X1 U602 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U603 ( .A(n540), .B(KEYINPUT112), .ZN(n558) );
  NAND2_X1 U604 ( .A1(n541), .A2(n558), .ZN(n542) );
  NOR2_X1 U605 ( .A1(n543), .A2(n542), .ZN(n554) );
  NAND2_X1 U606 ( .A1(n544), .A2(n554), .ZN(n545) );
  XNOR2_X1 U607 ( .A(G113GAT), .B(n545), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n547) );
  NAND2_X1 U609 ( .A1(n554), .A2(n512), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U611 ( .A(G120GAT), .B(n548), .Z(G1341GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n551) );
  NAND2_X1 U613 ( .A1(n554), .A2(n549), .ZN(n550) );
  XNOR2_X1 U614 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U615 ( .A(G127GAT), .B(n552), .Z(G1342GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n556) );
  NAND2_X1 U617 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U618 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U619 ( .A(G134GAT), .B(n557), .Z(G1343GAT) );
  NAND2_X1 U620 ( .A1(n577), .A2(n558), .ZN(n565) );
  NOR2_X1 U621 ( .A1(n579), .A2(n565), .ZN(n559) );
  XOR2_X1 U622 ( .A(G141GAT), .B(n559), .Z(G1344GAT) );
  NOR2_X1 U623 ( .A1(n570), .A2(n565), .ZN(n561) );
  XNOR2_X1 U624 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(n562), .ZN(G1345GAT) );
  NOR2_X1 U627 ( .A1(n586), .A2(n565), .ZN(n563) );
  XOR2_X1 U628 ( .A(KEYINPUT116), .B(n563), .Z(n564) );
  XNOR2_X1 U629 ( .A(G155GAT), .B(n564), .ZN(G1346GAT) );
  NOR2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n568) );
  XNOR2_X1 U631 ( .A(G162GAT), .B(KEYINPUT117), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n568), .B(n567), .ZN(G1347GAT) );
  NOR2_X1 U633 ( .A1(n574), .A2(n579), .ZN(n569) );
  XOR2_X1 U634 ( .A(G169GAT), .B(n569), .Z(G1348GAT) );
  XNOR2_X1 U635 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n572) );
  NOR2_X1 U636 ( .A1(n570), .A2(n574), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(G176GAT), .ZN(G1349GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n586), .ZN(n576) );
  XNOR2_X1 U640 ( .A(G183GAT), .B(KEYINPUT121), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1350GAT) );
  NAND2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n591) );
  NOR2_X1 U643 ( .A1(n579), .A2(n591), .ZN(n581) );
  XNOR2_X1 U644 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(n582), .ZN(G1352GAT) );
  NOR2_X1 U647 ( .A1(n470), .A2(n591), .ZN(n584) );
  XNOR2_X1 U648 ( .A(KEYINPUT123), .B(KEYINPUT61), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n585) );
  XOR2_X1 U650 ( .A(G204GAT), .B(n585), .Z(G1353GAT) );
  NOR2_X1 U651 ( .A1(n586), .A2(n591), .ZN(n587) );
  XOR2_X1 U652 ( .A(KEYINPUT124), .B(n587), .Z(n588) );
  XNOR2_X1 U653 ( .A(G211GAT), .B(n588), .ZN(G1354GAT) );
  XOR2_X1 U654 ( .A(KEYINPUT125), .B(KEYINPUT62), .Z(n590) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n589) );
  XNOR2_X1 U656 ( .A(n590), .B(n589), .ZN(n594) );
  NOR2_X1 U657 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U658 ( .A(n594), .B(n593), .Z(G1355GAT) );
endmodule

