//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 0 0 1 1 0 0 0 1 0 1 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n631,
    new_n632, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n789, new_n790, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n872, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914;
  XNOR2_X1  g000(.A(G113gat), .B(G120gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n203));
  XOR2_X1   g002(.A(G127gat), .B(G134gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT25), .ZN(new_n207));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT24), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n209), .A2(G183gat), .A3(G190gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT24), .ZN(new_n212));
  NOR2_X1   g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n208), .B(new_n210), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G169gat), .ZN(new_n215));
  INV_X1    g014(.A(G176gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT23), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(G169gat), .B2(G176gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  OAI211_X1 g019(.A(KEYINPUT64), .B(new_n207), .C1(new_n214), .C2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n223), .A2(new_n209), .B1(G169gat), .B2(G176gat), .ZN(new_n224));
  INV_X1    g023(.A(G183gat), .ZN(new_n225));
  INV_X1    g024(.A(G190gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(KEYINPUT24), .A3(new_n211), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n224), .A2(new_n228), .A3(new_n219), .A4(new_n217), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n207), .B1(new_n229), .B2(KEYINPUT64), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n222), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT26), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT26), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(G169gat), .B2(G176gat), .ZN(new_n234));
  INV_X1    g033(.A(new_n208), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n211), .B(new_n232), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT27), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT27), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(KEYINPUT65), .A3(G183gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n240), .A3(new_n226), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n238), .A2(new_n240), .A3(KEYINPUT66), .A4(new_n226), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT27), .B(G183gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n247), .A2(KEYINPUT28), .A3(new_n226), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n236), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n206), .B1(new_n231), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n246), .A2(new_n248), .ZN(new_n251));
  INV_X1    g050(.A(new_n236), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT64), .B1(new_n214), .B2(new_n220), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT25), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(new_n221), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n253), .A2(new_n205), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n250), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G227gat), .ZN(new_n259));
  INV_X1    g058(.A(G233gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT68), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n263));
  INV_X1    g062(.A(new_n261), .ZN(new_n264));
  AOI211_X1 g063(.A(new_n263), .B(new_n264), .C1(new_n250), .C2(new_n257), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT32), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT33), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n267), .B1(new_n262), .B2(new_n265), .ZN(new_n268));
  XOR2_X1   g067(.A(G15gat), .B(G43gat), .Z(new_n269));
  XNOR2_X1  g068(.A(G71gat), .B(G99gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n266), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT69), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n271), .A2(KEYINPUT33), .ZN(new_n274));
  OR2_X1    g073(.A1(new_n266), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n266), .A2(new_n268), .A3(new_n276), .A4(new_n271), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n273), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n250), .A2(new_n264), .A3(new_n257), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT34), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n280), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n273), .A2(new_n282), .A3(new_n275), .A4(new_n277), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n281), .A2(KEYINPUT36), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT70), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n281), .A2(new_n286), .A3(KEYINPUT36), .A4(new_n283), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT72), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n281), .A2(new_n289), .A3(new_n283), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n278), .A2(KEYINPUT72), .A3(new_n280), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT71), .B(KEYINPUT36), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n294));
  OR2_X1    g093(.A1(new_n294), .A2(KEYINPUT73), .ZN(new_n295));
  XNOR2_X1  g094(.A(G197gat), .B(G204gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(KEYINPUT73), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(G211gat), .B(G218gat), .Z(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G141gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G148gat), .ZN(new_n302));
  XOR2_X1   g101(.A(KEYINPUT76), .B(G148gat), .Z(new_n303));
  OAI21_X1  g102(.A(new_n302), .B1(new_n303), .B2(new_n301), .ZN(new_n304));
  NAND2_X1  g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305));
  INV_X1    g104(.A(G155gat), .ZN(new_n306));
  INV_X1    g105(.A(G162gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n305), .B1(new_n308), .B2(KEYINPUT2), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  XOR2_X1   g109(.A(KEYINPUT75), .B(KEYINPUT2), .Z(new_n311));
  XNOR2_X1  g110(.A(G141gat), .B(G148gat), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n305), .B(new_n308), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT3), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT29), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n300), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n319), .B1(G228gat), .B2(G233gat), .ZN(new_n320));
  INV_X1    g119(.A(new_n300), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT82), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n298), .A2(new_n299), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT82), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT29), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT3), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n320), .B1(new_n315), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n300), .A2(new_n318), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n315), .B1(new_n328), .B2(new_n316), .ZN(new_n329));
  OAI211_X1 g128(.A(G228gat), .B(G233gat), .C1(new_n319), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G78gat), .B(G106gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(G22gat), .ZN(new_n333));
  XOR2_X1   g132(.A(KEYINPUT31), .B(G50gat), .Z(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n331), .B(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(G57gat), .B(G85gat), .Z(new_n337));
  XNOR2_X1  g136(.A(G1gat), .B(G29gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n337), .B(new_n338), .ZN(new_n339));
  XOR2_X1   g138(.A(KEYINPUT79), .B(KEYINPUT0), .Z(new_n340));
  XNOR2_X1  g139(.A(new_n340), .B(KEYINPUT80), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n339), .B(new_n341), .Z(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(KEYINPUT83), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT84), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n344), .A2(KEYINPUT40), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G225gat), .A2(G233gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n347), .B(KEYINPUT77), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n315), .A2(new_n205), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n206), .A2(new_n314), .ZN(new_n351));
  OAI211_X1 g150(.A(KEYINPUT39), .B(new_n349), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n314), .A2(KEYINPUT3), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n317), .A2(new_n206), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT4), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n355), .B1(new_n206), .B2(new_n314), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n351), .A2(KEYINPUT4), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n354), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(KEYINPUT39), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n346), .B(new_n352), .C1(new_n359), .C2(new_n349), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n344), .A2(KEYINPUT40), .ZN(new_n361));
  OR2_X1    g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n354), .A2(new_n357), .A3(new_n349), .A4(new_n356), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT78), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n348), .B1(new_n350), .B2(new_n351), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT5), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n364), .A2(new_n367), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n343), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n360), .A2(new_n361), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n362), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  AOI22_X1  g174(.A1(new_n251), .A2(new_n252), .B1(new_n255), .B2(new_n221), .ZN(new_n376));
  INV_X1    g175(.A(G226gat), .ZN(new_n377));
  OAI22_X1  g176(.A1(new_n376), .A2(KEYINPUT29), .B1(new_n377), .B2(new_n260), .ZN(new_n378));
  OAI211_X1 g177(.A(G226gat), .B(G233gat), .C1(new_n231), .C2(new_n249), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(new_n300), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n300), .B1(new_n378), .B2(new_n379), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G8gat), .B(G36gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(G64gat), .B(G92gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT30), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT74), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n391), .B1(new_n381), .B2(new_n382), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n378), .A2(new_n379), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(new_n321), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n394), .A2(KEYINPUT74), .A3(new_n380), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n392), .A2(new_n386), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n383), .A2(KEYINPUT30), .A3(new_n387), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n390), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n336), .B1(new_n375), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n392), .A2(KEYINPUT37), .A3(new_n395), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n386), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT87), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT86), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT37), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n404), .B1(new_n383), .B2(new_n405), .ZN(new_n406));
  NOR4_X1   g205(.A1(new_n381), .A2(new_n382), .A3(KEYINPUT86), .A4(KEYINPUT37), .ZN(new_n407));
  OR2_X1    g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  XOR2_X1   g207(.A(KEYINPUT85), .B(KEYINPUT38), .Z(new_n409));
  NAND3_X1  g208(.A1(new_n400), .A2(KEYINPUT87), .A3(new_n386), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n403), .A2(new_n408), .A3(new_n409), .A4(new_n410), .ZN(new_n411));
  OAI221_X1 g210(.A(new_n386), .B1(new_n405), .B2(new_n383), .C1(new_n406), .C2(new_n407), .ZN(new_n412));
  INV_X1    g211(.A(new_n409), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n342), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT6), .B1(new_n371), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n369), .A2(new_n370), .A3(new_n342), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n373), .A2(new_n417), .B1(KEYINPUT6), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n415), .A2(new_n388), .A3(new_n420), .ZN(new_n421));
  AOI22_X1  g220(.A1(new_n288), .A2(new_n293), .B1(new_n399), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n417), .A2(KEYINPUT81), .A3(new_n418), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT81), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n372), .B(new_n342), .C1(new_n424), .C2(KEYINPUT6), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n398), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n336), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n281), .A2(new_n283), .ZN(new_n430));
  INV_X1    g229(.A(new_n336), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT35), .B1(new_n432), .B2(new_n428), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n290), .A2(new_n291), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n420), .A2(KEYINPUT35), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n434), .A2(new_n427), .A3(new_n435), .A4(new_n431), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n422), .A2(new_n429), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT95), .ZN(new_n440));
  INV_X1    g239(.A(G57gat), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n441), .A2(G64gat), .ZN(new_n442));
  INV_X1    g241(.A(G64gat), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n443), .A2(G57gat), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n440), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n443), .A2(G57gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n441), .A2(G64gat), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(new_n447), .A3(KEYINPUT95), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n445), .A2(KEYINPUT9), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(G71gat), .A2(G78gat), .ZN(new_n450));
  OR2_X1    g249(.A1(G71gat), .A2(G78gat), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT96), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n449), .A2(KEYINPUT96), .A3(new_n450), .A4(new_n451), .ZN(new_n455));
  AND2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT9), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n450), .B1(new_n451), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n458), .B1(new_n442), .B2(new_n444), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n456), .A2(KEYINPUT21), .A3(new_n459), .ZN(new_n460));
  NOR2_X1   g259(.A1(G15gat), .A2(G22gat), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT91), .ZN(new_n463));
  NAND2_X1  g262(.A1(G15gat), .A2(G22gat), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  AND2_X1   g264(.A1(G15gat), .A2(G22gat), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT91), .B1(new_n466), .B2(new_n461), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(G1gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT16), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n470), .B(KEYINPUT92), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n465), .A2(new_n467), .A3(new_n469), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(G8gat), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n475), .B1(new_n473), .B2(KEYINPUT93), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n472), .B(new_n473), .C1(KEYINPUT93), .C2(new_n475), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n460), .A2(new_n225), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n225), .B1(new_n460), .B2(new_n479), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n439), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n482), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n484), .A2(new_n480), .A3(new_n438), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n454), .A2(new_n459), .A3(new_n455), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT21), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  XOR2_X1   g288(.A(new_n489), .B(KEYINPUT97), .Z(new_n490));
  NAND2_X1  g289(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n490), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n483), .A2(new_n485), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G127gat), .B(G155gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(G211gat), .ZN(new_n496));
  AND2_X1   g295(.A1(G231gat), .A2(G233gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n491), .A2(new_n498), .A3(new_n493), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT7), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT98), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT98), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT7), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n504), .A2(new_n506), .A3(G85gat), .A4(G92gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(G99gat), .A2(G106gat), .ZN(new_n508));
  INV_X1    g307(.A(G85gat), .ZN(new_n509));
  INV_X1    g308(.A(G92gat), .ZN(new_n510));
  AOI22_X1  g309(.A1(KEYINPUT8), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI211_X1 g310(.A(KEYINPUT98), .B(new_n503), .C1(new_n509), .C2(new_n510), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n507), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(G99gat), .B(G106gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT88), .ZN(new_n517));
  INV_X1    g316(.A(G43gat), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n517), .B1(new_n518), .B2(G50gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(G50gat), .ZN(new_n520));
  INV_X1    g319(.A(G50gat), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n521), .A2(KEYINPUT88), .A3(G43gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT15), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT89), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT15), .B1(new_n518), .B2(G50gat), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n527), .B1(new_n518), .B2(G50gat), .ZN(new_n528));
  AND2_X1   g327(.A1(G29gat), .A2(G36gat), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR3_X1   g329(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n531), .A2(KEYINPUT90), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(KEYINPUT90), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT89), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n523), .A2(new_n536), .A3(new_n524), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n526), .A2(new_n530), .A3(new_n535), .A4(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT17), .ZN(new_n539));
  INV_X1    g338(.A(new_n534), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n540), .A2(new_n531), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n528), .B1(new_n541), .B2(new_n529), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n538), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n539), .B1(new_n538), .B2(new_n542), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n516), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n538), .A2(new_n542), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(new_n515), .ZN(new_n547));
  NAND3_X1  g346(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n545), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT41), .ZN(new_n550));
  NAND2_X1  g349(.A1(G232gat), .A2(G233gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n550), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n545), .A2(new_n553), .A3(new_n547), .A4(new_n548), .ZN(new_n554));
  XNOR2_X1  g353(.A(G134gat), .B(G162gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT99), .ZN(new_n556));
  XOR2_X1   g355(.A(G190gat), .B(G218gat), .Z(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n552), .A2(new_n554), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n558), .B1(new_n552), .B2(new_n554), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n502), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G230gat), .A2(G233gat), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n487), .A2(new_n516), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT10), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n515), .A2(new_n454), .A3(new_n459), .A4(new_n455), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n456), .A2(KEYINPUT10), .A3(new_n459), .A4(new_n515), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n565), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n564), .B1(new_n566), .B2(new_n568), .ZN(new_n572));
  OR2_X1    g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G176gat), .B(G204gat), .ZN(new_n574));
  INV_X1    g373(.A(G148gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(KEYINPUT100), .B(G120gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n573), .B(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n479), .B1(new_n543), .B2(new_n544), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n477), .A2(new_n478), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(new_n546), .ZN(new_n584));
  NAND2_X1  g383(.A1(G229gat), .A2(G233gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n582), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT18), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n585), .B(KEYINPUT13), .Z(new_n589));
  INV_X1    g388(.A(new_n584), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n583), .A2(new_n546), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n582), .A2(KEYINPUT18), .A3(new_n584), .A4(new_n585), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n588), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G113gat), .B(G141gat), .ZN(new_n595));
  INV_X1    g394(.A(G197gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT11), .B(G169gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT12), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n594), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT94), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n588), .A2(new_n600), .A3(new_n592), .A4(new_n593), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n594), .A2(KEYINPUT94), .A3(new_n601), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n581), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NOR3_X1   g408(.A1(new_n437), .A2(new_n563), .A3(new_n609), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n423), .A2(new_n425), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(KEYINPUT101), .B(G1gat), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(G1324gat));
  AND2_X1   g413(.A1(new_n610), .A2(new_n398), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT16), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n616), .A2(new_n475), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n475), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n615), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT42), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n622), .B(new_n623), .C1(new_n475), .C2(new_n615), .ZN(G1325gat));
  AOI21_X1  g423(.A(G15gat), .B1(new_n610), .B2(new_n434), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n290), .A2(new_n291), .ZN(new_n626));
  AOI22_X1  g425(.A1(new_n626), .A2(new_n292), .B1(new_n285), .B2(new_n287), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT102), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n628), .A2(G15gat), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n625), .B1(new_n610), .B2(new_n629), .ZN(G1326gat));
  NAND2_X1  g429(.A1(new_n610), .A2(new_n336), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT43), .B(G22gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(G1327gat));
  NAND2_X1  g432(.A1(new_n288), .A2(new_n293), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n421), .A2(new_n399), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n634), .A2(new_n429), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n433), .A2(new_n436), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n561), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n609), .A2(new_n502), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OR3_X1    g441(.A1(new_n642), .A2(G29gat), .A3(new_n426), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT45), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT44), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n645), .B1(new_n437), .B2(new_n562), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n638), .A2(KEYINPUT44), .A3(new_n561), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n641), .B(KEYINPUT103), .Z(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(G29gat), .B1(new_n650), .B2(new_n426), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n644), .A2(new_n651), .ZN(G1328gat));
  NOR3_X1   g451(.A1(new_n642), .A2(G36gat), .A3(new_n427), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT46), .ZN(new_n654));
  OAI21_X1  g453(.A(KEYINPUT104), .B1(new_n650), .B2(new_n427), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n648), .A2(new_n656), .A3(new_n398), .A4(new_n649), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n655), .A2(G36gat), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n654), .A2(new_n658), .ZN(G1329gat));
  OAI21_X1  g458(.A(G43gat), .B1(new_n650), .B2(new_n634), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n642), .A2(G43gat), .A3(new_n626), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n660), .A2(KEYINPUT47), .A3(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n648), .A2(new_n628), .A3(new_n649), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n661), .B1(new_n664), .B2(G43gat), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n663), .B1(KEYINPUT47), .B2(new_n665), .ZN(G1330gat));
  INV_X1    g465(.A(KEYINPUT48), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n640), .A2(new_n521), .A3(new_n336), .A4(new_n641), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n667), .B1(new_n668), .B2(KEYINPUT106), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n646), .A2(new_n647), .A3(new_n336), .A4(new_n649), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(G50gat), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n669), .B(new_n671), .C1(KEYINPUT106), .C2(new_n668), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(KEYINPUT105), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n670), .A2(new_n674), .A3(G50gat), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n673), .A2(new_n668), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n672), .B1(new_n676), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g476(.A(new_n607), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n563), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n638), .A2(new_n581), .A3(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n680), .A2(new_n426), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(new_n441), .ZN(G1332gat));
  XNOR2_X1  g481(.A(new_n680), .B(KEYINPUT107), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT108), .ZN(new_n684));
  NAND2_X1  g483(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n683), .A2(new_n684), .A3(new_n398), .A4(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n680), .A2(KEYINPUT107), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT107), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n580), .B1(new_n636), .B2(new_n637), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n688), .B1(new_n689), .B2(new_n679), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n398), .B(new_n685), .C1(new_n687), .C2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT108), .ZN(new_n692));
  NOR2_X1   g491(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n693));
  AND3_X1   g492(.A1(new_n686), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n693), .B1(new_n686), .B2(new_n692), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(G1333gat));
  NOR2_X1   g495(.A1(new_n687), .A2(new_n690), .ZN(new_n697));
  INV_X1    g496(.A(new_n628), .ZN(new_n698));
  OAI21_X1  g497(.A(G71gat), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT50), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT109), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(new_n680), .B2(new_n626), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n689), .A2(KEYINPUT109), .A3(new_n434), .A4(new_n679), .ZN(new_n703));
  AOI21_X1  g502(.A(G71gat), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n699), .A2(new_n700), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n700), .B1(new_n699), .B2(new_n705), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(G1334gat));
  NAND2_X1  g507(.A1(new_n683), .A2(new_n336), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g509(.A1(new_n611), .A2(new_n509), .A3(new_n581), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT111), .ZN(new_n712));
  NAND2_X1  g511(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n502), .A2(new_n678), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n714), .B1(new_n640), .B2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n715), .ZN(new_n717));
  NOR2_X1   g516(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n639), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n712), .B1(new_n716), .B2(new_n720), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n646), .A2(new_n647), .A3(new_n581), .A4(new_n715), .ZN(new_n722));
  OAI21_X1  g521(.A(G85gat), .B1(new_n722), .B2(new_n426), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT112), .ZN(G1336gat));
  OAI21_X1  g524(.A(G92gat), .B1(new_n722), .B2(new_n427), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT52), .B1(new_n726), .B2(KEYINPUT114), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n581), .A2(new_n510), .A3(new_n398), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT113), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n729), .B1(new_n716), .B2(new_n720), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n726), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n730), .B(new_n726), .C1(KEYINPUT114), .C2(KEYINPUT52), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(G1337gat));
  NOR2_X1   g533(.A1(new_n626), .A2(G99gat), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n581), .B(new_n735), .C1(new_n716), .C2(new_n720), .ZN(new_n736));
  OAI21_X1  g535(.A(G99gat), .B1(new_n722), .B2(new_n698), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(G1338gat));
  NOR2_X1   g537(.A1(new_n431), .A2(G106gat), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n581), .B(new_n739), .C1(new_n716), .C2(new_n720), .ZN(new_n740));
  OAI21_X1  g539(.A(G106gat), .B1(new_n722), .B2(new_n431), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g542(.A1(new_n569), .A2(new_n570), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT54), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n744), .A2(new_n745), .A3(new_n564), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n569), .A2(new_n570), .A3(new_n565), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT54), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n578), .B(new_n746), .C1(new_n748), .C2(new_n571), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT116), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT55), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n750), .B1(new_n749), .B2(new_n751), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT115), .B1(new_n749), .B2(new_n751), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n573), .A2(new_n578), .ZN(new_n756));
  INV_X1    g555(.A(new_n571), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n757), .A2(KEYINPUT54), .A3(new_n747), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n579), .B1(new_n571), .B2(new_n745), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n758), .A2(new_n759), .A3(new_n760), .A4(KEYINPUT55), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n755), .A2(new_n756), .A3(new_n761), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n754), .A2(new_n762), .A3(new_n607), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n590), .A2(new_n591), .A3(new_n589), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n585), .B1(new_n582), .B2(new_n584), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n599), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n604), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n580), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n562), .B1(new_n763), .B2(new_n768), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n755), .A2(new_n756), .A3(new_n761), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n749), .A2(new_n751), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT116), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n767), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n770), .A2(new_n561), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n502), .B1(new_n769), .B2(new_n776), .ZN(new_n777));
  AND4_X1   g576(.A1(new_n502), .A2(new_n562), .A3(new_n580), .A4(new_n607), .ZN(new_n778));
  OR2_X1    g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n779), .A2(new_n611), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n626), .A2(new_n336), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n780), .A2(new_n427), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(KEYINPUT117), .ZN(new_n783));
  OAI21_X1  g582(.A(G113gat), .B1(new_n783), .B2(new_n607), .ZN(new_n784));
  INV_X1    g583(.A(new_n432), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n780), .A2(new_n427), .A3(new_n785), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n786), .A2(G113gat), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n784), .B1(new_n607), .B2(new_n787), .ZN(G1340gat));
  OAI21_X1  g587(.A(G120gat), .B1(new_n783), .B2(new_n580), .ZN(new_n789));
  OR2_X1    g588(.A1(new_n580), .A2(G120gat), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n789), .B1(new_n786), .B2(new_n790), .ZN(G1341gat));
  INV_X1    g590(.A(G127gat), .ZN(new_n792));
  INV_X1    g591(.A(new_n502), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n783), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n786), .A2(new_n793), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n795), .A2(G127gat), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n794), .A2(new_n796), .ZN(G1342gat));
  NOR3_X1   g596(.A1(new_n786), .A2(G134gat), .A3(new_n562), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(KEYINPUT56), .ZN(new_n799));
  OAI21_X1  g598(.A(G134gat), .B1(new_n783), .B2(new_n562), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(G1343gat));
  INV_X1    g600(.A(KEYINPUT58), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n803), .B(new_n336), .C1(new_n777), .C2(new_n778), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n605), .A2(new_n606), .A3(new_n771), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n768), .B1(new_n770), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n776), .B1(new_n806), .B2(new_n561), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n778), .B1(new_n807), .B2(new_n793), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT57), .B1(new_n808), .B2(new_n431), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n611), .A2(new_n427), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT118), .B1(new_n627), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n812));
  INV_X1    g611(.A(new_n810), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n634), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n804), .A2(new_n809), .A3(new_n811), .A4(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(G141gat), .B1(new_n815), .B2(new_n607), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n628), .A2(new_n431), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n780), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT121), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT121), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n817), .A2(new_n820), .A3(new_n780), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n819), .A2(new_n427), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n607), .A2(G141gat), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n802), .B(new_n816), .C1(new_n822), .C2(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n817), .A2(new_n427), .A3(new_n780), .A4(new_n823), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n815), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n812), .B1(new_n634), .B2(new_n813), .ZN(new_n829));
  AOI211_X1 g628(.A(KEYINPUT118), .B(new_n810), .C1(new_n288), .C2(new_n293), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n831), .A2(KEYINPUT119), .A3(new_n809), .A4(new_n804), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n607), .B1(new_n828), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n826), .B1(new_n833), .B2(new_n301), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n834), .A2(KEYINPUT120), .A3(KEYINPUT58), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT120), .B1(new_n834), .B2(KEYINPUT58), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n825), .B1(new_n835), .B2(new_n836), .ZN(G1344gat));
  INV_X1    g636(.A(KEYINPUT59), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n580), .B1(new_n828), .B2(new_n832), .ZN(new_n839));
  INV_X1    g638(.A(new_n303), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n779), .A2(new_n336), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT57), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n754), .A2(new_n762), .A3(new_n562), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n844), .A2(KEYINPUT122), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(KEYINPUT122), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n845), .A2(new_n775), .A3(new_n846), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n806), .A2(new_n561), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n502), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n803), .B(new_n336), .C1(new_n849), .C2(new_n778), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n843), .A2(new_n581), .A3(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n831), .ZN(new_n852));
  OAI21_X1  g651(.A(KEYINPUT59), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n581), .A2(new_n840), .ZN(new_n854));
  OAI221_X1 g653(.A(new_n841), .B1(new_n853), .B2(new_n575), .C1(new_n822), .C2(new_n854), .ZN(G1345gat));
  AOI211_X1 g654(.A(new_n306), .B(new_n793), .C1(new_n828), .C2(new_n832), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n822), .A2(new_n793), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n856), .B1(new_n857), .B2(new_n306), .ZN(G1346gat));
  OR2_X1    g657(.A1(new_n822), .A2(G162gat), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n562), .B1(new_n828), .B2(new_n832), .ZN(new_n860));
  OAI22_X1  g659(.A1(new_n859), .A2(new_n562), .B1(new_n307), .B2(new_n860), .ZN(G1347gat));
  AND2_X1   g660(.A1(new_n779), .A2(new_n426), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n862), .A2(new_n398), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n863), .A2(G169gat), .A3(new_n781), .A4(new_n678), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT123), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n865), .B1(new_n432), .B2(new_n427), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n785), .A2(KEYINPUT123), .A3(new_n398), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n862), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n215), .B1(new_n868), .B2(new_n607), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n864), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(KEYINPUT124), .ZN(G1348gat));
  OAI21_X1  g670(.A(new_n216), .B1(new_n868), .B2(new_n580), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT125), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n863), .A2(G176gat), .A3(new_n781), .A4(new_n581), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(G1349gat));
  NAND3_X1  g674(.A1(new_n863), .A2(new_n502), .A3(new_n781), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(G183gat), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n502), .A2(new_n247), .ZN(new_n878));
  OR2_X1    g677(.A1(new_n868), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g678(.A(KEYINPUT126), .B(KEYINPUT60), .ZN(new_n880));
  AND3_X1   g679(.A1(new_n877), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n880), .B1(new_n877), .B2(new_n879), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(G1350gat));
  OR3_X1    g682(.A1(new_n868), .A2(G190gat), .A3(new_n562), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n863), .A2(new_n561), .A3(new_n781), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT61), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n885), .A2(new_n886), .A3(G190gat), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n885), .B2(G190gat), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n884), .B1(new_n887), .B2(new_n888), .ZN(G1351gat));
  NAND2_X1  g688(.A1(new_n863), .A2(new_n817), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n596), .A3(new_n678), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n843), .A2(new_n850), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n698), .A2(new_n426), .A3(new_n398), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n893), .A2(new_n607), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n892), .B1(new_n596), .B2(new_n895), .ZN(G1352gat));
  OR4_X1    g695(.A1(KEYINPUT62), .A2(new_n890), .A3(G204gat), .A4(new_n580), .ZN(new_n897));
  INV_X1    g696(.A(G204gat), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n891), .A2(new_n898), .A3(new_n581), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT62), .ZN(new_n900));
  OAI21_X1  g699(.A(G204gat), .B1(new_n851), .B2(new_n894), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n897), .A2(new_n900), .A3(new_n901), .ZN(G1353gat));
  OR3_X1    g701(.A1(new_n890), .A2(G211gat), .A3(new_n793), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n893), .A2(new_n894), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n502), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n905), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT63), .B1(new_n905), .B2(G211gat), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(G1354gat));
  INV_X1    g707(.A(KEYINPUT127), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n904), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT127), .B1(new_n893), .B2(new_n894), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(new_n561), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(G218gat), .ZN(new_n913));
  OR3_X1    g712(.A1(new_n890), .A2(G218gat), .A3(new_n562), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1355gat));
endmodule


