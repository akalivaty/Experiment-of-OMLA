//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 1 0 0 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1300, new_n1301, new_n1302;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n204), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G13), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT0), .Z(new_n215));
  INV_X1    g0015(.A(KEYINPUT1), .ZN(new_n216));
  XOR2_X1   g0016(.A(KEYINPUT69), .B(G238), .Z(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT68), .B(G68), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G107), .A2(G264), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n224));
  AND4_X1   g0024(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n210), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n215), .B1(new_n216), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n227), .B1(new_n216), .B2(new_n226), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G20), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT65), .ZN(new_n232));
  INV_X1    g0032(.A(G50), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n204), .A2(new_n205), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n233), .B1(new_n234), .B2(KEYINPUT66), .ZN(new_n235));
  OAI21_X1  g0035(.A(new_n235), .B1(KEYINPUT66), .B2(new_n234), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(KEYINPUT67), .Z(new_n237));
  AOI21_X1  g0037(.A(new_n228), .B1(new_n232), .B2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  INV_X1    g0039(.A(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT2), .B(G226), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G264), .B(G270), .Z(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G50), .B(G68), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G58), .B(G77), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  AOI21_X1  g0058(.A(G1698), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G222), .ZN(new_n260));
  INV_X1    g0060(.A(G77), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n257), .A2(new_n258), .ZN(new_n262));
  INV_X1    g0062(.A(G223), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(G1698), .ZN(new_n264));
  OAI221_X1 g0064(.A(new_n260), .B1(new_n261), .B2(new_n262), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G41), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(new_n229), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(KEYINPUT70), .B1(new_n267), .B2(new_n229), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT70), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n266), .A2(new_n273), .A3(G1), .A4(G13), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n270), .A2(G274), .A3(new_n272), .A4(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n270), .A2(new_n274), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(new_n272), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n276), .B1(G226), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n269), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT71), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n269), .A2(new_n279), .A3(KEYINPUT71), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G179), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n287), .A2(new_n229), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n208), .A2(G20), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G50), .ZN(new_n292));
  OAI22_X1  g0092(.A1(new_n290), .A2(new_n292), .B1(G50), .B2(new_n289), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n209), .B1(new_n234), .B2(new_n233), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT72), .ZN(new_n296));
  XOR2_X1   g0096(.A(KEYINPUT8), .B(G58), .Z(new_n297));
  NAND2_X1  g0097(.A1(new_n209), .A2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(G20), .A2(G33), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n297), .A2(new_n299), .B1(G150), .B2(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n296), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n294), .B1(new_n302), .B2(new_n288), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n282), .A2(new_n304), .A3(new_n283), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n286), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n284), .A2(G190), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT9), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n282), .A2(G200), .A3(new_n283), .ZN(new_n310));
  OAI211_X1 g0110(.A(KEYINPUT9), .B(new_n294), .C1(new_n302), .C2(new_n288), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n307), .A2(new_n309), .A3(new_n310), .A4(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT10), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n312), .A2(KEYINPUT10), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n306), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n290), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n317), .A2(G77), .A3(new_n291), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n297), .A2(new_n300), .B1(G20), .B2(G77), .ZN(new_n319));
  XOR2_X1   g0119(.A(KEYINPUT15), .B(G87), .Z(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n299), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n288), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n289), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT73), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n323), .A2(new_n324), .A3(new_n261), .ZN(new_n325));
  OAI21_X1  g0125(.A(KEYINPUT73), .B1(new_n289), .B2(G77), .ZN(new_n326));
  AOI211_X1 g0126(.A(new_n318), .B(new_n322), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n276), .B1(G244), .B2(new_n278), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n262), .A2(G232), .ZN(new_n329));
  INV_X1    g0129(.A(G107), .ZN(new_n330));
  OAI22_X1  g0130(.A1(new_n329), .A2(G1698), .B1(new_n330), .B2(new_n262), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n264), .A2(new_n217), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n268), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n327), .B1(new_n334), .B2(new_n304), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(G179), .B2(new_n334), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(G200), .ZN(new_n337));
  INV_X1    g0137(.A(G190), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n327), .B(new_n337), .C1(new_n338), .C2(new_n334), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n297), .A2(new_n291), .ZN(new_n341));
  OAI22_X1  g0141(.A1(new_n341), .A2(new_n290), .B1(new_n289), .B2(new_n297), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT77), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n342), .B(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n203), .A2(KEYINPUT68), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT68), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G68), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n202), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(G20), .B1(new_n348), .B2(new_n234), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n300), .A2(G159), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n257), .A2(new_n209), .A3(new_n258), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT7), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n257), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n258), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n203), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n288), .B1(new_n357), .B2(KEYINPUT16), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n354), .A2(KEYINPUT76), .A3(new_n355), .ZN(new_n359));
  INV_X1    g0159(.A(new_n218), .ZN(new_n360));
  OR2_X1    g0160(.A1(new_n355), .A2(KEYINPUT76), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n204), .B(new_n205), .C1(new_n218), .C2(new_n202), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n363), .A2(G20), .B1(G159), .B2(new_n300), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT16), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n344), .B1(new_n358), .B2(new_n367), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n270), .A2(G232), .A3(new_n271), .A4(new_n274), .ZN(new_n369));
  NOR2_X1   g0169(.A1(G223), .A2(G1698), .ZN(new_n370));
  INV_X1    g0170(.A(G226), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n370), .B1(new_n371), .B2(G1698), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n372), .A2(new_n262), .B1(G33), .B2(G87), .ZN(new_n373));
  INV_X1    g0173(.A(new_n268), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n275), .B(new_n369), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G169), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n371), .A2(G1698), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(G223), .B2(G1698), .ZN(new_n378));
  AND2_X1   g0178(.A1(KEYINPUT3), .A2(G33), .ZN(new_n379));
  NOR2_X1   g0179(.A1(KEYINPUT3), .A2(G33), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G87), .ZN(new_n382));
  OAI22_X1  g0182(.A1(new_n378), .A2(new_n381), .B1(new_n256), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n268), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n384), .A2(G179), .A3(new_n275), .A4(new_n369), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n376), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT18), .B1(new_n368), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g0188(.A(new_n342), .B(KEYINPUT77), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT7), .B1(new_n381), .B2(new_n209), .ZN(new_n390));
  INV_X1    g0190(.A(new_n355), .ZN(new_n391));
  OAI21_X1  g0191(.A(G68), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n364), .A2(KEYINPUT16), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n287), .A2(new_n229), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT16), .B1(new_n362), .B2(new_n364), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n389), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT18), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(new_n386), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G200), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n375), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n384), .A2(new_n338), .A3(new_n275), .A4(new_n369), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n403), .B(new_n389), .C1(new_n395), .C2(new_n396), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT17), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n358), .A2(new_n367), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n407), .A2(KEYINPUT17), .A3(new_n389), .A4(new_n403), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n388), .A2(new_n399), .A3(new_n406), .A4(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n340), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n360), .A2(new_n209), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n300), .A2(G50), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n261), .B2(new_n298), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n394), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT11), .ZN(new_n416));
  OR2_X1    g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n415), .A2(new_n416), .ZN(new_n418));
  XNOR2_X1  g0218(.A(KEYINPUT75), .B(KEYINPUT12), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n360), .B2(new_n289), .ZN(new_n420));
  OR3_X1    g0220(.A1(new_n289), .A2(KEYINPUT12), .A3(G68), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n203), .B1(new_n208), .B2(G20), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n420), .A2(new_n421), .B1(new_n317), .B2(new_n422), .ZN(new_n423));
  AND3_X1   g0223(.A1(new_n417), .A2(new_n418), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n259), .A2(KEYINPUT74), .A3(G226), .ZN(new_n426));
  INV_X1    g0226(.A(G1698), .ZN(new_n427));
  OAI211_X1 g0227(.A(G226), .B(new_n427), .C1(new_n379), .C2(new_n380), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT74), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G97), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(new_n329), .B2(new_n427), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n268), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT13), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n270), .A2(G238), .A3(new_n271), .A4(new_n274), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n275), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n434), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n381), .A2(new_n240), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n440), .A2(G1698), .B1(G33), .B2(G97), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n426), .A2(new_n430), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n374), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT13), .B1(new_n443), .B2(new_n437), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n439), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT14), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(new_n446), .A3(G169), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n439), .A2(new_n444), .A3(G179), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n446), .B1(new_n445), .B2(G169), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n425), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n424), .B1(new_n445), .B2(new_n338), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n400), .B1(new_n439), .B2(new_n444), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n316), .A2(new_n411), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n208), .A2(G45), .ZN(new_n458));
  NOR2_X1   g0258(.A1(KEYINPUT5), .A2(G41), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(KEYINPUT5), .A2(G41), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n458), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n462), .A2(G274), .A3(new_n270), .A4(new_n274), .ZN(new_n463));
  INV_X1    g0263(.A(G45), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(G1), .ZN(new_n465));
  INV_X1    g0265(.A(new_n461), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n465), .B1(new_n466), .B2(new_n459), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n270), .A2(new_n467), .A3(G270), .A4(new_n274), .ZN(new_n468));
  AND2_X1   g0268(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g0269(.A(G264), .B(G1698), .C1(new_n379), .C2(new_n380), .ZN(new_n470));
  OAI211_X1 g0270(.A(G257), .B(new_n427), .C1(new_n379), .C2(new_n380), .ZN(new_n471));
  INV_X1    g0271(.A(G303), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n470), .B(new_n471), .C1(new_n472), .C2(new_n262), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n268), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT82), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G283), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n209), .ZN(new_n478));
  OR2_X1    g0278(.A1(KEYINPUT78), .A2(G97), .ZN(new_n479));
  NAND2_X1  g0279(.A1(KEYINPUT78), .A2(G97), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n478), .B1(new_n481), .B2(new_n256), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT20), .ZN(new_n483));
  INV_X1    g0283(.A(G116), .ZN(new_n484));
  AOI22_X1  g0284(.A1(KEYINPUT82), .A2(new_n483), .B1(new_n484), .B2(G20), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n394), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n476), .B(KEYINPUT20), .C1(new_n482), .C2(new_n486), .ZN(new_n487));
  AND2_X1   g0287(.A1(KEYINPUT78), .A2(G97), .ZN(new_n488));
  NOR2_X1   g0288(.A1(KEYINPUT78), .A2(G97), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n209), .B(new_n477), .C1(new_n490), .C2(G33), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n476), .A2(KEYINPUT20), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n491), .A2(new_n394), .A3(new_n485), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n289), .A2(new_n484), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n208), .A2(G33), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n289), .A2(new_n495), .A3(new_n229), .A4(new_n287), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n494), .B1(new_n497), .B2(new_n484), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n487), .A2(new_n493), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n475), .A2(new_n499), .A3(G169), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT21), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n469), .A2(G179), .A3(new_n474), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n500), .A2(new_n501), .B1(new_n502), .B2(new_n499), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT83), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(new_n500), .B2(new_n501), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n304), .B1(new_n469), .B2(new_n474), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n506), .A2(KEYINPUT83), .A3(KEYINPUT21), .A4(new_n499), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n503), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n270), .A2(new_n467), .A3(G264), .A4(new_n274), .ZN(new_n509));
  OAI211_X1 g0309(.A(G257), .B(G1698), .C1(new_n379), .C2(new_n380), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G294), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n259), .A2(KEYINPUT86), .A3(G250), .ZN(new_n513));
  OAI211_X1 g0313(.A(G250), .B(new_n427), .C1(new_n379), .C2(new_n380), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT86), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n512), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n463), .B(new_n509), .C1(new_n517), .C2(new_n374), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n304), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n510), .A2(new_n511), .ZN(new_n520));
  AOI21_X1  g0320(.A(KEYINPUT86), .B1(new_n259), .B2(G250), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n514), .A2(new_n515), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n268), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n524), .A2(new_n285), .A3(new_n463), .A4(new_n509), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT24), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n209), .B(G87), .C1(new_n379), .C2(new_n380), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT22), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT22), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n262), .A2(new_n529), .A3(new_n209), .A4(G87), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G33), .A2(G116), .ZN(new_n532));
  OR3_X1    g0332(.A1(new_n532), .A2(KEYINPUT84), .A3(G20), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT23), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n209), .B2(G107), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n330), .A2(KEYINPUT23), .A3(G20), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(KEYINPUT84), .B1(new_n532), .B2(G20), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n533), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n526), .B1(new_n531), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n531), .A2(new_n526), .A3(new_n539), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n288), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n323), .A2(new_n330), .ZN(new_n544));
  NOR2_X1   g0344(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n545));
  OR2_X1    g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AND2_X1   g0346(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n547), .B1(new_n544), .B2(new_n545), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n546), .A2(new_n548), .B1(G107), .B2(new_n497), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n519), .B(new_n525), .C1(new_n543), .C2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n508), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n542), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n394), .B1(new_n554), .B2(new_n540), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n518), .A2(G200), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n524), .A2(G190), .A3(new_n463), .A4(new_n509), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n555), .A2(new_n556), .A3(new_n557), .A4(new_n549), .ZN(new_n558));
  OAI211_X1 g0358(.A(G244), .B(new_n427), .C1(new_n379), .C2(new_n380), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT79), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT4), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n561), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n262), .A2(G244), .A3(new_n427), .A4(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n262), .A2(G250), .A3(G1698), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n562), .A2(new_n477), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n268), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n270), .A2(new_n467), .A3(G257), .A4(new_n274), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n463), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  AND3_X1   g0370(.A1(new_n567), .A2(G179), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n304), .B1(new_n567), .B2(new_n570), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n359), .A2(G107), .A3(new_n361), .ZN(new_n573));
  XOR2_X1   g0373(.A(G97), .B(G107), .Z(new_n574));
  NAND2_X1  g0374(.A1(new_n330), .A2(KEYINPUT6), .ZN(new_n575));
  OAI22_X1  g0375(.A1(new_n574), .A2(KEYINPUT6), .B1(new_n490), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n576), .A2(G20), .B1(G77), .B2(new_n300), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n288), .B1(new_n573), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(G97), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n323), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n496), .B2(new_n579), .ZN(new_n581));
  OAI22_X1  g0381(.A1(new_n571), .A2(new_n572), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n567), .A2(new_n570), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(G200), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n573), .A2(new_n577), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n581), .B1(new_n585), .B2(new_n394), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n569), .B1(new_n268), .B2(new_n566), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(G190), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n584), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n558), .A2(new_n582), .A3(new_n589), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n474), .A2(new_n468), .A3(new_n463), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n499), .B1(new_n591), .B2(G190), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(new_n400), .B2(new_n591), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT19), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n209), .B1(new_n432), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n479), .A2(new_n330), .A3(new_n480), .ZN(new_n596));
  XNOR2_X1  g0396(.A(KEYINPUT80), .B(G87), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n262), .A2(new_n209), .A3(G68), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n594), .B1(new_n490), .B2(new_n298), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT81), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT81), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n598), .A2(new_n600), .A3(new_n603), .A4(new_n599), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n602), .A2(new_n394), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n497), .A2(new_n320), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n320), .A2(new_n289), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(G244), .B(G1698), .C1(new_n379), .C2(new_n380), .ZN(new_n610));
  OAI211_X1 g0410(.A(G238), .B(new_n427), .C1(new_n379), .C2(new_n380), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(new_n611), .A3(new_n532), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n268), .ZN(new_n613));
  OR2_X1    g0413(.A1(new_n465), .A2(G250), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n458), .A2(G274), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n614), .A2(new_n615), .A3(new_n270), .A4(new_n274), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(G169), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n613), .A2(G179), .A3(new_n616), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n609), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n400), .B1(new_n613), .B2(new_n616), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n613), .A2(new_n616), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n622), .B1(G190), .B2(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n496), .A2(new_n382), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n624), .A2(new_n608), .A3(new_n605), .A4(new_n626), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n593), .A2(new_n621), .A3(new_n627), .ZN(new_n628));
  AND4_X1   g0428(.A1(new_n457), .A2(new_n553), .A3(new_n590), .A4(new_n628), .ZN(G372));
  INV_X1    g0429(.A(new_n306), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n388), .A2(new_n399), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n336), .A2(new_n454), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n445), .A2(G169), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT14), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n635), .A2(new_n448), .A3(new_n447), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n633), .B1(new_n425), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n408), .A2(new_n406), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n632), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n315), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n313), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n630), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n457), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n613), .A2(G179), .A3(new_n616), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n304), .B1(new_n613), .B2(new_n616), .ZN(new_n645));
  OAI21_X1  g0445(.A(KEYINPUT87), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT87), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n618), .A2(new_n647), .A3(new_n619), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n649), .A2(new_n609), .ZN(new_n650));
  INV_X1    g0450(.A(new_n586), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n567), .A2(G179), .A3(new_n570), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n304), .B2(new_n587), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n627), .A2(new_n621), .A3(new_n651), .A4(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n650), .B1(new_n654), .B2(KEYINPUT26), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT89), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n288), .B1(new_n601), .B2(KEYINPUT81), .ZN(new_n657));
  AOI211_X1 g0457(.A(new_n607), .B(new_n625), .C1(new_n657), .C2(new_n604), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n649), .A2(new_n609), .B1(new_n658), .B2(new_n624), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT26), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n652), .B(KEYINPUT88), .C1(new_n304), .C2(new_n587), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT88), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n586), .B1(new_n653), .B2(new_n662), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n659), .A2(new_n660), .A3(new_n661), .A4(new_n663), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n655), .A2(new_n656), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n656), .B1(new_n655), .B2(new_n664), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n551), .A2(new_n505), .A3(new_n503), .A4(new_n507), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n590), .A2(new_n667), .A3(new_n659), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n665), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n642), .B1(new_n643), .B2(new_n669), .ZN(G369));
  NAND3_X1  g0470(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(G213), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(G343), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n499), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g0477(.A(new_n508), .B(new_n677), .Z(new_n678));
  AND2_X1   g0478(.A1(new_n678), .A2(new_n593), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n679), .A2(G330), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n551), .A2(new_n676), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n676), .B1(new_n543), .B2(new_n550), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n558), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n681), .B1(new_n551), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT90), .ZN(new_n686));
  INV_X1    g0486(.A(new_n508), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(new_n676), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n551), .B2(new_n676), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n686), .A2(new_n690), .ZN(G399));
  NOR2_X1   g0491(.A1(new_n212), .A2(G41), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G1), .ZN(new_n694));
  OR3_X1    g0494(.A1(new_n596), .A2(new_n597), .A3(G116), .ZN(new_n695));
  OAI22_X1  g0495(.A1(new_n694), .A2(new_n695), .B1(new_n236), .B2(new_n693), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n696), .B(KEYINPUT28), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n663), .A2(new_n661), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n660), .B1(new_n698), .B2(new_n659), .ZN(new_n699));
  INV_X1    g0499(.A(new_n650), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n654), .B2(KEYINPUT26), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n687), .A2(KEYINPUT91), .A3(new_n551), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT91), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n667), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n703), .A2(new_n705), .A3(new_n590), .A4(new_n659), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n676), .B1(new_n702), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(KEYINPUT29), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n669), .A2(new_n676), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n708), .B1(new_n709), .B2(KEYINPUT29), .ZN(new_n710));
  INV_X1    g0510(.A(new_n676), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n553), .A2(new_n590), .A3(new_n628), .A4(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT30), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n591), .A2(new_n509), .A3(new_n524), .A4(new_n623), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(new_n652), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n591), .A2(G179), .A3(new_n623), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(new_n518), .A3(new_n583), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n524), .A2(new_n509), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n475), .A2(new_n617), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n718), .A2(new_n571), .A3(new_n719), .A4(KEYINPUT30), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n715), .A2(new_n717), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n676), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT31), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n721), .A2(KEYINPUT31), .A3(new_n676), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n712), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G330), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n710), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n697), .B1(new_n728), .B2(G1), .ZN(G364));
  NOR2_X1   g0529(.A1(new_n211), .A2(G20), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n208), .B1(new_n730), .B2(G45), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n692), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n680), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n679), .A2(G330), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G13), .A2(G33), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n679), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n212), .A2(new_n381), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G355), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(G116), .B2(new_n213), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n237), .A2(new_n464), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n212), .A2(new_n262), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n747), .B1(new_n253), .B2(G45), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n744), .B1(new_n745), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n209), .B1(KEYINPUT92), .B2(new_n304), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n304), .A2(KEYINPUT92), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n229), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n739), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n733), .B1(new_n749), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n209), .A2(new_n285), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n756), .A2(G190), .A3(G200), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT93), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n209), .A2(G179), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(G190), .A3(G200), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT94), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n762), .A2(G326), .B1(new_n769), .B2(G303), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G190), .A2(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n756), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G311), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n763), .A2(new_n771), .ZN(new_n774));
  INV_X1    g0574(.A(G329), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n772), .A2(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n756), .A2(G190), .A3(new_n400), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n262), .B(new_n776), .C1(G322), .C2(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n763), .A2(new_n338), .A3(G200), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G283), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n338), .A2(G179), .A3(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n209), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(KEYINPUT33), .B(G317), .ZN(new_n786));
  NOR4_X1   g0586(.A1(new_n209), .A2(new_n285), .A3(new_n400), .A4(G190), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n785), .A2(G294), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n770), .A2(new_n779), .A3(new_n782), .A4(new_n788), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n777), .A2(new_n202), .B1(new_n772), .B2(new_n261), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n785), .A2(G97), .B1(G68), .B2(new_n787), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT32), .ZN(new_n792));
  INV_X1    g0592(.A(G159), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n774), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n791), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n790), .B(new_n795), .C1(new_n792), .C2(new_n794), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(new_n233), .B2(new_n761), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n781), .A2(G107), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(new_n262), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(new_n769), .B2(new_n597), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT95), .Z(new_n801));
  OAI21_X1  g0601(.A(new_n789), .B1(new_n797), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n755), .B1(new_n802), .B2(new_n752), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n734), .A2(new_n736), .B1(new_n741), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(G396));
  NOR2_X1   g0605(.A1(new_n336), .A2(new_n676), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n339), .B1(new_n327), .B2(new_n711), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n806), .B1(new_n807), .B2(new_n336), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n340), .A2(new_n711), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n709), .A2(new_n808), .B1(new_n669), .B2(new_n809), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n810), .A2(new_n727), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n733), .B1(new_n810), .B2(new_n727), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n381), .B1(new_n768), .B2(new_n330), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT96), .ZN(new_n815));
  INV_X1    g0615(.A(G294), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n784), .A2(new_n579), .B1(new_n777), .B2(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT97), .ZN(new_n818));
  INV_X1    g0618(.A(new_n772), .ZN(new_n819));
  INV_X1    g0619(.A(new_n774), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G116), .A2(new_n819), .B1(new_n820), .B2(G311), .ZN(new_n821));
  INV_X1    g0621(.A(G283), .ZN(new_n822));
  INV_X1    g0622(.A(new_n787), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n821), .B1(new_n382), .B2(new_n780), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(G303), .B2(new_n762), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n815), .A2(new_n818), .A3(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(KEYINPUT98), .B(G143), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n778), .A2(new_n828), .B1(new_n819), .B2(G159), .ZN(new_n829));
  INV_X1    g0629(.A(G150), .ZN(new_n830));
  INV_X1    g0630(.A(G137), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n829), .B1(new_n830), .B2(new_n823), .C1(new_n761), .C2(new_n831), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT99), .Z(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(KEYINPUT34), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n381), .B1(new_n820), .B2(G132), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT100), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n769), .A2(G50), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n780), .A2(new_n203), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(G58), .B2(new_n785), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n834), .A2(new_n836), .A3(new_n837), .A4(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n833), .A2(KEYINPUT34), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n826), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n752), .ZN(new_n843));
  INV_X1    g0643(.A(new_n733), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n752), .A2(new_n737), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n844), .B1(new_n845), .B2(new_n261), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n808), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n847), .B1(new_n737), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n813), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(G384));
  OR2_X1    g0651(.A1(new_n576), .A2(KEYINPUT35), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n576), .A2(KEYINPUT35), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n852), .A2(G116), .A3(new_n232), .A4(new_n853), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT36), .Z(new_n855));
  OAI21_X1  g0655(.A(G77), .B1(new_n218), .B2(new_n202), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n236), .A2(new_n856), .B1(G50), .B2(new_n203), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n208), .A2(G13), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n855), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n425), .A2(new_n676), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n451), .A2(new_n455), .A3(new_n860), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n425), .B(new_n676), .C1(new_n636), .C2(new_n454), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n655), .A2(new_n664), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n668), .B1(new_n864), .B2(KEYINPUT89), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n655), .A2(new_n656), .A3(new_n664), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n809), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n863), .B1(new_n867), .B2(new_n806), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n358), .B1(KEYINPUT16), .B2(new_n357), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n674), .B1(new_n869), .B2(new_n389), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n409), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT101), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n409), .A2(KEYINPUT101), .A3(new_n870), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n368), .A2(new_n674), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT37), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n397), .A2(new_n386), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n877), .A2(new_n878), .A3(new_n879), .A4(new_n404), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n869), .A2(new_n389), .B1(new_n387), .B2(new_n674), .ZN(new_n881));
  INV_X1    g0681(.A(new_n404), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT37), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT38), .B1(new_n875), .B2(new_n884), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n409), .A2(KEYINPUT101), .A3(new_n870), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT101), .B1(new_n409), .B2(new_n870), .ZN(new_n887));
  OAI211_X1 g0687(.A(KEYINPUT38), .B(new_n884), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n674), .ZN(new_n891));
  OAI22_X1  g0691(.A1(new_n868), .A2(new_n890), .B1(new_n632), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n884), .B1(new_n886), .B2(new_n887), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n895), .A2(KEYINPUT39), .A3(new_n888), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n410), .A2(new_n877), .ZN(new_n898));
  INV_X1    g0698(.A(new_n880), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n387), .B1(new_n407), .B2(new_n389), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT102), .B1(new_n900), .B2(new_n882), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT102), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n879), .A2(new_n902), .A3(new_n404), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n901), .A2(new_n877), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT37), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n899), .B1(new_n905), .B2(KEYINPUT103), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT103), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n904), .A2(new_n907), .A3(KEYINPUT37), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n898), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n888), .B1(new_n909), .B2(KEYINPUT38), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n896), .B1(new_n897), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n636), .A2(new_n425), .A3(new_n711), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n892), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n457), .B(new_n708), .C1(new_n709), .C2(KEYINPUT29), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n915), .A2(new_n642), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n914), .B(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n457), .A2(new_n726), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n918), .B(KEYINPUT104), .Z(new_n919));
  INV_X1    g0719(.A(new_n898), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n879), .A2(new_n404), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n876), .B1(new_n921), .B2(KEYINPUT102), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n878), .B1(new_n922), .B2(new_n903), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n880), .B1(new_n923), .B2(new_n907), .ZN(new_n924));
  INV_X1    g0724(.A(new_n908), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n920), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n889), .B1(new_n926), .B2(new_n894), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n863), .A2(new_n726), .A3(new_n808), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(KEYINPUT40), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n863), .A2(new_n726), .A3(new_n808), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n895), .B2(new_n888), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n927), .A2(new_n929), .B1(new_n931), .B2(KEYINPUT40), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n919), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n919), .A2(new_n932), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n933), .A2(G330), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n917), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n208), .B2(new_n730), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n917), .A2(new_n935), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n859), .B1(new_n937), .B2(new_n938), .ZN(G367));
  INV_X1    g0739(.A(new_n728), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n698), .A2(new_n676), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n582), .B(new_n589), .C1(new_n586), .C2(new_n711), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n690), .A2(new_n943), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT44), .Z(new_n945));
  NOR2_X1   g0745(.A1(new_n690), .A2(new_n943), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT45), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n686), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n686), .A2(new_n948), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n684), .B(new_n688), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n680), .B(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n940), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n692), .B(KEYINPUT41), .Z(new_n956));
  OAI21_X1  g0756(.A(new_n731), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n943), .A2(new_n689), .ZN(new_n958));
  XOR2_X1   g0758(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n959));
  OR2_X1    g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n959), .ZN(new_n961));
  INV_X1    g0761(.A(new_n943), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n962), .A2(new_n552), .B1(new_n651), .B2(new_n653), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n960), .B(new_n961), .C1(new_n676), .C2(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT106), .ZN(new_n965));
  OR3_X1    g0765(.A1(new_n700), .A2(new_n658), .A3(new_n711), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n659), .B1(new_n658), .B2(new_n711), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(KEYINPUT43), .Z(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n965), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n965), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n686), .A2(new_n962), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n957), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n246), .A2(new_n747), .ZN(new_n978));
  INV_X1    g0778(.A(new_n320), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n753), .B1(new_n213), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n733), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n823), .A2(new_n816), .B1(new_n780), .B2(new_n490), .ZN(new_n982));
  AOI22_X1  g0782(.A1(G283), .A2(new_n819), .B1(new_n820), .B2(G317), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n983), .B(new_n381), .C1(new_n472), .C2(new_n777), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n982), .B(new_n984), .C1(G107), .C2(new_n785), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n773), .B2(new_n761), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n768), .A2(new_n484), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT46), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n785), .A2(G68), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n989), .B1(new_n830), .B2(new_n777), .C1(new_n761), .C2(new_n827), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(KEYINPUT107), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n262), .B1(new_n772), .B2(new_n233), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n823), .A2(new_n793), .B1(new_n261), .B2(new_n780), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(G137), .C2(new_n820), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n991), .B(new_n994), .C1(new_n202), .C2(new_n768), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n990), .A2(KEYINPUT107), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n986), .A2(new_n988), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT47), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n981), .B1(new_n998), .B2(new_n752), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n966), .A2(new_n739), .A3(new_n967), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n977), .A2(new_n1001), .ZN(G387));
  OR2_X1    g0802(.A1(new_n243), .A2(new_n464), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n1003), .A2(new_n746), .B1(new_n695), .B2(new_n742), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n297), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1005), .A2(G50), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT50), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n464), .B1(new_n203), .B2(new_n261), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n695), .B(new_n1008), .C1(new_n1007), .C2(new_n1006), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n1004), .A2(new_n1009), .B1(G107), .B2(new_n213), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n844), .B1(new_n1010), .B2(new_n753), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n769), .A2(G77), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n793), .B2(new_n761), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n778), .A2(G50), .B1(new_n820), .B2(G150), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1014), .B(new_n262), .C1(new_n203), .C2(new_n772), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n785), .A2(new_n320), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n579), .B2(new_n780), .C1(new_n1005), .C2(new_n823), .ZN(new_n1017));
  NOR3_X1   g0817(.A1(new_n1013), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(G326), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n381), .B1(new_n774), .B2(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n778), .A2(G317), .B1(new_n819), .B2(G303), .ZN(new_n1021));
  INV_X1    g0821(.A(G322), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1021), .B1(new_n773), .B2(new_n823), .C1(new_n761), .C2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT48), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n769), .A2(G294), .B1(G283), .B2(new_n785), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT49), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n1020), .B(new_n1030), .C1(G116), .C2(new_n781), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1018), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n752), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1011), .B1(new_n684), .B2(new_n740), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT108), .Z(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n954), .B2(new_n732), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n728), .A2(new_n954), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n692), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n728), .A2(new_n954), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1037), .B1(new_n1039), .B2(new_n1040), .ZN(G393));
  INV_X1    g0841(.A(KEYINPUT109), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n949), .A2(new_n1042), .A3(new_n950), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n686), .A2(KEYINPUT109), .A3(new_n948), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n732), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n762), .A2(G317), .B1(G311), .B2(new_n778), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT52), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n768), .A2(new_n822), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n381), .B1(new_n774), .B2(new_n1022), .C1(new_n816), .C2(new_n772), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n798), .B1(new_n484), .B2(new_n784), .C1(new_n472), .C2(new_n823), .ZN(new_n1051));
  NOR4_X1   g0851(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT112), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n761), .A2(new_n830), .B1(new_n793), .B2(new_n777), .ZN(new_n1054));
  XOR2_X1   g0854(.A(KEYINPUT110), .B(KEYINPUT51), .Z(new_n1055));
  XNOR2_X1  g0855(.A(new_n1054), .B(new_n1055), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n262), .B1(new_n774), .B2(new_n827), .C1(new_n1005), .C2(new_n772), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n785), .A2(G77), .B1(new_n781), .B2(G87), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n233), .B2(new_n823), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1057), .B(new_n1059), .C1(new_n360), .C2(new_n769), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT111), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1034), .B1(new_n1053), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n250), .A2(new_n746), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n754), .B1(new_n212), .B2(new_n481), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n844), .B(new_n1063), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n943), .A2(new_n739), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1043), .A2(new_n1038), .A3(new_n1044), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n692), .B1(new_n951), .B2(new_n1038), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1046), .B(new_n1068), .C1(new_n1070), .C2(new_n1071), .ZN(G390));
  NAND4_X1  g0872(.A1(new_n863), .A2(new_n726), .A3(new_n808), .A4(G330), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n806), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n669), .B2(new_n809), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n913), .B1(new_n1076), .B2(new_n863), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n905), .A2(KEYINPUT103), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1078), .A2(new_n880), .A3(new_n908), .ZN(new_n1079));
  AOI21_X1  g0879(.A(KEYINPUT38), .B1(new_n1079), .B2(new_n920), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n897), .B1(new_n1080), .B2(new_n889), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n896), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1077), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n863), .B(KEYINPUT113), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n336), .A2(new_n807), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n806), .B1(new_n707), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n912), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1087), .A2(new_n927), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1074), .B1(new_n1083), .B2(new_n1088), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n910), .B(new_n912), .C1(new_n1086), .C2(new_n1084), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1090), .B(new_n1073), .C1(new_n911), .C2(new_n1077), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1086), .A2(new_n1073), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1084), .B1(new_n727), .B2(new_n848), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n861), .B(new_n862), .C1(new_n727), .C2(new_n848), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n1073), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n1093), .A2(new_n1094), .B1(new_n1096), .B2(new_n1076), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n457), .A2(G330), .A3(new_n726), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n915), .A2(new_n642), .A3(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n693), .B1(new_n1092), .B2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1089), .A2(new_n1091), .A3(new_n1100), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1089), .A2(new_n732), .A3(new_n1091), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n844), .B1(new_n845), .B2(new_n1005), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n481), .A2(new_n819), .B1(new_n787), .B2(G107), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n761), .B2(new_n822), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT116), .Z(new_n1109));
  OAI22_X1  g0909(.A1(new_n784), .A2(new_n261), .B1(new_n777), .B2(new_n484), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT118), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n838), .B(new_n1111), .C1(G294), .C2(new_n820), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n381), .B1(new_n768), .B2(new_n382), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n1113), .A2(KEYINPUT117), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(KEYINPUT117), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1109), .A2(new_n1112), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n785), .A2(G159), .B1(G137), .B2(new_n787), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(KEYINPUT54), .B(G143), .ZN(new_n1118));
  XOR2_X1   g0918(.A(new_n1118), .B(KEYINPUT114), .Z(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1117), .B1(new_n1120), .B2(new_n772), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT115), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n768), .A2(new_n830), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT53), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n381), .B1(new_n778), .B2(G132), .ZN(new_n1125));
  INV_X1    g0925(.A(G125), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1125), .B1(new_n233), .B2(new_n780), .C1(new_n1126), .C2(new_n774), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(G128), .B2(new_n762), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1122), .A2(new_n1124), .A3(new_n1128), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1116), .A2(new_n1129), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1106), .B1(new_n1034), .B2(new_n1130), .C1(new_n911), .C2(new_n738), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1104), .A2(new_n1105), .A3(new_n1131), .ZN(G378));
  XNOR2_X1  g0932(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n303), .A2(new_n891), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n316), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1135), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(new_n641), .B2(new_n306), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1134), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n316), .A2(new_n1135), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n641), .A2(new_n306), .A3(new_n1137), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1140), .A2(new_n1141), .A3(new_n1133), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(G330), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1144), .B1(new_n932), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n928), .B1(new_n885), .B2(new_n889), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT40), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n930), .A2(new_n1148), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n1080), .B2(new_n889), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1149), .A2(new_n1151), .A3(new_n1143), .A4(G330), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n914), .A2(new_n1146), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1081), .A2(new_n1082), .A3(new_n913), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n892), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n1146), .A2(new_n1152), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n732), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n262), .A2(G41), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n989), .B1(new_n761), .B2(new_n484), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT120), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n823), .A2(new_n579), .B1(new_n979), .B2(new_n772), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT119), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1158), .B1(new_n822), .B2(new_n774), .C1(new_n330), .C2(new_n777), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(G58), .B2(new_n781), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1162), .A2(new_n1012), .A3(new_n1164), .A4(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT58), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1160), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n784), .A2(new_n830), .ZN(new_n1170));
  INV_X1    g0970(.A(G128), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n777), .A2(new_n1171), .B1(new_n772), .B2(new_n831), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1170), .B(new_n1172), .C1(G132), .C2(new_n787), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1173), .B1(new_n1126), .B2(new_n761), .C1(new_n768), .C2(new_n1120), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1174), .A2(KEYINPUT59), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(KEYINPUT59), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n781), .A2(G159), .ZN(new_n1177));
  AOI211_X1 g0977(.A(G33), .B(G41), .C1(new_n820), .C2(G124), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1169), .B1(new_n1168), .B2(new_n1167), .C1(new_n1175), .C2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n752), .ZN(new_n1181));
  XOR2_X1   g0981(.A(new_n1181), .B(KEYINPUT121), .Z(new_n1182));
  AOI21_X1  g0982(.A(new_n844), .B1(new_n845), .B2(new_n233), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1182), .B(new_n1183), .C1(new_n738), .C2(new_n1143), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n1157), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT57), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1155), .A2(new_n1154), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n910), .A2(new_n1150), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1143), .B1(new_n1188), .B2(G330), .ZN(new_n1189));
  AND4_X1   g0989(.A1(G330), .A2(new_n1149), .A3(new_n1151), .A4(new_n1143), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1187), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n914), .A2(new_n1146), .A3(new_n1152), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1186), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1099), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1103), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(new_n692), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1198));
  AOI21_X1  g0998(.A(KEYINPUT57), .B1(new_n1195), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1185), .B1(new_n1197), .B2(new_n1199), .ZN(G375));
  INV_X1    g1000(.A(new_n956), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1101), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n1084), .A2(new_n737), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n844), .B1(new_n845), .B2(new_n203), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n768), .A2(new_n579), .B1(new_n472), .B2(new_n774), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT122), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n381), .B1(new_n772), .B2(new_n330), .C1(new_n822), .C2(new_n777), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1016), .B1(new_n261), .B2(new_n780), .C1(new_n484), .C2(new_n823), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1208), .B(new_n1209), .C1(G294), .C2(new_n762), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n784), .A2(new_n233), .B1(new_n780), .B2(new_n202), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n381), .B1(new_n820), .B2(G128), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1212), .B1(new_n831), .B2(new_n777), .C1(new_n830), .C2(new_n772), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1211), .B(new_n1213), .C1(new_n787), .C2(new_n1119), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n762), .A2(G132), .B1(new_n769), .B2(G159), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1207), .A2(new_n1210), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1205), .B1(new_n1216), .B2(new_n1034), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n1097), .A2(new_n731), .B1(new_n1204), .B2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1203), .A2(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT123), .ZN(G381));
  OAI211_X1 g1021(.A(new_n1069), .B(new_n692), .C1(new_n1038), .C2(new_n951), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1045), .A2(new_n732), .B1(new_n1067), .B2(new_n1066), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1037), .B(new_n804), .C1(new_n1040), .C2(new_n1039), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1222), .A2(new_n850), .A3(new_n1223), .A4(new_n1225), .ZN(new_n1226));
  NOR3_X1   g1026(.A1(G387), .A2(G381), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1105), .A2(new_n1131), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1229));
  INV_X1    g1029(.A(G375), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1227), .A2(new_n1229), .A3(new_n1230), .ZN(G407));
  INV_X1    g1031(.A(G213), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1232), .A2(G343), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(G375), .A2(G378), .A3(new_n1234), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1235), .B(KEYINPUT124), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1236), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1037(.A(KEYINPUT125), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1103), .A2(new_n1194), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1201), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1238), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n956), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1242), .A2(KEYINPUT125), .A3(new_n1195), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1241), .A2(new_n1185), .A3(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1229), .ZN(new_n1245));
  OAI211_X1 g1045(.A(G378), .B(new_n1185), .C1(new_n1197), .C2(new_n1199), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1233), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1097), .A2(KEYINPUT60), .A3(new_n1099), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1248), .A2(new_n692), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT60), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1202), .B1(new_n1100), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1219), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n850), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1252), .A2(G384), .A3(new_n1219), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  AOI211_X1 g1056(.A(KEYINPUT126), .B(KEYINPUT63), .C1(new_n1247), .C2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT126), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1157), .A2(new_n1184), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1199), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n693), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n1259), .B(new_n1229), .C1(new_n1260), .C2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT125), .B1(new_n1242), .B2(new_n1195), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1263), .A2(new_n1259), .ZN(new_n1264));
  AOI21_X1  g1064(.A(G378), .B1(new_n1264), .B2(new_n1243), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1234), .B(new_n1256), .C1(new_n1262), .C2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT63), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1258), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1257), .A2(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1234), .B1(new_n1262), .B2(new_n1265), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1233), .A2(G2897), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(new_n1256), .B(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(KEYINPUT61), .B1(new_n1270), .B2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1247), .A2(KEYINPUT63), .A3(new_n1256), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n957), .A2(new_n976), .B1(new_n1000), .B2(new_n999), .ZN(new_n1275));
  AND2_X1   g1075(.A1(G393), .A2(G396), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1276), .A2(new_n1225), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(G390), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1222), .B(new_n1223), .C1(new_n1276), .C2(new_n1225), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1275), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1275), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1273), .A2(new_n1274), .A3(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT61), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(new_n1286), .B(new_n1271), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1285), .B1(new_n1247), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT62), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1266), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1247), .A2(KEYINPUT62), .A3(new_n1256), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1288), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT127), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1293), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(G387), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1296), .A2(KEYINPUT127), .A3(new_n1280), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1294), .A2(new_n1297), .ZN(new_n1298));
  OAI22_X1  g1098(.A1(new_n1269), .A2(new_n1284), .B1(new_n1292), .B2(new_n1298), .ZN(G405));
  NAND2_X1  g1099(.A1(G375), .A2(new_n1229), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1246), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1301), .B(new_n1286), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(new_n1302), .B(new_n1283), .ZN(G402));
endmodule


