

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582;

  XNOR2_X1 U323 ( .A(KEYINPUT54), .B(KEYINPUT118), .ZN(n409) );
  XOR2_X1 U324 ( .A(n385), .B(KEYINPUT32), .Z(n291) );
  XOR2_X1 U325 ( .A(n393), .B(n392), .Z(n292) );
  XNOR2_X1 U326 ( .A(KEYINPUT109), .B(KEYINPUT47), .ZN(n400) );
  XNOR2_X1 U327 ( .A(n401), .B(n400), .ZN(n406) );
  XNOR2_X1 U328 ( .A(n394), .B(n292), .ZN(n395) );
  XNOR2_X1 U329 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U330 ( .A(n396), .B(n395), .ZN(n572) );
  INV_X1 U331 ( .A(G190GAT), .ZN(n449) );
  XOR2_X1 U332 ( .A(KEYINPUT98), .B(n458), .Z(n533) );
  XNOR2_X1 U333 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U334 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XOR2_X1 U335 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n294) );
  XNOR2_X1 U336 ( .A(G92GAT), .B(KEYINPUT9), .ZN(n293) );
  XNOR2_X1 U337 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U338 ( .A(G134GAT), .B(KEYINPUT77), .Z(n314) );
  XOR2_X1 U339 ( .A(n295), .B(n314), .Z(n297) );
  XNOR2_X1 U340 ( .A(G218GAT), .B(G106GAT), .ZN(n296) );
  XNOR2_X1 U341 ( .A(n297), .B(n296), .ZN(n302) );
  XNOR2_X1 U342 ( .A(G99GAT), .B(G85GAT), .ZN(n298) );
  XNOR2_X1 U343 ( .A(n298), .B(KEYINPUT74), .ZN(n391) );
  XOR2_X1 U344 ( .A(KEYINPUT78), .B(n391), .Z(n300) );
  NAND2_X1 U345 ( .A1(G232GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U347 ( .A(n302), .B(n301), .Z(n312) );
  XOR2_X1 U348 ( .A(G43GAT), .B(G29GAT), .Z(n304) );
  XNOR2_X1 U349 ( .A(KEYINPUT7), .B(G50GAT), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U351 ( .A(n305), .B(KEYINPUT68), .Z(n307) );
  XNOR2_X1 U352 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n306) );
  XNOR2_X1 U353 ( .A(n307), .B(n306), .ZN(n382) );
  XOR2_X1 U354 ( .A(KEYINPUT76), .B(KEYINPUT75), .Z(n309) );
  XNOR2_X1 U355 ( .A(G190GAT), .B(G162GAT), .ZN(n308) );
  XNOR2_X1 U356 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U357 ( .A(n382), .B(n310), .ZN(n311) );
  XOR2_X1 U358 ( .A(n312), .B(n311), .Z(n527) );
  XNOR2_X1 U359 ( .A(G1GAT), .B(G127GAT), .ZN(n313) );
  XNOR2_X1 U360 ( .A(n313), .B(G57GAT), .ZN(n357) );
  XOR2_X1 U361 ( .A(n357), .B(n314), .Z(n316) );
  NAND2_X1 U362 ( .A1(G225GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U363 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U364 ( .A(n317), .B(KEYINPUT6), .Z(n320) );
  XNOR2_X1 U365 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n318) );
  XNOR2_X1 U366 ( .A(n318), .B(G120GAT), .ZN(n438) );
  XNOR2_X1 U367 ( .A(n438), .B(KEYINPUT4), .ZN(n319) );
  XNOR2_X1 U368 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U369 ( .A(KEYINPUT96), .B(G85GAT), .Z(n322) );
  XNOR2_X1 U370 ( .A(G29GAT), .B(G148GAT), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U372 ( .A(n324), .B(n323), .Z(n334) );
  XOR2_X1 U373 ( .A(KEYINPUT3), .B(KEYINPUT94), .Z(n326) );
  XNOR2_X1 U374 ( .A(G162GAT), .B(KEYINPUT93), .ZN(n325) );
  XNOR2_X1 U375 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U376 ( .A(n327), .B(KEYINPUT2), .Z(n329) );
  XNOR2_X1 U377 ( .A(G141GAT), .B(G155GAT), .ZN(n328) );
  XNOR2_X1 U378 ( .A(n329), .B(n328), .ZN(n426) );
  XOR2_X1 U379 ( .A(KEYINPUT5), .B(KEYINPUT95), .Z(n331) );
  XNOR2_X1 U380 ( .A(KEYINPUT1), .B(KEYINPUT97), .ZN(n330) );
  XNOR2_X1 U381 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U382 ( .A(n426), .B(n332), .ZN(n333) );
  XNOR2_X1 U383 ( .A(n334), .B(n333), .ZN(n458) );
  INV_X1 U384 ( .A(n533), .ZN(n478) );
  XNOR2_X1 U385 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n335) );
  XNOR2_X1 U386 ( .A(n335), .B(KEYINPUT86), .ZN(n336) );
  XOR2_X1 U387 ( .A(n336), .B(KEYINPUT87), .Z(n338) );
  XNOR2_X1 U388 ( .A(KEYINPUT19), .B(G190GAT), .ZN(n337) );
  XNOR2_X1 U389 ( .A(n338), .B(n337), .ZN(n439) );
  XOR2_X1 U390 ( .A(G64GAT), .B(G92GAT), .Z(n340) );
  XNOR2_X1 U391 ( .A(G176GAT), .B(G204GAT), .ZN(n339) );
  XNOR2_X1 U392 ( .A(n340), .B(n339), .ZN(n386) );
  XOR2_X1 U393 ( .A(G169GAT), .B(G8GAT), .Z(n372) );
  XOR2_X1 U394 ( .A(n386), .B(n372), .Z(n342) );
  NAND2_X1 U395 ( .A1(G226GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U396 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U397 ( .A(n343), .B(KEYINPUT99), .Z(n345) );
  XOR2_X1 U398 ( .A(G183GAT), .B(G211GAT), .Z(n364) );
  XNOR2_X1 U399 ( .A(G36GAT), .B(n364), .ZN(n344) );
  XNOR2_X1 U400 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U401 ( .A(n439), .B(n346), .ZN(n350) );
  XOR2_X1 U402 ( .A(KEYINPUT21), .B(G218GAT), .Z(n348) );
  XNOR2_X1 U403 ( .A(KEYINPUT92), .B(KEYINPUT91), .ZN(n347) );
  XNOR2_X1 U404 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U405 ( .A(G197GAT), .B(n349), .Z(n422) );
  XOR2_X1 U406 ( .A(n350), .B(n422), .Z(n482) );
  XNOR2_X1 U407 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n408) );
  XOR2_X1 U408 ( .A(KEYINPUT12), .B(KEYINPUT79), .Z(n352) );
  XNOR2_X1 U409 ( .A(KEYINPUT80), .B(KEYINPUT14), .ZN(n351) );
  XNOR2_X1 U410 ( .A(n352), .B(n351), .ZN(n368) );
  XOR2_X1 U411 ( .A(KEYINPUT81), .B(KEYINPUT15), .Z(n354) );
  NAND2_X1 U412 ( .A1(G231GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U414 ( .A(n355), .B(KEYINPUT82), .Z(n359) );
  XNOR2_X1 U415 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n356) );
  XNOR2_X1 U416 ( .A(n356), .B(KEYINPUT70), .ZN(n387) );
  XNOR2_X1 U417 ( .A(n357), .B(n387), .ZN(n358) );
  XNOR2_X1 U418 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U419 ( .A(G64GAT), .B(G78GAT), .Z(n361) );
  XNOR2_X1 U420 ( .A(G8GAT), .B(G155GAT), .ZN(n360) );
  XNOR2_X1 U421 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U422 ( .A(n363), .B(n362), .Z(n366) );
  XOR2_X1 U423 ( .A(G15GAT), .B(G22GAT), .Z(n377) );
  XNOR2_X1 U424 ( .A(n377), .B(n364), .ZN(n365) );
  XNOR2_X1 U425 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U426 ( .A(n368), .B(n367), .ZN(n543) );
  XOR2_X1 U427 ( .A(KEYINPUT108), .B(n543), .Z(n560) );
  INV_X1 U428 ( .A(n527), .ZN(n546) );
  XOR2_X1 U429 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n370) );
  XNOR2_X1 U430 ( .A(G197GAT), .B(G1GAT), .ZN(n369) );
  XNOR2_X1 U431 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U432 ( .A(n371), .B(KEYINPUT29), .ZN(n376) );
  XOR2_X1 U433 ( .A(KEYINPUT66), .B(n372), .Z(n374) );
  NAND2_X1 U434 ( .A1(G229GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U435 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U436 ( .A(n376), .B(n375), .ZN(n378) );
  XOR2_X1 U437 ( .A(n378), .B(n377), .Z(n380) );
  XNOR2_X1 U438 ( .A(G113GAT), .B(G141GAT), .ZN(n379) );
  XNOR2_X1 U439 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U440 ( .A(n382), .B(n381), .ZN(n566) );
  XOR2_X1 U441 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n384) );
  NAND2_X1 U442 ( .A1(G230GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U443 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U444 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U445 ( .A(n291), .B(n388), .ZN(n396) );
  XOR2_X1 U446 ( .A(G78GAT), .B(G148GAT), .Z(n390) );
  XNOR2_X1 U447 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n390), .B(n389), .ZN(n418) );
  XNOR2_X1 U449 ( .A(n418), .B(n391), .ZN(n394) );
  XOR2_X1 U450 ( .A(KEYINPUT71), .B(KEYINPUT72), .Z(n393) );
  XNOR2_X1 U451 ( .A(G120GAT), .B(G57GAT), .ZN(n392) );
  XOR2_X1 U452 ( .A(KEYINPUT41), .B(n572), .Z(n538) );
  INV_X1 U453 ( .A(n538), .ZN(n553) );
  NOR2_X1 U454 ( .A1(n566), .A2(n553), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n397), .B(KEYINPUT46), .ZN(n398) );
  NOR2_X1 U456 ( .A1(n546), .A2(n398), .ZN(n399) );
  NAND2_X1 U457 ( .A1(n560), .A2(n399), .ZN(n401) );
  INV_X1 U458 ( .A(n543), .ZN(n577) );
  XNOR2_X1 U459 ( .A(n527), .B(KEYINPUT36), .ZN(n580) );
  NOR2_X1 U460 ( .A1(n577), .A2(n580), .ZN(n402) );
  XOR2_X1 U461 ( .A(KEYINPUT45), .B(n402), .Z(n403) );
  NOR2_X1 U462 ( .A1(n572), .A2(n403), .ZN(n404) );
  XOR2_X1 U463 ( .A(n566), .B(KEYINPUT69), .Z(n550) );
  NAND2_X1 U464 ( .A1(n404), .A2(n550), .ZN(n405) );
  NAND2_X1 U465 ( .A1(n406), .A2(n405), .ZN(n407) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n530) );
  NAND2_X1 U467 ( .A1(n482), .A2(n530), .ZN(n410) );
  NOR2_X1 U468 ( .A1(n478), .A2(n411), .ZN(n565) );
  XOR2_X1 U469 ( .A(KEYINPUT23), .B(KEYINPUT75), .Z(n413) );
  XNOR2_X1 U470 ( .A(G50GAT), .B(G22GAT), .ZN(n412) );
  XNOR2_X1 U471 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U472 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n415) );
  XNOR2_X1 U473 ( .A(KEYINPUT22), .B(G211GAT), .ZN(n414) );
  XNOR2_X1 U474 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U475 ( .A(n417), .B(n416), .Z(n424) );
  XOR2_X1 U476 ( .A(n418), .B(G204GAT), .Z(n420) );
  NAND2_X1 U477 ( .A1(G228GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U478 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U479 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U480 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n459) );
  NAND2_X1 U482 ( .A1(n565), .A2(n459), .ZN(n427) );
  XNOR2_X1 U483 ( .A(KEYINPUT55), .B(n427), .ZN(n448) );
  XOR2_X1 U484 ( .A(G176GAT), .B(G71GAT), .Z(n429) );
  XNOR2_X1 U485 ( .A(G169GAT), .B(G183GAT), .ZN(n428) );
  XNOR2_X1 U486 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U487 ( .A(KEYINPUT84), .B(KEYINPUT88), .Z(n431) );
  XNOR2_X1 U488 ( .A(KEYINPUT85), .B(KEYINPUT89), .ZN(n430) );
  XNOR2_X1 U489 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n447) );
  XOR2_X1 U491 ( .A(KEYINPUT20), .B(KEYINPUT65), .Z(n435) );
  XNOR2_X1 U492 ( .A(G134GAT), .B(G127GAT), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(n437) );
  XOR2_X1 U494 ( .A(G43GAT), .B(G99GAT), .Z(n436) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n443) );
  XOR2_X1 U496 ( .A(KEYINPUT83), .B(n438), .Z(n441) );
  XNOR2_X1 U497 ( .A(G15GAT), .B(n439), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U499 ( .A(n443), .B(n442), .ZN(n445) );
  NAND2_X1 U500 ( .A1(G227GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U501 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U502 ( .A(n447), .B(n446), .Z(n516) );
  INV_X1 U503 ( .A(n516), .ZN(n487) );
  NAND2_X1 U504 ( .A1(n448), .A2(n487), .ZN(n559) );
  NOR2_X1 U505 ( .A1(n527), .A2(n559), .ZN(n452) );
  XNOR2_X1 U506 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n450) );
  NOR2_X1 U507 ( .A1(n572), .A2(n550), .ZN(n476) );
  INV_X1 U508 ( .A(n482), .ZN(n507) );
  XOR2_X1 U509 ( .A(KEYINPUT27), .B(n507), .Z(n460) );
  NOR2_X1 U510 ( .A1(n459), .A2(n487), .ZN(n453) );
  XNOR2_X1 U511 ( .A(n453), .B(KEYINPUT26), .ZN(n564) );
  AND2_X1 U512 ( .A1(n460), .A2(n564), .ZN(n531) );
  NAND2_X1 U513 ( .A1(n487), .A2(n482), .ZN(n454) );
  NAND2_X1 U514 ( .A1(n459), .A2(n454), .ZN(n455) );
  XNOR2_X1 U515 ( .A(KEYINPUT25), .B(n455), .ZN(n456) );
  NOR2_X1 U516 ( .A1(n531), .A2(n456), .ZN(n457) );
  NOR2_X1 U517 ( .A1(n458), .A2(n457), .ZN(n463) );
  XNOR2_X1 U518 ( .A(KEYINPUT28), .B(n459), .ZN(n512) );
  AND2_X1 U519 ( .A1(n512), .A2(n460), .ZN(n461) );
  NAND2_X1 U520 ( .A1(n461), .A2(n478), .ZN(n515) );
  NOR2_X1 U521 ( .A1(n487), .A2(n515), .ZN(n462) );
  NOR2_X1 U522 ( .A1(n463), .A2(n462), .ZN(n473) );
  NOR2_X1 U523 ( .A1(n546), .A2(n577), .ZN(n464) );
  XOR2_X1 U524 ( .A(KEYINPUT16), .B(n464), .Z(n465) );
  NOR2_X1 U525 ( .A1(n473), .A2(n465), .ZN(n495) );
  NAND2_X1 U526 ( .A1(n476), .A2(n495), .ZN(n471) );
  NOR2_X1 U527 ( .A1(n533), .A2(n471), .ZN(n466) );
  XOR2_X1 U528 ( .A(KEYINPUT34), .B(n466), .Z(n467) );
  XNOR2_X1 U529 ( .A(G1GAT), .B(n467), .ZN(G1324GAT) );
  NOR2_X1 U530 ( .A1(n507), .A2(n471), .ZN(n468) );
  XOR2_X1 U531 ( .A(G8GAT), .B(n468), .Z(G1325GAT) );
  NOR2_X1 U532 ( .A1(n516), .A2(n471), .ZN(n470) );
  XNOR2_X1 U533 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n469) );
  XNOR2_X1 U534 ( .A(n470), .B(n469), .ZN(G1326GAT) );
  NOR2_X1 U535 ( .A1(n512), .A2(n471), .ZN(n472) );
  XOR2_X1 U536 ( .A(G22GAT), .B(n472), .Z(G1327GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT39), .B(KEYINPUT100), .Z(n480) );
  NOR2_X1 U538 ( .A1(n580), .A2(n473), .ZN(n474) );
  NAND2_X1 U539 ( .A1(n577), .A2(n474), .ZN(n475) );
  XNOR2_X1 U540 ( .A(KEYINPUT37), .B(n475), .ZN(n505) );
  NAND2_X1 U541 ( .A1(n476), .A2(n505), .ZN(n477) );
  XOR2_X1 U542 ( .A(KEYINPUT38), .B(n477), .Z(n492) );
  NAND2_X1 U543 ( .A1(n492), .A2(n478), .ZN(n479) );
  XNOR2_X1 U544 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U545 ( .A(G29GAT), .B(n481), .ZN(G1328GAT) );
  XOR2_X1 U546 ( .A(G36GAT), .B(KEYINPUT101), .Z(n484) );
  NAND2_X1 U547 ( .A1(n492), .A2(n482), .ZN(n483) );
  XNOR2_X1 U548 ( .A(n484), .B(n483), .ZN(G1329GAT) );
  XOR2_X1 U549 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n486) );
  XNOR2_X1 U550 ( .A(G43GAT), .B(KEYINPUT103), .ZN(n485) );
  XNOR2_X1 U551 ( .A(n486), .B(n485), .ZN(n490) );
  NAND2_X1 U552 ( .A1(n492), .A2(n487), .ZN(n488) );
  XNOR2_X1 U553 ( .A(n488), .B(KEYINPUT102), .ZN(n489) );
  XNOR2_X1 U554 ( .A(n490), .B(n489), .ZN(G1330GAT) );
  XOR2_X1 U555 ( .A(G50GAT), .B(KEYINPUT105), .Z(n494) );
  INV_X1 U556 ( .A(n512), .ZN(n491) );
  NAND2_X1 U557 ( .A1(n492), .A2(n491), .ZN(n493) );
  XNOR2_X1 U558 ( .A(n494), .B(n493), .ZN(G1331GAT) );
  INV_X1 U559 ( .A(n566), .ZN(n534) );
  NOR2_X1 U560 ( .A1(n534), .A2(n553), .ZN(n504) );
  NAND2_X1 U561 ( .A1(n504), .A2(n495), .ZN(n501) );
  NOR2_X1 U562 ( .A1(n533), .A2(n501), .ZN(n497) );
  XNOR2_X1 U563 ( .A(KEYINPUT42), .B(KEYINPUT106), .ZN(n496) );
  XNOR2_X1 U564 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U565 ( .A(G57GAT), .B(n498), .Z(G1332GAT) );
  NOR2_X1 U566 ( .A1(n507), .A2(n501), .ZN(n499) );
  XOR2_X1 U567 ( .A(G64GAT), .B(n499), .Z(G1333GAT) );
  NOR2_X1 U568 ( .A1(n516), .A2(n501), .ZN(n500) );
  XOR2_X1 U569 ( .A(G71GAT), .B(n500), .Z(G1334GAT) );
  NOR2_X1 U570 ( .A1(n512), .A2(n501), .ZN(n503) );
  XNOR2_X1 U571 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n502) );
  XNOR2_X1 U572 ( .A(n503), .B(n502), .ZN(G1335GAT) );
  NAND2_X1 U573 ( .A1(n505), .A2(n504), .ZN(n511) );
  NOR2_X1 U574 ( .A1(n533), .A2(n511), .ZN(n506) );
  XOR2_X1 U575 ( .A(G85GAT), .B(n506), .Z(G1336GAT) );
  NOR2_X1 U576 ( .A1(n507), .A2(n511), .ZN(n509) );
  XNOR2_X1 U577 ( .A(G92GAT), .B(KEYINPUT107), .ZN(n508) );
  XNOR2_X1 U578 ( .A(n509), .B(n508), .ZN(G1337GAT) );
  NOR2_X1 U579 ( .A1(n516), .A2(n511), .ZN(n510) );
  XOR2_X1 U580 ( .A(G99GAT), .B(n510), .Z(G1338GAT) );
  NOR2_X1 U581 ( .A1(n512), .A2(n511), .ZN(n513) );
  XOR2_X1 U582 ( .A(KEYINPUT44), .B(n513), .Z(n514) );
  XNOR2_X1 U583 ( .A(G106GAT), .B(n514), .ZN(G1339GAT) );
  NOR2_X1 U584 ( .A1(n516), .A2(n515), .ZN(n517) );
  NAND2_X1 U585 ( .A1(n517), .A2(n530), .ZN(n526) );
  NOR2_X1 U586 ( .A1(n550), .A2(n526), .ZN(n518) );
  XOR2_X1 U587 ( .A(G113GAT), .B(n518), .Z(n519) );
  XNOR2_X1 U588 ( .A(KEYINPUT110), .B(n519), .ZN(G1340GAT) );
  NOR2_X1 U589 ( .A1(n553), .A2(n526), .ZN(n521) );
  XNOR2_X1 U590 ( .A(KEYINPUT111), .B(KEYINPUT49), .ZN(n520) );
  XNOR2_X1 U591 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U592 ( .A(G120GAT), .B(n522), .Z(G1341GAT) );
  NOR2_X1 U593 ( .A1(n560), .A2(n526), .ZN(n524) );
  XNOR2_X1 U594 ( .A(KEYINPUT50), .B(KEYINPUT112), .ZN(n523) );
  XNOR2_X1 U595 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U596 ( .A(G127GAT), .B(n525), .Z(G1342GAT) );
  NOR2_X1 U597 ( .A1(n527), .A2(n526), .ZN(n529) );
  XNOR2_X1 U598 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n528) );
  XNOR2_X1 U599 ( .A(n529), .B(n528), .ZN(G1343GAT) );
  NAND2_X1 U600 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U601 ( .A1(n533), .A2(n532), .ZN(n547) );
  NAND2_X1 U602 ( .A1(n534), .A2(n547), .ZN(n535) );
  XNOR2_X1 U603 ( .A(G141GAT), .B(n535), .ZN(G1344GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT115), .B(KEYINPUT114), .Z(n537) );
  XNOR2_X1 U605 ( .A(KEYINPUT52), .B(KEYINPUT53), .ZN(n536) );
  XNOR2_X1 U606 ( .A(n537), .B(n536), .ZN(n542) );
  XOR2_X1 U607 ( .A(G148GAT), .B(KEYINPUT113), .Z(n540) );
  NAND2_X1 U608 ( .A1(n547), .A2(n538), .ZN(n539) );
  XNOR2_X1 U609 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U610 ( .A(n542), .B(n541), .Z(G1345GAT) );
  XNOR2_X1 U611 ( .A(G155GAT), .B(KEYINPUT116), .ZN(n545) );
  NAND2_X1 U612 ( .A1(n547), .A2(n543), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(G1346GAT) );
  XOR2_X1 U614 ( .A(G162GAT), .B(KEYINPUT117), .Z(n549) );
  NAND2_X1 U615 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(G1347GAT) );
  NOR2_X1 U617 ( .A1(n550), .A2(n559), .ZN(n552) );
  XNOR2_X1 U618 ( .A(G169GAT), .B(KEYINPUT119), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(G1348GAT) );
  NOR2_X1 U620 ( .A1(n553), .A2(n559), .ZN(n558) );
  XOR2_X1 U621 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n555) );
  XNOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT120), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U624 ( .A(KEYINPUT56), .B(n556), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(G1349GAT) );
  NOR2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n562) );
  XNOR2_X1 U627 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G183GAT), .B(n563), .ZN(G1350GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n579) );
  NOR2_X1 U631 ( .A1(n566), .A2(n579), .ZN(n571) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n568) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(KEYINPUT59), .B(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n575) );
  INV_X1 U638 ( .A(n579), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XOR2_X1 U641 ( .A(G204GAT), .B(n576), .Z(G1353GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n579), .ZN(n578) );
  XOR2_X1 U643 ( .A(G211GAT), .B(n578), .Z(G1354GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(KEYINPUT62), .B(n581), .Z(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

