//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n440, new_n441, new_n448, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n565,
    new_n567, new_n568, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n628, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1275,
    new_n1276, new_n1277, new_n1278;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  AND2_X1   g014(.A1(KEYINPUT64), .A2(G57), .ZN(new_n440));
  NOR2_X1   g015(.A1(KEYINPUT64), .A2(G57), .ZN(new_n441));
  NOR2_X1   g016(.A1(new_n440), .A2(new_n441), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  INV_X1    g025(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g026(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n451), .A2(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT66), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n457), .A2(G567), .ZN(new_n460));
  AND2_X1   g035(.A1(new_n460), .A2(KEYINPUT67), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(KEYINPUT67), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n455), .A2(G2106), .ZN(new_n463));
  NOR3_X1   g038(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(G319));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n468), .A3(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n471), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT69), .B1(new_n467), .B2(KEYINPUT3), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n479), .A2(new_n465), .A3(G2104), .ZN(new_n480));
  AND4_X1   g055(.A1(new_n477), .A2(new_n478), .A3(new_n480), .A4(new_n468), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n467), .A2(G2105), .ZN(new_n482));
  AOI22_X1  g057(.A1(new_n481), .A2(G137), .B1(G101), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n476), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G160));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n477), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n478), .A2(new_n480), .A3(new_n477), .A4(new_n468), .ZN(new_n488));
  INV_X1    g063(.A(G136), .ZN(new_n489));
  INV_X1    g064(.A(G124), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n478), .A2(new_n480), .A3(G2105), .A4(new_n468), .ZN(new_n491));
  OAI221_X1 g066(.A(new_n487), .B1(new_n488), .B2(new_n489), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n478), .A2(new_n480), .A3(new_n468), .A4(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n466), .A2(new_n468), .ZN(new_n497));
  NOR3_X1   g072(.A1(new_n494), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n496), .A2(KEYINPUT4), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n500), .B(G2104), .C1(G114), .C2(new_n477), .ZN(new_n501));
  INV_X1    g076(.A(G126), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n501), .B1(new_n491), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n499), .A2(new_n503), .ZN(G164));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT70), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G651), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n506), .A2(new_n508), .A3(KEYINPUT6), .ZN(new_n509));
  OR2_X1    g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n509), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G88), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT70), .B(G651), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n512), .A2(G62), .ZN(new_n520));
  AND2_X1   g095(.A1(G75), .A2(G543), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g097(.A(G543), .B1(new_n505), .B2(KEYINPUT6), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n523), .B1(new_n518), .B2(KEYINPUT6), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G50), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n517), .A2(new_n522), .A3(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT72), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT72), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n530), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT7), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n529), .A2(new_n534), .A3(new_n531), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n524), .A2(G51), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT71), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n510), .A2(new_n538), .A3(new_n511), .ZN(new_n539));
  AND2_X1   g114(.A1(KEYINPUT5), .A2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(KEYINPUT5), .A2(G543), .ZN(new_n541));
  OAI21_X1  g116(.A(KEYINPUT71), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n539), .A2(new_n542), .A3(G63), .A4(G651), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n509), .A2(new_n512), .A3(G89), .A4(new_n514), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n536), .A2(new_n537), .A3(new_n543), .A4(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  NAND3_X1  g121(.A1(new_n539), .A2(new_n542), .A3(G64), .ZN(new_n547));
  NAND2_X1  g122(.A1(G77), .A2(G543), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n518), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  XNOR2_X1  g124(.A(KEYINPUT73), .B(G90), .ZN(new_n550));
  NAND4_X1  g125(.A1(new_n509), .A2(new_n512), .A3(new_n514), .A4(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n523), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n509), .A2(new_n552), .A3(G52), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n549), .A2(new_n554), .ZN(G171));
  INV_X1    g130(.A(G81), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n509), .A2(new_n552), .ZN(new_n557));
  INV_X1    g132(.A(G43), .ZN(new_n558));
  OAI22_X1  g133(.A1(new_n515), .A2(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n539), .A2(new_n542), .A3(G56), .ZN(new_n560));
  NAND2_X1  g135(.A1(G68), .A2(G543), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n518), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT74), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  INV_X1    g144(.A(G53), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT9), .B1(new_n557), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n524), .A2(new_n572), .A3(G53), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n540), .A2(new_n541), .ZN(new_n576));
  INV_X1    g151(.A(G65), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G651), .ZN(new_n579));
  INV_X1    g154(.A(G91), .ZN(new_n580));
  AND3_X1   g155(.A1(new_n506), .A2(new_n508), .A3(KEYINPUT6), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n514), .B1(new_n540), .B2(new_n541), .ZN(new_n582));
  OAI21_X1  g157(.A(KEYINPUT75), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT75), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n509), .A2(new_n512), .A3(new_n584), .A4(new_n514), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g161(.A(new_n574), .B(new_n579), .C1(new_n580), .C2(new_n586), .ZN(G299));
  INV_X1    g162(.A(G171), .ZN(G301));
  AND2_X1   g163(.A1(new_n583), .A2(new_n585), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G87), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n539), .A2(new_n542), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n591), .B2(G74), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n524), .A2(G49), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n590), .A2(new_n592), .A3(new_n593), .ZN(G288));
  NAND3_X1  g169(.A1(new_n583), .A2(G86), .A3(new_n585), .ZN(new_n595));
  OAI21_X1  g170(.A(G61), .B1(new_n540), .B2(new_n541), .ZN(new_n596));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(G48), .A2(new_n524), .B1(new_n598), .B2(new_n519), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(G305));
  NAND2_X1  g175(.A1(new_n591), .A2(G60), .ZN(new_n601));
  NAND2_X1  g176(.A1(G72), .A2(G543), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n518), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(G85), .ZN(new_n604));
  INV_X1    g179(.A(G47), .ZN(new_n605));
  OAI22_X1  g180(.A1(new_n515), .A2(new_n604), .B1(new_n557), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(G290));
  NAND2_X1  g183(.A1(G301), .A2(G868), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n583), .A2(G92), .A3(new_n585), .ZN(new_n610));
  XOR2_X1   g185(.A(KEYINPUT76), .B(KEYINPUT10), .Z(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g188(.A1(new_n583), .A2(G92), .A3(new_n585), .A4(new_n611), .ZN(new_n614));
  NAND2_X1  g189(.A1(G79), .A2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G66), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n576), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G651), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n524), .A2(G54), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n613), .A2(new_n614), .A3(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n609), .B1(new_n623), .B2(G868), .ZN(G284));
  OAI21_X1  g199(.A(new_n609), .B1(new_n623), .B2(G868), .ZN(G321));
  MUX2_X1   g200(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g201(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n623), .B1(new_n628), .B2(G860), .ZN(G148));
  OR2_X1    g204(.A1(new_n559), .A2(new_n562), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n623), .A2(new_n628), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT77), .ZN(new_n632));
  MUX2_X1   g207(.A(new_n630), .B(new_n632), .S(G868), .Z(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g209(.A1(new_n477), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT12), .Z(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT13), .ZN(new_n638));
  AOI22_X1  g213(.A1(new_n637), .A2(new_n638), .B1(KEYINPUT78), .B2(G2100), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(new_n638), .B2(new_n637), .ZN(new_n640));
  NOR2_X1   g215(.A1(KEYINPUT78), .A2(G2100), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT79), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(new_n477), .B2(G111), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n644), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n645));
  NOR3_X1   g220(.A1(new_n643), .A2(new_n477), .A3(G111), .ZN(new_n646));
  INV_X1    g221(.A(G123), .ZN(new_n647));
  OAI22_X1  g222(.A1(new_n645), .A2(new_n646), .B1(new_n491), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n648), .B1(G135), .B2(new_n481), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2096), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n642), .A2(new_n650), .ZN(G156));
  INV_X1    g226(.A(KEYINPUT14), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2427), .B(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2430), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n652), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n656), .B1(new_n655), .B2(new_n654), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n657), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2443), .B(G2446), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(G14), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(G401));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2072), .B(G2078), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT80), .ZN(new_n671));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  OR3_X1    g247(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n671), .B1(new_n670), .B2(new_n672), .ZN(new_n674));
  INV_X1    g249(.A(new_n668), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n669), .B(KEYINPUT17), .Z(new_n676));
  OAI211_X1 g251(.A(new_n673), .B(new_n674), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n672), .A2(new_n668), .A3(new_n669), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT18), .Z(new_n679));
  NAND3_X1  g254(.A1(new_n676), .A2(new_n672), .A3(new_n675), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n677), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G2096), .B(G2100), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G227));
  INV_X1    g259(.A(G1986), .ZN(new_n685));
  XOR2_X1   g260(.A(G1971), .B(G1976), .Z(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT81), .B(KEYINPUT19), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT81), .B(KEYINPUT19), .Z(new_n689));
  XNOR2_X1  g264(.A(G1971), .B(G1976), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1956), .B(G2474), .Z(new_n693));
  XOR2_X1   g268(.A(G1961), .B(G1966), .Z(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT83), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n693), .A2(new_n694), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NOR3_X1   g275(.A1(new_n692), .A2(new_n700), .A3(new_n695), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G1981), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n700), .A2(KEYINPUT82), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT82), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n699), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n704), .A2(new_n692), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT20), .ZN(new_n708));
  AND3_X1   g283(.A1(new_n702), .A2(new_n703), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n703), .B1(new_n702), .B2(new_n708), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n685), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n702), .A2(new_n708), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G1981), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n702), .A2(new_n708), .A3(new_n703), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n713), .A2(G1986), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT84), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n711), .A2(new_n715), .A3(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n718), .B1(new_n711), .B2(new_n715), .ZN(new_n721));
  XNOR2_X1  g296(.A(G1991), .B(G1996), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  NOR3_X1   g298(.A1(new_n720), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n711), .A2(new_n715), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(new_n717), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n722), .B1(new_n726), .B2(new_n719), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n724), .A2(new_n727), .ZN(G229));
  INV_X1    g303(.A(G16), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G22), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT87), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G303), .B2(G16), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G1971), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n729), .A2(G23), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(G288), .B2(G16), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT33), .B(G1976), .Z(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n729), .A2(G6), .ZN(new_n740));
  INV_X1    g315(.A(G305), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(new_n729), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT32), .B(G1981), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n735), .A2(new_n737), .ZN(new_n745));
  NOR3_X1   g320(.A1(new_n739), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT34), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT88), .Z(new_n749));
  INV_X1    g324(.A(G29), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G25), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT85), .Z(new_n752));
  AND2_X1   g327(.A1(new_n481), .A2(G131), .ZN(new_n753));
  INV_X1    g328(.A(G119), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n477), .A2(G107), .ZN(new_n755));
  OAI21_X1  g330(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n756));
  OAI22_X1  g331(.A1(new_n491), .A2(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n752), .B1(new_n758), .B2(new_n750), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT35), .B(G1991), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT86), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n759), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n729), .A2(G24), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n607), .B2(new_n729), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G1986), .ZN(new_n765));
  AOI211_X1 g340(.A(new_n762), .B(new_n765), .C1(new_n746), .C2(new_n747), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n749), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(KEYINPUT36), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT36), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n749), .A2(new_n769), .A3(new_n766), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n750), .B1(KEYINPUT24), .B2(G34), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(KEYINPUT24), .B2(G34), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n484), .B2(G29), .ZN(new_n774));
  INV_X1    g349(.A(G2084), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT93), .Z(new_n777));
  INV_X1    g352(.A(G2090), .ZN(new_n778));
  NOR2_X1   g353(.A1(G29), .A2(G35), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G162), .B2(G29), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n777), .B1(new_n778), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(G4), .A2(G16), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n623), .B2(G16), .ZN(new_n785));
  OAI22_X1  g360(.A1(new_n782), .A2(new_n778), .B1(G1348), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G1348), .B2(new_n785), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n729), .A2(G5), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G171), .B2(new_n729), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G1961), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT92), .Z(new_n791));
  NAND2_X1  g366(.A1(G299), .A2(G16), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n729), .A2(G20), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT23), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(G1956), .Z(new_n796));
  NAND4_X1  g371(.A1(new_n783), .A2(new_n787), .A3(new_n791), .A4(new_n796), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n477), .A2(G103), .A3(G2104), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT25), .ZN(new_n799));
  INV_X1    g374(.A(G139), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n488), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n497), .A2(G127), .ZN(new_n802));
  INV_X1    g377(.A(G115), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(new_n467), .ZN(new_n804));
  AOI211_X1 g379(.A(new_n799), .B(new_n801), .C1(new_n804), .C2(G2105), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n805), .A2(new_n750), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n750), .B2(G33), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n808), .A2(G2072), .ZN(new_n809));
  NOR2_X1   g384(.A1(G16), .A2(G19), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n563), .B2(G16), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT89), .B(G1341), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(G27), .A2(G29), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G164), .B2(G29), .ZN(new_n815));
  INV_X1    g390(.A(G2078), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT30), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n819), .A2(G28), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n750), .B1(new_n819), .B2(G28), .ZN(new_n821));
  AND2_X1   g396(.A1(KEYINPUT31), .A2(G11), .ZN(new_n822));
  NOR2_X1   g397(.A1(KEYINPUT31), .A2(G11), .ZN(new_n823));
  OAI22_X1  g398(.A1(new_n820), .A2(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(new_n649), .B2(G29), .ZN(new_n825));
  INV_X1    g400(.A(G2072), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n807), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n750), .A2(G32), .ZN(new_n828));
  NAND3_X1  g403(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT26), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n830), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n831), .A2(new_n832), .B1(G105), .B2(new_n482), .ZN(new_n833));
  INV_X1    g408(.A(G129), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n491), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(G141), .B2(new_n481), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n828), .B1(new_n836), .B2(new_n750), .ZN(new_n837));
  XOR2_X1   g412(.A(KEYINPUT27), .B(G1996), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NOR4_X1   g414(.A1(new_n809), .A2(new_n818), .A3(new_n827), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n750), .A2(G26), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT28), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n481), .A2(G140), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n480), .A2(new_n468), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n844), .A2(G128), .A3(G2105), .A4(new_n478), .ZN(new_n845));
  OR2_X1    g420(.A1(G104), .A2(G2105), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n846), .B(G2104), .C1(G116), .C2(new_n477), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n843), .A2(new_n845), .A3(KEYINPUT90), .A4(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT90), .ZN(new_n849));
  INV_X1    g424(.A(G128), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n847), .B1(new_n491), .B2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(G140), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n488), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n849), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n848), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n842), .B1(new_n856), .B2(new_n750), .ZN(new_n857));
  INV_X1    g432(.A(G2067), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n729), .A2(G21), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(G168), .B2(new_n729), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(G1966), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT91), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n789), .A2(G1961), .ZN(new_n864));
  OAI221_X1 g439(.A(new_n864), .B1(G1966), .B2(new_n861), .C1(new_n775), .C2(new_n774), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n840), .A2(new_n859), .A3(new_n863), .A4(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n797), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n771), .A2(new_n868), .ZN(G150));
  INV_X1    g444(.A(G150), .ZN(G311));
  NAND2_X1  g445(.A1(new_n623), .A2(G559), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT38), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n539), .A2(new_n542), .A3(G67), .ZN(new_n873));
  NAND2_X1  g448(.A1(G80), .A2(G543), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n518), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(KEYINPUT95), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n509), .A2(new_n512), .A3(G93), .A4(new_n514), .ZN(new_n878));
  XOR2_X1   g453(.A(KEYINPUT96), .B(G55), .Z(new_n879));
  NAND3_X1  g454(.A1(new_n879), .A2(new_n509), .A3(new_n552), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(new_n875), .B2(KEYINPUT95), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n630), .B1(new_n877), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT95), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n873), .A2(new_n874), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n884), .B1(new_n885), .B2(new_n518), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n886), .A2(new_n563), .A3(new_n876), .A4(new_n881), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n872), .B(new_n888), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n889), .A2(KEYINPUT39), .ZN(new_n890));
  INV_X1    g465(.A(G860), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(KEYINPUT39), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n877), .A2(new_n882), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n894), .A2(new_n891), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT37), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(new_n896), .ZN(G145));
  INV_X1    g472(.A(KEYINPUT99), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n649), .B(G162), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(G160), .ZN(new_n900));
  INV_X1    g475(.A(new_n836), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n848), .A2(new_n854), .A3(G164), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(G164), .B1(new_n848), .B2(new_n854), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n903), .A2(new_n904), .A3(new_n805), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n799), .B1(new_n804), .B2(G2105), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(new_n800), .B2(new_n488), .ZN(new_n907));
  INV_X1    g482(.A(G164), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n855), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n907), .B1(new_n909), .B2(new_n902), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n901), .B1(new_n905), .B2(new_n910), .ZN(new_n911));
  OR2_X1    g486(.A1(G106), .A2(G2105), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n912), .B(G2104), .C1(G118), .C2(new_n477), .ZN(new_n913));
  INV_X1    g488(.A(G142), .ZN(new_n914));
  INV_X1    g489(.A(G130), .ZN(new_n915));
  OAI221_X1 g490(.A(new_n913), .B1(new_n488), .B2(new_n914), .C1(new_n915), .C2(new_n491), .ZN(new_n916));
  OR2_X1    g491(.A1(new_n916), .A2(new_n636), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n636), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n917), .A2(new_n758), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n758), .B1(new_n917), .B2(new_n918), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n805), .B1(new_n903), .B2(new_n904), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n909), .A2(new_n907), .A3(new_n902), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n923), .A3(new_n836), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n911), .A2(new_n921), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT98), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT98), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n911), .A2(new_n927), .A3(new_n921), .A4(new_n924), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT97), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n911), .A2(new_n924), .ZN(new_n931));
  INV_X1    g506(.A(new_n921), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI211_X1 g508(.A(KEYINPUT97), .B(new_n921), .C1(new_n911), .C2(new_n924), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n900), .B1(new_n929), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n931), .A2(new_n932), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n937), .A2(new_n900), .A3(new_n925), .ZN(new_n938));
  INV_X1    g513(.A(G37), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n898), .B1(new_n936), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n937), .A2(KEYINPUT97), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n931), .A2(new_n930), .A3(new_n932), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n942), .A2(new_n926), .A3(new_n928), .A4(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n900), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n940), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n946), .A2(KEYINPUT99), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n941), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n949), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g525(.A1(new_n883), .A2(new_n887), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n632), .B(new_n951), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n589), .A2(G91), .B1(G651), .B2(new_n578), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n620), .B1(new_n610), .B2(new_n612), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n953), .A2(new_n954), .A3(new_n574), .A4(new_n614), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n622), .A2(G299), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n952), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(KEYINPUT41), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT41), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n955), .A2(new_n956), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT100), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT100), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n964), .B1(new_n957), .B2(KEYINPUT41), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n959), .B1(new_n966), .B2(new_n952), .ZN(new_n967));
  NAND2_X1  g542(.A1(G290), .A2(new_n741), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n607), .A2(G305), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(G288), .A2(G166), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n590), .A2(G303), .A3(new_n592), .A4(new_n593), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OR2_X1    g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  AOI22_X1  g549(.A1(new_n968), .A2(new_n969), .B1(new_n971), .B2(new_n972), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n977), .B(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n967), .B(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(G868), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(G868), .B2(new_n894), .ZN(G295));
  OAI21_X1  g557(.A(new_n981), .B1(G868), .B2(new_n894), .ZN(G331));
  NAND3_X1  g558(.A1(new_n974), .A2(KEYINPUT106), .A3(new_n976), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n970), .A2(new_n973), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n985), .B1(new_n986), .B2(new_n975), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n960), .A2(new_n962), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n551), .A2(new_n553), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT102), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n547), .A2(new_n548), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n991), .B(new_n992), .C1(new_n993), .C2(new_n518), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT102), .B1(new_n549), .B2(new_n554), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n994), .A2(G168), .A3(new_n995), .ZN(new_n996));
  OAI211_X1 g571(.A(G286), .B(KEYINPUT102), .C1(new_n549), .C2(new_n554), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n883), .A2(new_n887), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n998), .B(KEYINPUT105), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n996), .A2(new_n997), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n951), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT104), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT104), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n951), .A2(new_n1000), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n990), .B1(new_n999), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1001), .A2(KEYINPUT103), .A3(new_n998), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1000), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT103), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(new_n888), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT107), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(new_n1012), .A3(new_n958), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1006), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1012), .B1(new_n1011), .B2(new_n958), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n989), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT43), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1010), .B(new_n1007), .C1(new_n963), .C2(new_n965), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1008), .A2(new_n888), .A3(KEYINPUT105), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT105), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n998), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1022), .A2(new_n958), .A3(new_n1002), .A4(new_n1004), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1018), .A2(new_n977), .A3(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1016), .A2(new_n1017), .A3(new_n939), .A4(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n939), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n988), .B1(new_n1018), .B2(new_n1023), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT43), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1017), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1016), .A2(new_n939), .A3(new_n1024), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1030), .B1(new_n1031), .B2(new_n1017), .ZN(new_n1032));
  MUX2_X1   g607(.A(new_n1029), .B(new_n1032), .S(KEYINPUT44), .Z(G397));
  XNOR2_X1  g608(.A(new_n855), .B(new_n858), .ZN(new_n1034));
  INV_X1    g609(.A(G101), .ZN(new_n1035));
  INV_X1    g610(.A(new_n482), .ZN(new_n1036));
  INV_X1    g611(.A(G137), .ZN(new_n1037));
  OAI221_X1 g612(.A(G40), .B1(new_n1035), .B2(new_n1036), .C1(new_n488), .C2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n476), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G1384), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(new_n499), .B2(new_n503), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT45), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1034), .A2(new_n1046), .ZN(new_n1047));
  XOR2_X1   g622(.A(new_n1047), .B(KEYINPUT108), .Z(new_n1048));
  INV_X1    g623(.A(G1996), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n836), .B(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1048), .B1(new_n1045), .B2(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n758), .B(new_n761), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1051), .B1(new_n1046), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(G290), .A2(G1986), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n607), .A2(new_n685), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1046), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  XOR2_X1   g632(.A(G299), .B(KEYINPUT57), .Z(new_n1058));
  OAI211_X1 g633(.A(KEYINPUT45), .B(new_n1041), .C1(new_n499), .C2(new_n503), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1044), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1038), .B1(new_n474), .B2(new_n475), .ZN(new_n1061));
  XNOR2_X1  g636(.A(KEYINPUT56), .B(G2072), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1042), .A2(KEYINPUT50), .ZN(new_n1064));
  NOR2_X1   g639(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1065), .B1(new_n499), .B2(new_n503), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT114), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT114), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1068), .B(new_n1065), .C1(new_n499), .C2(new_n503), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1064), .A2(new_n1067), .A3(new_n1061), .A4(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT117), .B(G1956), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(KEYINPUT118), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT118), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1058), .B(new_n1063), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT119), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n1072), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1080), .A2(new_n1081), .A3(new_n1058), .A4(new_n1063), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1076), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1064), .A2(KEYINPUT109), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT109), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1042), .A2(new_n1085), .A3(KEYINPUT50), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1084), .A2(new_n1061), .A3(new_n1086), .A4(new_n1066), .ZN(new_n1087));
  INV_X1    g662(.A(G1348), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n858), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n622), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1058), .B1(new_n1080), .B2(new_n1063), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1083), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1089), .A2(KEYINPUT60), .A3(new_n1091), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n623), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1089), .A2(KEYINPUT60), .A3(new_n622), .A4(new_n1091), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT60), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n630), .A2(KEYINPUT121), .ZN(new_n1102));
  XOR2_X1   g677(.A(KEYINPUT58), .B(G1341), .Z(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1044), .A2(new_n1061), .A3(new_n1049), .A4(new_n1059), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1106), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1102), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(KEYINPUT59), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1111), .B(new_n1102), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1098), .A2(new_n1101), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1093), .B1(new_n1076), .B2(new_n1082), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1113), .B1(KEYINPUT61), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1063), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1058), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT122), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1075), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT61), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NOR3_X1   g695(.A1(new_n1116), .A2(KEYINPUT122), .A3(new_n1117), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1094), .B1(new_n1115), .B2(new_n1122), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1064), .A2(KEYINPUT109), .B1(new_n908), .B2(new_n1065), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1040), .A2(G2090), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1124), .A2(new_n1086), .A3(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1044), .A2(new_n1061), .A3(new_n1059), .ZN(new_n1127));
  INV_X1    g702(.A(G1971), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT110), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(G303), .A2(G8), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT55), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1126), .A2(KEYINPUT110), .A3(new_n1129), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1132), .A2(G8), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n595), .A2(new_n703), .A3(new_n599), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT111), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n595), .A2(new_n599), .A3(KEYINPUT111), .A4(new_n703), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n516), .A2(G86), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n703), .B1(new_n599), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1142), .A2(KEYINPUT49), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT113), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1144), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1149), .A2(KEYINPUT113), .A3(KEYINPUT49), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT112), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT49), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT112), .B1(new_n1149), .B2(KEYINPUT49), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(G8), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1090), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1151), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1160));
  AND2_X1   g735(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT115), .ZN(new_n1162));
  AOI21_X1  g737(.A(G2090), .B1(new_n1070), .B2(new_n1162), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1064), .A2(new_n1061), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1164), .A2(KEYINPUT115), .A3(new_n1067), .A4(new_n1069), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1161), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1134), .B1(new_n1166), .B2(new_n1158), .ZN(new_n1167));
  INV_X1    g742(.A(G288), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(G1976), .ZN(new_n1169));
  INV_X1    g744(.A(G1976), .ZN(new_n1170));
  AOI21_X1  g745(.A(KEYINPUT52), .B1(G288), .B2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1169), .A2(new_n1159), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1061), .A2(new_n1041), .A3(new_n908), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n1173), .B(G8), .C1(G288), .C2(new_n1170), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(KEYINPUT52), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1176), .ZN(new_n1177));
  AND4_X1   g752(.A1(new_n1137), .A2(new_n1160), .A3(new_n1167), .A4(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(G1961), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1087), .A2(new_n1179), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1044), .A2(new_n1061), .A3(new_n816), .A4(new_n1059), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT53), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1060), .A2(KEYINPUT53), .A3(new_n816), .A4(new_n1061), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1180), .A2(G301), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(KEYINPUT54), .ZN(new_n1186));
  AOI22_X1  g761(.A1(new_n1087), .A2(new_n1179), .B1(new_n1182), .B2(new_n1181), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1182), .A2(G2078), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1060), .A2(new_n472), .A3(new_n1039), .A4(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(G301), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(KEYINPUT123), .B1(new_n1186), .B2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1180), .A2(new_n1183), .A3(new_n1189), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1192), .A2(G171), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT123), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1193), .A2(new_n1194), .A3(KEYINPUT54), .A4(new_n1185), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1191), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(G1966), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1127), .A2(new_n1197), .ZN(new_n1198));
  OAI211_X1 g773(.A(G168), .B(new_n1198), .C1(new_n1087), .C2(G2084), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(G8), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1124), .A2(new_n775), .A3(new_n1061), .A4(new_n1086), .ZN(new_n1201));
  AOI21_X1  g776(.A(G168), .B1(new_n1201), .B2(new_n1198), .ZN(new_n1202));
  OAI21_X1  g777(.A(KEYINPUT51), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT51), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1199), .A2(new_n1204), .A3(G8), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1187), .A2(new_n1184), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1207), .A2(G171), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1187), .A2(G301), .A3(new_n1189), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT54), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND4_X1  g787(.A1(new_n1178), .A2(new_n1196), .A3(new_n1206), .A4(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1213), .A2(KEYINPUT124), .ZN(new_n1214));
  INV_X1    g789(.A(new_n1159), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1215), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1176), .B1(new_n1216), .B2(new_n1151), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n1217), .A2(new_n1137), .A3(new_n1167), .ZN(new_n1218));
  AOI21_X1  g793(.A(KEYINPUT54), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1219));
  NOR2_X1   g794(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g795(.A(KEYINPUT124), .ZN(new_n1221));
  NAND4_X1  g796(.A1(new_n1220), .A2(new_n1221), .A3(new_n1196), .A4(new_n1206), .ZN(new_n1222));
  AND3_X1   g797(.A1(new_n1123), .A2(new_n1214), .A3(new_n1222), .ZN(new_n1223));
  NAND3_X1  g798(.A1(new_n1132), .A2(G8), .A3(new_n1136), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1224), .A2(new_n1134), .ZN(new_n1225));
  AOI211_X1 g800(.A(new_n1158), .B(G286), .C1(new_n1201), .C2(new_n1198), .ZN(new_n1226));
  AND2_X1   g801(.A1(new_n1226), .A2(KEYINPUT63), .ZN(new_n1227));
  NAND4_X1  g802(.A1(new_n1225), .A2(new_n1227), .A3(new_n1137), .A4(new_n1217), .ZN(new_n1228));
  NAND4_X1  g803(.A1(new_n1217), .A2(new_n1137), .A3(new_n1167), .A4(new_n1226), .ZN(new_n1229));
  AND2_X1   g804(.A1(new_n1229), .A2(KEYINPUT116), .ZN(new_n1230));
  INV_X1    g805(.A(KEYINPUT63), .ZN(new_n1231));
  OAI21_X1  g806(.A(new_n1231), .B1(new_n1229), .B2(KEYINPUT116), .ZN(new_n1232));
  OAI21_X1  g807(.A(new_n1228), .B1(new_n1230), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g808(.A(KEYINPUT62), .ZN(new_n1234));
  AND3_X1   g809(.A1(new_n1203), .A2(new_n1234), .A3(new_n1205), .ZN(new_n1235));
  AOI21_X1  g810(.A(G301), .B1(new_n1187), .B2(new_n1184), .ZN(new_n1236));
  NAND4_X1  g811(.A1(new_n1217), .A2(new_n1137), .A3(new_n1167), .A4(new_n1236), .ZN(new_n1237));
  OAI21_X1  g812(.A(KEYINPUT125), .B1(new_n1235), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g813(.A(KEYINPUT125), .ZN(new_n1239));
  NAND3_X1  g814(.A1(new_n1203), .A2(new_n1234), .A3(new_n1205), .ZN(new_n1240));
  NAND4_X1  g815(.A1(new_n1178), .A2(new_n1239), .A3(new_n1236), .A4(new_n1240), .ZN(new_n1241));
  NAND2_X1  g816(.A1(new_n1206), .A2(KEYINPUT62), .ZN(new_n1242));
  NAND3_X1  g817(.A1(new_n1238), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  NAND3_X1  g818(.A1(new_n1160), .A2(new_n1170), .A3(new_n1168), .ZN(new_n1244));
  AOI21_X1  g819(.A(new_n1215), .B1(new_n1244), .B2(new_n1142), .ZN(new_n1245));
  INV_X1    g820(.A(new_n1137), .ZN(new_n1246));
  AOI21_X1  g821(.A(new_n1245), .B1(new_n1246), .B2(new_n1217), .ZN(new_n1247));
  NAND3_X1  g822(.A1(new_n1233), .A2(new_n1243), .A3(new_n1247), .ZN(new_n1248));
  OAI21_X1  g823(.A(new_n1057), .B1(new_n1223), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g824(.A1(new_n1045), .A2(new_n1049), .ZN(new_n1250));
  XOR2_X1   g825(.A(new_n1250), .B(KEYINPUT46), .Z(new_n1251));
  AOI21_X1  g826(.A(new_n1046), .B1(new_n1034), .B2(new_n836), .ZN(new_n1252));
  NOR2_X1   g827(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  XOR2_X1   g828(.A(new_n1253), .B(KEYINPUT47), .Z(new_n1254));
  NOR2_X1   g829(.A1(new_n1046), .A2(new_n1055), .ZN(new_n1255));
  XNOR2_X1  g830(.A(new_n1255), .B(KEYINPUT48), .ZN(new_n1256));
  OAI21_X1  g831(.A(new_n1254), .B1(new_n1053), .B2(new_n1256), .ZN(new_n1257));
  NOR3_X1   g832(.A1(new_n753), .A2(new_n761), .A3(new_n757), .ZN(new_n1258));
  NAND2_X1  g833(.A1(new_n1051), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g834(.A1(new_n856), .A2(new_n858), .ZN(new_n1260));
  AOI21_X1  g835(.A(new_n1046), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NOR2_X1   g836(.A1(new_n1257), .A2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g837(.A1(new_n1249), .A2(new_n1262), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g838(.A1(new_n683), .A2(G319), .ZN(new_n1265));
  OAI22_X1  g839(.A1(new_n1265), .A2(KEYINPUT126), .B1(new_n665), .B2(new_n666), .ZN(new_n1266));
  AND2_X1   g840(.A1(new_n1265), .A2(KEYINPUT126), .ZN(new_n1267));
  NOR2_X1   g841(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g842(.A(new_n1268), .B1(new_n724), .B2(new_n727), .ZN(new_n1269));
  INV_X1    g843(.A(new_n1269), .ZN(new_n1270));
  AND4_X1   g844(.A1(KEYINPUT127), .A2(new_n949), .A3(new_n1029), .A4(new_n1270), .ZN(new_n1271));
  AOI21_X1  g845(.A(new_n1269), .B1(new_n941), .B2(new_n948), .ZN(new_n1272));
  AOI21_X1  g846(.A(KEYINPUT127), .B1(new_n1272), .B2(new_n1029), .ZN(new_n1273));
  NOR2_X1   g847(.A1(new_n1271), .A2(new_n1273), .ZN(G308));
  NAND2_X1  g848(.A1(new_n1272), .A2(new_n1029), .ZN(new_n1275));
  INV_X1    g849(.A(KEYINPUT127), .ZN(new_n1276));
  NAND2_X1  g850(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g851(.A1(new_n1272), .A2(KEYINPUT127), .A3(new_n1029), .ZN(new_n1278));
  NAND2_X1  g852(.A1(new_n1277), .A2(new_n1278), .ZN(G225));
endmodule


