//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n748, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G146), .ZN(new_n192));
  NOR3_X1   g006(.A1(new_n188), .A2(KEYINPUT64), .A3(G143), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n189), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  AND2_X1   g008(.A1(KEYINPUT0), .A2(G128), .ZN(new_n195));
  NOR2_X1   g009(.A1(KEYINPUT0), .A2(G128), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(G143), .B(G146), .ZN(new_n198));
  AOI22_X1  g012(.A1(new_n194), .A2(new_n197), .B1(new_n198), .B2(new_n195), .ZN(new_n199));
  INV_X1    g013(.A(G137), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(KEYINPUT11), .A3(G134), .ZN(new_n201));
  INV_X1    g015(.A(G134), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G137), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n200), .A2(G134), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT11), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n207), .B1(new_n202), .B2(G137), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT65), .ZN(new_n210));
  AOI211_X1 g024(.A(G131), .B(new_n204), .C1(new_n208), .C2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n208), .ZN(new_n213));
  INV_X1    g027(.A(new_n204), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n199), .B1(new_n211), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT67), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT2), .ZN(new_n218));
  INV_X1    g032(.A(G113), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT67), .B1(KEYINPUT2), .B2(G113), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(KEYINPUT2), .A2(G113), .ZN(new_n223));
  XNOR2_X1  g037(.A(G116), .B(G119), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n224), .B1(new_n222), .B2(new_n223), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n191), .A2(G146), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT1), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n189), .A2(new_n228), .A3(new_n229), .A4(G128), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT66), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n191), .A2(G146), .ZN(new_n233));
  OAI21_X1  g047(.A(G128), .B1(new_n233), .B2(new_n229), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n194), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT64), .B1(new_n188), .B2(G143), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n190), .A2(new_n191), .A3(G146), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n233), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G128), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n239), .B1(new_n189), .B2(KEYINPUT1), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT66), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n231), .B1(new_n235), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n213), .A2(new_n212), .A3(new_n214), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n203), .A2(new_n205), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G131), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n216), .B(new_n227), .C1(new_n242), .C2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n232), .B1(new_n194), .B2(new_n234), .ZN(new_n250));
  NOR3_X1   g064(.A1(new_n238), .A2(KEYINPUT66), .A3(new_n240), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n230), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(new_n245), .A3(new_n243), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n253), .A2(KEYINPUT68), .A3(new_n227), .A4(new_n216), .ZN(new_n254));
  NOR2_X1   g068(.A1(G237), .A2(G953), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G210), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n256), .B(KEYINPUT27), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(G101), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n257), .B(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n249), .A2(new_n254), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT31), .ZN(new_n263));
  INV_X1    g077(.A(new_n227), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT30), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n265), .B1(new_n253), .B2(new_n216), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n242), .A2(new_n246), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n198), .A2(new_n195), .ZN(new_n268));
  INV_X1    g082(.A(new_n197), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n268), .B1(new_n238), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n213), .A2(new_n214), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G131), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n270), .B1(new_n272), .B2(new_n243), .ZN(new_n273));
  NOR3_X1   g087(.A1(new_n267), .A2(new_n273), .A3(KEYINPUT30), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n264), .B1(new_n266), .B2(new_n274), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n249), .A2(new_n254), .A3(KEYINPUT69), .A4(new_n259), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n262), .A2(new_n263), .A3(new_n275), .A4(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT28), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n247), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n264), .B1(new_n267), .B2(new_n273), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n249), .A2(new_n254), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n280), .B1(new_n282), .B2(KEYINPUT28), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n277), .B1(new_n259), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n276), .A2(new_n275), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n263), .B1(new_n286), .B2(new_n262), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n187), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT32), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n260), .A2(new_n261), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT31), .B1(new_n291), .B2(new_n285), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n282), .A2(KEYINPUT28), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n279), .ZN(new_n294));
  INV_X1    g108(.A(new_n259), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n292), .A2(new_n296), .A3(new_n277), .ZN(new_n297));
  INV_X1    g111(.A(new_n187), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n298), .A2(new_n289), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n253), .A2(new_n265), .A3(new_n216), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT30), .B1(new_n267), .B2(new_n273), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n227), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n249), .A2(new_n254), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n295), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT70), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n293), .A2(new_n259), .A3(new_n279), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT70), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n309), .B(new_n295), .C1(new_n303), .C2(new_n304), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n306), .A2(new_n307), .A3(new_n308), .A4(new_n310), .ZN(new_n311));
  XOR2_X1   g125(.A(KEYINPUT71), .B(G902), .Z(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  AOI211_X1 g127(.A(new_n295), .B(new_n280), .C1(new_n282), .C2(KEYINPUT28), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n313), .B1(new_n314), .B2(KEYINPUT29), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G472), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n290), .A2(new_n300), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n239), .A2(G119), .ZN(new_n319));
  INV_X1    g133(.A(G119), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G128), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT23), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n323), .A2(KEYINPUT23), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n324), .B1(new_n327), .B2(new_n319), .ZN(new_n328));
  XOR2_X1   g142(.A(KEYINPUT74), .B(G110), .Z(new_n329));
  NAND3_X1  g143(.A1(new_n326), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT24), .B(G110), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n322), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n334), .B1(new_n322), .B2(new_n333), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n326), .A2(KEYINPUT75), .A3(new_n328), .A4(new_n329), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n332), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G140), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G125), .ZN(new_n341));
  INV_X1    g155(.A(G125), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G140), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n343), .A3(KEYINPUT16), .ZN(new_n344));
  OR3_X1    g158(.A1(new_n342), .A2(KEYINPUT16), .A3(G140), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT73), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n341), .A2(new_n343), .A3(KEYINPUT73), .A4(KEYINPUT16), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n188), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n341), .A2(new_n343), .A3(KEYINPUT77), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT77), .B1(new_n341), .B2(new_n343), .ZN(new_n351));
  NOR3_X1   g165(.A1(new_n350), .A2(new_n351), .A3(G146), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n339), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n322), .A2(new_n333), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n326), .A2(new_n328), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n355), .B1(new_n356), .B2(G110), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n341), .A2(new_n343), .A3(KEYINPUT16), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n346), .B1(new_n341), .B2(KEYINPUT16), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n188), .B(new_n348), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n357), .B1(new_n361), .B2(new_n349), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n354), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G953), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n364), .A2(G221), .A3(G234), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n365), .B(KEYINPUT78), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT22), .B(G137), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n366), .B(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n363), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n354), .A2(new_n362), .A3(new_n368), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  XOR2_X1   g186(.A(new_n372), .B(KEYINPUT80), .Z(new_n373));
  INV_X1    g187(.A(G217), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n374), .B1(new_n312), .B2(G234), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(G902), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(KEYINPUT25), .B1(new_n372), .B2(new_n312), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n354), .A2(new_n362), .A3(new_n368), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n368), .B1(new_n354), .B2(new_n362), .ZN(new_n380));
  OAI211_X1 g194(.A(KEYINPUT25), .B(new_n312), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n375), .B1(new_n378), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT79), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT79), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n385), .B(new_n375), .C1(new_n378), .C2(new_n382), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n377), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT97), .ZN(new_n389));
  INV_X1    g203(.A(G116), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G122), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(KEYINPUT14), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n390), .A2(G122), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n391), .B1(new_n393), .B2(KEYINPUT14), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n392), .B1(new_n394), .B2(KEYINPUT96), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n395), .B1(KEYINPUT96), .B2(new_n394), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G107), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n191), .A2(G128), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n239), .A2(G143), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G134), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n398), .A2(new_n399), .A3(new_n202), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G122), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G116), .ZN(new_n405));
  INV_X1    g219(.A(G107), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n391), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n397), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n407), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n406), .B1(new_n405), .B2(new_n391), .ZN(new_n412));
  OR2_X1    g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n413), .A2(new_n402), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT13), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n398), .A2(KEYINPUT95), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(KEYINPUT13), .B1(new_n191), .B2(G128), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n418), .A2(KEYINPUT95), .ZN(new_n419));
  OAI221_X1 g233(.A(new_n399), .B1(new_n415), .B2(new_n398), .C1(new_n417), .C2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(G134), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n414), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT9), .B(G234), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n423), .A2(new_n374), .A3(G953), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n410), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n424), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n408), .B1(new_n396), .B2(G107), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n402), .B1(new_n411), .B2(new_n412), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n428), .B1(new_n420), .B2(G134), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n426), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n389), .B1(new_n431), .B2(new_n312), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(G478), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(KEYINPUT15), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n431), .A2(new_n389), .A3(new_n312), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n433), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n431), .A2(new_n312), .ZN(new_n438));
  OR2_X1    g252(.A1(new_n438), .A2(new_n435), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT93), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n442), .B1(new_n361), .B2(new_n349), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n348), .B1(new_n358), .B2(new_n359), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G146), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(KEYINPUT93), .A3(new_n360), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n255), .A2(G214), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT91), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(G143), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n255), .B(G214), .C1(new_n448), .C2(G143), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT92), .B1(new_n452), .B2(G131), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(G131), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT17), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT92), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n450), .A2(new_n451), .A3(new_n456), .A4(new_n212), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n453), .A2(new_n454), .A3(new_n455), .A4(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n452), .A2(KEYINPUT17), .A3(G131), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n443), .A2(new_n446), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(G113), .B(G122), .ZN(new_n461));
  INV_X1    g275(.A(G104), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n461), .B(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(KEYINPUT18), .A2(G131), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n452), .B(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n188), .B1(new_n341), .B2(new_n343), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n465), .B1(new_n352), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n460), .A2(new_n463), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT94), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n460), .A2(KEYINPUT94), .A3(new_n463), .A4(new_n467), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n453), .A2(new_n454), .A3(new_n457), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n350), .A2(new_n351), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n341), .A2(new_n343), .ZN(new_n475));
  MUX2_X1   g289(.A(new_n474), .B(new_n475), .S(KEYINPUT19), .Z(new_n476));
  OAI211_X1 g290(.A(new_n445), .B(new_n473), .C1(new_n476), .C2(G146), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n467), .ZN(new_n478));
  INV_X1    g292(.A(new_n463), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n472), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT20), .ZN(new_n482));
  NOR2_X1   g296(.A1(G475), .A2(G902), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n470), .A2(new_n471), .B1(new_n479), .B2(new_n478), .ZN(new_n485));
  INV_X1    g299(.A(new_n483), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT20), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n460), .A2(new_n467), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n470), .A2(new_n471), .B1(new_n479), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(G475), .B1(new_n490), .B2(G902), .ZN(new_n491));
  NAND2_X1  g305(.A1(G234), .A2(G237), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n492), .A2(G952), .A3(new_n364), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n313), .A2(G953), .A3(new_n492), .ZN(new_n494));
  XOR2_X1   g308(.A(new_n494), .B(KEYINPUT98), .Z(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT21), .B(G898), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(KEYINPUT99), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n493), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n441), .A2(new_n488), .A3(new_n491), .A4(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(G214), .B1(G237), .B2(G902), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(G110), .B(G122), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(KEYINPUT8), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n320), .A2(G116), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n390), .A2(G119), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n508), .A3(KEYINPUT5), .ZN(new_n509));
  OR3_X1    g323(.A1(new_n390), .A2(KEYINPUT5), .A3(G119), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n510), .A3(G113), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT82), .B(G101), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT3), .B1(new_n462), .B2(G107), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT3), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(new_n406), .A3(G104), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n462), .A2(G107), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n512), .A2(new_n513), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n462), .A2(G107), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n406), .A2(G104), .ZN(new_n519));
  OAI21_X1  g333(.A(G101), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AND4_X1   g334(.A1(new_n506), .A2(new_n511), .A3(new_n517), .A4(new_n520), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n506), .A2(new_n511), .B1(new_n517), .B2(new_n520), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n505), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT89), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n506), .A2(new_n511), .A3(new_n517), .A4(new_n520), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n513), .A2(new_n515), .A3(new_n516), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT4), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(new_n528), .A3(G101), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n529), .B1(new_n225), .B2(new_n226), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n527), .A2(G101), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n531), .A2(KEYINPUT4), .A3(new_n517), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n504), .B(new_n526), .C1(new_n530), .C2(new_n532), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n342), .B(new_n230), .C1(new_n250), .C2(new_n251), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n270), .A2(G125), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT87), .ZN(new_n536));
  INV_X1    g350(.A(G224), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n536), .B1(new_n537), .B2(G953), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n364), .A2(KEYINPUT87), .A3(G224), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(KEYINPUT7), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n534), .A2(new_n535), .A3(new_n541), .ZN(new_n542));
  OAI211_X1 g356(.A(KEYINPUT89), .B(new_n505), .C1(new_n521), .C2(new_n522), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n525), .A2(new_n533), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n199), .A2(new_n342), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n342), .B2(new_n242), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT90), .B1(new_n547), .B2(new_n541), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n534), .A2(new_n535), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT90), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(new_n550), .A3(new_n540), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(G902), .B1(new_n545), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n538), .A2(new_n539), .ZN(new_n554));
  XOR2_X1   g368(.A(new_n554), .B(KEYINPUT86), .Z(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  AOI211_X1 g370(.A(G125), .B(new_n231), .C1(new_n235), .C2(new_n241), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n556), .B1(new_n557), .B2(new_n546), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n534), .A2(new_n535), .A3(new_n555), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n526), .B1(new_n530), .B2(new_n532), .ZN(new_n561));
  INV_X1    g375(.A(new_n504), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(KEYINPUT6), .A3(new_n533), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT6), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n561), .A2(new_n565), .A3(new_n562), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n560), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT88), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n560), .A2(new_n564), .A3(KEYINPUT88), .A4(new_n566), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n553), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(G210), .B1(G237), .B2(G902), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n553), .A2(new_n569), .A3(new_n572), .A4(new_n570), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n503), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(G221), .B1(new_n423), .B2(G902), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n364), .A2(G227), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(KEYINPUT81), .ZN(new_n579));
  XNOR2_X1  g393(.A(G110), .B(G140), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n579), .B(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n211), .A2(new_n215), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n517), .A2(new_n520), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n252), .A2(KEYINPUT10), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n189), .A2(new_n228), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n234), .A2(KEYINPUT84), .A3(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT84), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n587), .B1(new_n240), .B2(new_n198), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n230), .A2(KEYINPUT83), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT83), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n198), .A2(new_n590), .A3(new_n229), .A4(G128), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n586), .A2(new_n588), .A3(new_n589), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n583), .ZN(new_n593));
  XOR2_X1   g407(.A(KEYINPUT85), .B(KEYINPUT10), .Z(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n529), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(new_n270), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n531), .A2(KEYINPUT4), .A3(new_n517), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AND4_X1   g413(.A1(new_n582), .A2(new_n584), .A3(new_n595), .A4(new_n599), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n593), .A2(new_n594), .B1(new_n598), .B2(new_n597), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n582), .B1(new_n601), .B2(new_n584), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n581), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n581), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n584), .A2(new_n595), .A3(new_n582), .A4(new_n599), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT12), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n517), .A2(new_n520), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n230), .B(new_n607), .C1(new_n250), .C2(new_n251), .ZN(new_n608));
  AOI211_X1 g422(.A(new_n606), .B(new_n582), .C1(new_n593), .C2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n593), .ZN(new_n610));
  INV_X1    g424(.A(new_n582), .ZN(new_n611));
  AOI21_X1  g425(.A(KEYINPUT12), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n604), .B(new_n605), .C1(new_n609), .C2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n603), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(G469), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n614), .A2(new_n615), .A3(new_n312), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n605), .B1(new_n609), .B2(new_n612), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n581), .ZN(new_n618));
  INV_X1    g432(.A(new_n602), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n619), .A2(new_n604), .A3(new_n605), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n618), .A2(new_n620), .A3(G469), .ZN(new_n621));
  INV_X1    g435(.A(G902), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n616), .A2(new_n621), .A3(new_n624), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n576), .A2(new_n577), .A3(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n318), .A2(new_n388), .A3(new_n501), .A4(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(new_n627), .B(new_n512), .Z(G3));
  AOI21_X1  g442(.A(new_n482), .B1(new_n481), .B2(new_n483), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n485), .A2(KEYINPUT20), .A3(new_n486), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n491), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI211_X1 g445(.A(KEYINPUT97), .B(new_n313), .C1(new_n425), .C2(new_n430), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n432), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT101), .B(G478), .Z(new_n634));
  INV_X1    g448(.A(KEYINPUT33), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n430), .B2(KEYINPUT100), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n431), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n425), .B(new_n430), .C1(KEYINPUT100), .C2(new_n635), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n313), .A2(new_n434), .ZN(new_n640));
  AOI22_X1  g454(.A1(new_n633), .A2(new_n634), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n631), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n550), .B1(new_n549), .B2(new_n540), .ZN(new_n644));
  AOI211_X1 g458(.A(KEYINPUT90), .B(new_n541), .C1(new_n534), .C2(new_n535), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n622), .B1(new_n646), .B2(new_n544), .ZN(new_n647));
  AND4_X1   g461(.A1(KEYINPUT88), .A2(new_n560), .A3(new_n564), .A4(new_n566), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n572), .B1(new_n649), .B2(new_n569), .ZN(new_n650));
  INV_X1    g464(.A(new_n575), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n499), .B(new_n502), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n643), .A2(new_n652), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n625), .A2(new_n577), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n297), .A2(new_n312), .ZN(new_n655));
  AOI22_X1  g469(.A1(new_n655), .A2(G472), .B1(new_n187), .B2(new_n297), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n653), .A2(new_n388), .A3(new_n654), .A4(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT34), .B(G104), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G6));
  INV_X1    g473(.A(G472), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(new_n297), .B2(new_n312), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n259), .B1(new_n293), .B2(new_n279), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n291), .A2(new_n285), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n662), .B1(new_n663), .B2(new_n263), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n298), .B1(new_n664), .B2(new_n292), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n661), .A2(new_n665), .A3(new_n387), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n489), .A2(new_n479), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n472), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n622), .ZN(new_n669));
  AOI21_X1  g483(.A(KEYINPUT102), .B1(new_n669), .B2(G475), .ZN(new_n670));
  OAI211_X1 g484(.A(KEYINPUT102), .B(G475), .C1(new_n490), .C2(G902), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n488), .B(new_n440), .C1(new_n670), .C2(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n652), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n666), .A2(new_n654), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G107), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT103), .B(KEYINPUT35), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G9));
  NOR2_X1   g492(.A1(new_n368), .A2(KEYINPUT36), .ZN(new_n679));
  XOR2_X1   g493(.A(new_n679), .B(KEYINPUT104), .Z(new_n680));
  AND2_X1   g494(.A1(new_n680), .A2(new_n363), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(new_n363), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n376), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n384), .A2(new_n386), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT105), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n384), .A2(new_n686), .A3(new_n386), .A4(new_n683), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n688), .A2(new_n501), .A3(new_n626), .A4(new_n656), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT37), .B(G110), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G12));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n688), .A2(new_n318), .A3(new_n626), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT102), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n491), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n671), .ZN(new_n696));
  INV_X1    g510(.A(G900), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n495), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n493), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n696), .A2(new_n488), .A3(new_n440), .A4(new_n700), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n692), .B1(new_n693), .B2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n300), .ZN(new_n703));
  AOI21_X1  g517(.A(KEYINPUT32), .B1(new_n297), .B2(new_n187), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n660), .B1(new_n311), .B2(new_n315), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n685), .A2(new_n576), .A3(new_n654), .A4(new_n687), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n701), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n708), .A2(KEYINPUT106), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n702), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G128), .ZN(G30));
  XOR2_X1   g526(.A(new_n699), .B(KEYINPUT39), .Z(new_n713));
  NAND2_X1  g527(.A1(new_n654), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(new_n714), .B(KEYINPUT40), .Z(new_n715));
  AND2_X1   g529(.A1(new_n282), .A2(new_n295), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n622), .B1(new_n663), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n703), .B1(new_n717), .B2(G472), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n290), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n631), .A2(new_n440), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(new_n503), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n574), .A2(new_n575), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT107), .B(KEYINPUT38), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(new_n684), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n715), .A2(new_n719), .A3(new_n721), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G143), .ZN(G45));
  AOI211_X1 g541(.A(new_n699), .B(new_n641), .C1(new_n488), .C2(new_n491), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n708), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G146), .ZN(G48));
  AOI21_X1  g544(.A(new_n615), .B1(new_n614), .B2(new_n312), .ZN(new_n731));
  AOI211_X1 g545(.A(G469), .B(new_n313), .C1(new_n603), .C2(new_n613), .ZN(new_n732));
  INV_X1    g546(.A(new_n577), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n318), .A2(new_n653), .A3(new_n388), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT41), .B(G113), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(KEYINPUT108), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n735), .B(new_n737), .ZN(G15));
  NAND4_X1  g552(.A1(new_n318), .A2(new_n674), .A3(new_n388), .A4(new_n734), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G116), .ZN(G18));
  AND2_X1   g554(.A1(new_n576), .A2(new_n734), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n688), .A2(new_n318), .A3(new_n501), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G119), .ZN(G21));
  INV_X1    g557(.A(new_n720), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n576), .A2(new_n734), .A3(new_n499), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n666), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G122), .ZN(G24));
  AND4_X1   g561(.A1(new_n656), .A2(new_n741), .A3(new_n684), .A4(new_n728), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(new_n342), .ZN(G27));
  NOR2_X1   g563(.A1(new_n722), .A2(new_n503), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n641), .B1(new_n488), .B2(new_n491), .ZN(new_n751));
  AND4_X1   g565(.A1(new_n654), .A2(new_n750), .A3(new_n751), .A4(new_n700), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n752), .A2(KEYINPUT42), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT111), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n300), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n297), .A2(KEYINPUT111), .A3(new_n299), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n755), .A2(new_n290), .A3(new_n317), .A4(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n757), .A2(new_n758), .A3(new_n388), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n758), .B1(new_n757), .B2(new_n388), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n753), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT109), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n317), .A2(new_n300), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n388), .B1(new_n763), .B2(new_n704), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n625), .A2(new_n577), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n765), .A2(new_n503), .A3(new_n722), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n728), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n762), .B1(new_n764), .B2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n752), .A2(KEYINPUT109), .A3(new_n318), .A4(new_n388), .ZN(new_n769));
  XOR2_X1   g583(.A(KEYINPUT110), .B(KEYINPUT42), .Z(new_n770));
  NAND3_X1  g584(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n761), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G131), .ZN(G33));
  NAND3_X1  g587(.A1(new_n318), .A2(new_n388), .A3(new_n766), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n701), .B(KEYINPUT113), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  INV_X1    g592(.A(new_n631), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n642), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT43), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n782), .B(new_n684), .C1(new_n665), .C2(new_n661), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT44), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(new_n750), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n618), .A2(new_n620), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n790), .A2(KEYINPUT45), .ZN(new_n791));
  OAI21_X1  g605(.A(G469), .B1(new_n790), .B2(KEYINPUT45), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n623), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT46), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n616), .B1(new_n794), .B2(KEYINPUT46), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n798), .A2(new_n577), .A3(new_n713), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n799), .B1(new_n787), .B2(new_n788), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n789), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(new_n200), .ZN(G39));
  OAI21_X1  g616(.A(new_n577), .B1(new_n796), .B2(new_n797), .ZN(new_n803));
  XOR2_X1   g617(.A(new_n803), .B(KEYINPUT47), .Z(new_n804));
  AND4_X1   g618(.A1(new_n706), .A2(new_n387), .A3(new_n728), .A4(new_n750), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G140), .ZN(G42));
  NOR2_X1   g621(.A1(new_n731), .A2(new_n732), .ZN(new_n808));
  XOR2_X1   g622(.A(new_n808), .B(KEYINPUT49), .Z(new_n809));
  NOR4_X1   g623(.A1(new_n809), .A2(new_n387), .A3(new_n503), .A4(new_n733), .ZN(new_n810));
  INV_X1    g624(.A(new_n719), .ZN(new_n811));
  INV_X1    g625(.A(new_n780), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n810), .A2(new_n811), .A3(new_n724), .A4(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n689), .A2(new_n742), .A3(new_n627), .A4(new_n746), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n440), .B(new_n491), .C1(new_n629), .C2(new_n630), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n816), .A2(KEYINPUT115), .A3(new_n499), .A4(new_n576), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n818), .B1(new_n652), .B2(new_n815), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n666), .A2(new_n817), .A3(new_n819), .A4(new_n654), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n820), .A2(new_n739), .A3(new_n735), .A4(new_n657), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n814), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n656), .A2(new_n684), .A3(new_n728), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n696), .A2(new_n488), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n440), .A2(new_n699), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n824), .A2(new_n685), .A3(new_n687), .A4(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n823), .B1(new_n826), .B2(new_n706), .ZN(new_n827));
  AOI22_X1  g641(.A1(new_n766), .A2(new_n827), .B1(new_n775), .B2(new_n776), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n772), .A2(new_n822), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(KEYINPUT116), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n748), .B1(new_n708), .B2(new_n728), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n684), .A2(new_n699), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT117), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n721), .A2(new_n722), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n833), .A2(new_n719), .A3(new_n834), .A4(new_n654), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT106), .B1(new_n708), .B2(new_n709), .ZN(new_n836));
  NOR4_X1   g650(.A1(new_n706), .A2(new_n707), .A3(new_n692), .A4(new_n701), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n831), .B(new_n835), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n711), .A2(KEYINPUT52), .A3(new_n831), .A4(new_n835), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n772), .A2(new_n822), .A3(new_n843), .A4(new_n828), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n830), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n848));
  INV_X1    g662(.A(new_n829), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n842), .A2(new_n849), .A3(KEYINPUT53), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n847), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n845), .A2(new_n852), .A3(new_n846), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n852), .B1(new_n845), .B2(new_n846), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n845), .A2(new_n846), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n851), .B1(new_n856), .B2(new_n848), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n782), .A2(new_n493), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n750), .A2(new_n734), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n656), .A2(new_n684), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n811), .A2(new_n388), .A3(new_n493), .A4(new_n859), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n779), .A2(new_n641), .ZN(new_n863));
  OAI22_X1  g677(.A1(new_n860), .A2(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n858), .A2(new_n666), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n724), .A2(new_n503), .A3(new_n734), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n867), .A2(KEYINPUT50), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(KEYINPUT50), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n864), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n731), .A2(new_n732), .A3(new_n577), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n750), .B(new_n865), .C1(new_n804), .C2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT51), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n873), .B(new_n874), .ZN(new_n875));
  OR2_X1    g689(.A1(new_n759), .A2(new_n760), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n876), .A2(new_n859), .A3(new_n858), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT48), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n862), .A2(new_n643), .ZN(new_n879));
  INV_X1    g693(.A(G952), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n879), .A2(new_n880), .A3(G953), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n865), .A2(new_n741), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n882), .A2(KEYINPUT119), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n882), .A2(KEYINPUT119), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n878), .B(new_n881), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n885), .B(KEYINPUT120), .Z(new_n886));
  NOR3_X1   g700(.A1(new_n857), .A2(new_n875), .A3(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(G952), .A2(G953), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n813), .B1(new_n887), .B2(new_n888), .ZN(G75));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT56), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n847), .A2(new_n850), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n313), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n891), .B1(new_n893), .B2(new_n572), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n564), .A2(new_n566), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(new_n560), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT55), .Z(new_n897));
  NAND2_X1  g711(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n364), .A2(G952), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n894), .A2(new_n897), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n890), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n899), .B1(new_n894), .B2(new_n897), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n904), .B(KEYINPUT121), .C1(new_n894), .C2(new_n897), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n903), .A2(new_n905), .ZN(G51));
  NAND3_X1  g720(.A1(new_n892), .A2(new_n313), .A3(new_n793), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT122), .Z(new_n908));
  NAND2_X1  g722(.A1(new_n892), .A2(KEYINPUT54), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n851), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n623), .B(KEYINPUT57), .Z(new_n912));
  OAI21_X1  g726(.A(new_n614), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n899), .B1(new_n908), .B2(new_n913), .ZN(G54));
  NAND4_X1  g728(.A1(new_n892), .A2(KEYINPUT58), .A3(G475), .A4(new_n313), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n915), .A2(new_n485), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n915), .A2(new_n485), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n916), .A2(new_n917), .A3(new_n899), .ZN(G60));
  NAND2_X1  g732(.A1(G478), .A2(G902), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT59), .Z(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n639), .B1(new_n857), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n920), .B1(new_n637), .B2(new_n638), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n899), .B1(new_n910), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(KEYINPUT123), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT123), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n845), .A2(new_n846), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n845), .A2(new_n846), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n928), .B1(new_n929), .B2(new_n852), .ZN(new_n930));
  OAI21_X1  g744(.A(KEYINPUT54), .B1(new_n930), .B2(new_n853), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n920), .B1(new_n931), .B2(new_n851), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n927), .B(new_n924), .C1(new_n932), .C2(new_n639), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n926), .A2(new_n933), .ZN(G63));
  NAND2_X1  g748(.A1(G217), .A2(G902), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT60), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n936), .B1(new_n847), .B2(new_n850), .ZN(new_n937));
  OR2_X1    g751(.A1(new_n937), .A2(new_n373), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n681), .A2(new_n682), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n899), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(KEYINPUT124), .B1(new_n937), .B2(new_n939), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n942), .A2(KEYINPUT61), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n941), .B(new_n943), .ZN(G66));
  OAI21_X1  g758(.A(G953), .B1(new_n497), .B2(new_n537), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n945), .B1(new_n822), .B2(G953), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n895), .B1(G898), .B2(new_n364), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(G69));
  NOR2_X1   g762(.A1(new_n266), .A2(new_n274), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(new_n476), .Z(new_n950));
  AND2_X1   g764(.A1(new_n711), .A2(new_n831), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n726), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT62), .ZN(new_n953));
  INV_X1    g767(.A(new_n806), .ZN(new_n954));
  INV_X1    g768(.A(new_n764), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n714), .A2(new_n503), .A3(new_n722), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n955), .B(new_n956), .C1(new_n751), .C2(new_n816), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT125), .ZN(new_n958));
  NOR4_X1   g772(.A1(new_n801), .A2(new_n953), .A3(new_n954), .A4(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n950), .B1(new_n959), .B2(G953), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n806), .A2(new_n777), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n799), .A2(new_n876), .A3(new_n834), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n961), .A2(new_n772), .A3(new_n951), .A4(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n963), .A2(new_n801), .ZN(new_n964));
  MUX2_X1   g778(.A(G900), .B(new_n964), .S(new_n364), .Z(new_n965));
  OAI21_X1  g779(.A(new_n960), .B1(new_n965), .B2(new_n950), .ZN(new_n966));
  INV_X1    g780(.A(G227), .ZN(new_n967));
  OAI21_X1  g781(.A(G953), .B1(new_n967), .B2(new_n697), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT126), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n969), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n971), .B(new_n960), .C1(new_n965), .C2(new_n950), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n970), .A2(new_n972), .ZN(G72));
  NAND3_X1  g787(.A1(new_n275), .A2(new_n249), .A3(new_n254), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n974), .A2(new_n259), .ZN(new_n975));
  NOR4_X1   g789(.A1(new_n963), .A2(new_n801), .A3(new_n814), .A4(new_n821), .ZN(new_n976));
  NAND2_X1  g790(.A1(G472), .A2(G902), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT63), .Z(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n975), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n979), .B1(new_n959), .B2(new_n822), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n974), .A2(new_n259), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n980), .B(new_n900), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n856), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n306), .B(new_n310), .C1(new_n291), .C2(new_n285), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n985), .A2(new_n978), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n983), .B1(new_n984), .B2(new_n986), .ZN(G57));
endmodule


