

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U548 ( .A1(n523), .A2(G2104), .ZN(n878) );
  NOR2_X1 U549 ( .A1(G651), .A2(G543), .ZN(n649) );
  NOR2_X1 U550 ( .A1(G651), .A2(n645), .ZN(n653) );
  INV_X1 U551 ( .A(KEYINPUT86), .ZN(n531) );
  NOR2_X1 U552 ( .A1(n527), .A2(n526), .ZN(G160) );
  XOR2_X1 U553 ( .A(KEYINPUT68), .B(n580), .Z(n516) );
  NOR2_X1 U554 ( .A1(n691), .A2(n913), .ZN(n693) );
  NOR2_X1 U555 ( .A1(n693), .A2(n928), .ZN(n692) );
  XNOR2_X1 U556 ( .A(KEYINPUT100), .B(KEYINPUT30), .ZN(n720) );
  XNOR2_X1 U557 ( .A(n721), .B(n720), .ZN(n722) );
  INV_X1 U558 ( .A(KEYINPUT29), .ZN(n709) );
  XNOR2_X1 U559 ( .A(n710), .B(n709), .ZN(n716) );
  INV_X1 U560 ( .A(n712), .ZN(n731) );
  NOR2_X1 U561 ( .A1(G164), .A2(G1384), .ZN(n798) );
  NAND2_X1 U562 ( .A1(n877), .A2(G138), .ZN(n530) );
  INV_X1 U563 ( .A(KEYINPUT17), .ZN(n521) );
  XNOR2_X1 U564 ( .A(n584), .B(KEYINPUT15), .ZN(n928) );
  AND2_X1 U565 ( .A1(G2105), .A2(G2104), .ZN(n882) );
  NAND2_X1 U566 ( .A1(G113), .A2(n882), .ZN(n517) );
  XNOR2_X1 U567 ( .A(n517), .B(KEYINPUT64), .ZN(n520) );
  INV_X1 U568 ( .A(G2105), .ZN(n523) );
  NAND2_X1 U569 ( .A1(G101), .A2(n878), .ZN(n518) );
  XOR2_X1 U570 ( .A(KEYINPUT23), .B(n518), .Z(n519) );
  NAND2_X1 U571 ( .A1(n520), .A2(n519), .ZN(n527) );
  NOR2_X1 U572 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  XNOR2_X2 U573 ( .A(n522), .B(n521), .ZN(n877) );
  NAND2_X1 U574 ( .A1(G137), .A2(n877), .ZN(n525) );
  NOR2_X2 U575 ( .A1(G2104), .A2(n523), .ZN(n881) );
  NAND2_X1 U576 ( .A1(G125), .A2(n881), .ZN(n524) );
  NAND2_X1 U577 ( .A1(n525), .A2(n524), .ZN(n526) );
  NAND2_X1 U578 ( .A1(n881), .A2(G126), .ZN(n528) );
  XNOR2_X1 U579 ( .A(n528), .B(KEYINPUT84), .ZN(n534) );
  NAND2_X1 U580 ( .A1(G102), .A2(n878), .ZN(n529) );
  NAND2_X1 U581 ( .A1(n530), .A2(n529), .ZN(n532) );
  XNOR2_X1 U582 ( .A(n532), .B(n531), .ZN(n533) );
  NAND2_X1 U583 ( .A1(n534), .A2(n533), .ZN(n537) );
  NAND2_X1 U584 ( .A1(G114), .A2(n882), .ZN(n535) );
  XNOR2_X1 U585 ( .A(KEYINPUT85), .B(n535), .ZN(n536) );
  NOR2_X1 U586 ( .A1(n537), .A2(n536), .ZN(G164) );
  XOR2_X1 U587 ( .A(G2443), .B(G2446), .Z(n539) );
  XNOR2_X1 U588 ( .A(G2427), .B(G2451), .ZN(n538) );
  XNOR2_X1 U589 ( .A(n539), .B(n538), .ZN(n545) );
  XOR2_X1 U590 ( .A(G2430), .B(G2454), .Z(n541) );
  XNOR2_X1 U591 ( .A(G1348), .B(G1341), .ZN(n540) );
  XNOR2_X1 U592 ( .A(n541), .B(n540), .ZN(n543) );
  XOR2_X1 U593 ( .A(G2435), .B(G2438), .Z(n542) );
  XNOR2_X1 U594 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U595 ( .A(n545), .B(n544), .Z(n546) );
  AND2_X1 U596 ( .A1(G14), .A2(n546), .ZN(G401) );
  AND2_X1 U597 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U598 ( .A1(G123), .A2(n881), .ZN(n547) );
  XNOR2_X1 U599 ( .A(n547), .B(KEYINPUT18), .ZN(n555) );
  NAND2_X1 U600 ( .A1(G111), .A2(n882), .ZN(n548) );
  XNOR2_X1 U601 ( .A(n548), .B(KEYINPUT74), .ZN(n550) );
  NAND2_X1 U602 ( .A1(n877), .A2(G135), .ZN(n549) );
  NAND2_X1 U603 ( .A1(n550), .A2(n549), .ZN(n553) );
  NAND2_X1 U604 ( .A1(G99), .A2(n878), .ZN(n551) );
  XNOR2_X1 U605 ( .A(KEYINPUT75), .B(n551), .ZN(n552) );
  NOR2_X1 U606 ( .A1(n553), .A2(n552), .ZN(n554) );
  NAND2_X1 U607 ( .A1(n555), .A2(n554), .ZN(n993) );
  XNOR2_X1 U608 ( .A(G2096), .B(n993), .ZN(n556) );
  OR2_X1 U609 ( .A1(G2100), .A2(n556), .ZN(G156) );
  INV_X1 U610 ( .A(G57), .ZN(G237) );
  INV_X1 U611 ( .A(G132), .ZN(G219) );
  INV_X1 U612 ( .A(G82), .ZN(G220) );
  INV_X1 U613 ( .A(G96), .ZN(G221) );
  INV_X1 U614 ( .A(G651), .ZN(n560) );
  NOR2_X1 U615 ( .A1(G543), .A2(n560), .ZN(n557) );
  XOR2_X2 U616 ( .A(KEYINPUT1), .B(n557), .Z(n652) );
  NAND2_X1 U617 ( .A1(G64), .A2(n652), .ZN(n559) );
  XOR2_X1 U618 ( .A(G543), .B(KEYINPUT0), .Z(n645) );
  NAND2_X1 U619 ( .A1(G52), .A2(n653), .ZN(n558) );
  NAND2_X1 U620 ( .A1(n559), .A2(n558), .ZN(n565) );
  NOR2_X1 U621 ( .A1(n645), .A2(n560), .ZN(n648) );
  NAND2_X1 U622 ( .A1(G77), .A2(n648), .ZN(n562) );
  NAND2_X1 U623 ( .A1(G90), .A2(n649), .ZN(n561) );
  NAND2_X1 U624 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U625 ( .A(KEYINPUT9), .B(n563), .Z(n564) );
  NOR2_X1 U626 ( .A1(n565), .A2(n564), .ZN(G171) );
  NAND2_X1 U627 ( .A1(G7), .A2(G661), .ZN(n566) );
  XNOR2_X1 U628 ( .A(n566), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U629 ( .A(G223), .ZN(n829) );
  NAND2_X1 U630 ( .A1(n829), .A2(G567), .ZN(n567) );
  XOR2_X1 U631 ( .A(KEYINPUT11), .B(n567), .Z(G234) );
  NAND2_X1 U632 ( .A1(n649), .A2(G81), .ZN(n568) );
  XNOR2_X1 U633 ( .A(n568), .B(KEYINPUT12), .ZN(n570) );
  NAND2_X1 U634 ( .A1(G68), .A2(n648), .ZN(n569) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(KEYINPUT13), .B(n571), .ZN(n577) );
  NAND2_X1 U637 ( .A1(G56), .A2(n652), .ZN(n572) );
  XOR2_X1 U638 ( .A(KEYINPUT14), .B(n572), .Z(n575) );
  NAND2_X1 U639 ( .A1(G43), .A2(n653), .ZN(n573) );
  XNOR2_X1 U640 ( .A(KEYINPUT67), .B(n573), .ZN(n574) );
  NOR2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n913) );
  INV_X1 U643 ( .A(G860), .ZN(n608) );
  OR2_X1 U644 ( .A1(n913), .A2(n608), .ZN(G153) );
  INV_X1 U645 ( .A(G171), .ZN(G301) );
  NAND2_X1 U646 ( .A1(G868), .A2(G301), .ZN(n586) );
  NAND2_X1 U647 ( .A1(G54), .A2(n653), .ZN(n583) );
  NAND2_X1 U648 ( .A1(G79), .A2(n648), .ZN(n579) );
  NAND2_X1 U649 ( .A1(G92), .A2(n649), .ZN(n578) );
  NAND2_X1 U650 ( .A1(n579), .A2(n578), .ZN(n581) );
  NAND2_X1 U651 ( .A1(n652), .A2(G66), .ZN(n580) );
  NOR2_X1 U652 ( .A1(n581), .A2(n516), .ZN(n582) );
  NAND2_X1 U653 ( .A1(n583), .A2(n582), .ZN(n584) );
  OR2_X1 U654 ( .A1(n928), .A2(G868), .ZN(n585) );
  NAND2_X1 U655 ( .A1(n586), .A2(n585), .ZN(G284) );
  NAND2_X1 U656 ( .A1(G63), .A2(n652), .ZN(n588) );
  NAND2_X1 U657 ( .A1(G51), .A2(n653), .ZN(n587) );
  NAND2_X1 U658 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U659 ( .A(KEYINPUT6), .B(n589), .ZN(n595) );
  NAND2_X1 U660 ( .A1(n649), .A2(G89), .ZN(n590) );
  XNOR2_X1 U661 ( .A(n590), .B(KEYINPUT4), .ZN(n592) );
  NAND2_X1 U662 ( .A1(G76), .A2(n648), .ZN(n591) );
  NAND2_X1 U663 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U664 ( .A(n593), .B(KEYINPUT5), .Z(n594) );
  NOR2_X1 U665 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U666 ( .A(KEYINPUT69), .B(n596), .Z(n597) );
  XOR2_X1 U667 ( .A(KEYINPUT7), .B(n597), .Z(G168) );
  XOR2_X1 U668 ( .A(G168), .B(KEYINPUT8), .Z(n598) );
  XNOR2_X1 U669 ( .A(KEYINPUT70), .B(n598), .ZN(G286) );
  NAND2_X1 U670 ( .A1(G65), .A2(n652), .ZN(n600) );
  NAND2_X1 U671 ( .A1(G53), .A2(n653), .ZN(n599) );
  NAND2_X1 U672 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U673 ( .A1(G78), .A2(n648), .ZN(n602) );
  NAND2_X1 U674 ( .A1(G91), .A2(n649), .ZN(n601) );
  NAND2_X1 U675 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U676 ( .A1(n604), .A2(n603), .ZN(n916) );
  INV_X1 U677 ( .A(n916), .ZN(G299) );
  XNOR2_X1 U678 ( .A(KEYINPUT71), .B(G868), .ZN(n605) );
  NOR2_X1 U679 ( .A1(G286), .A2(n605), .ZN(n607) );
  NOR2_X1 U680 ( .A1(G868), .A2(G299), .ZN(n606) );
  NOR2_X1 U681 ( .A1(n607), .A2(n606), .ZN(G297) );
  NAND2_X1 U682 ( .A1(G559), .A2(n608), .ZN(n609) );
  XNOR2_X1 U683 ( .A(KEYINPUT72), .B(n609), .ZN(n610) );
  NAND2_X1 U684 ( .A1(n610), .A2(n928), .ZN(n611) );
  XNOR2_X1 U685 ( .A(KEYINPUT16), .B(n611), .ZN(G148) );
  NAND2_X1 U686 ( .A1(n928), .A2(G868), .ZN(n612) );
  NOR2_X1 U687 ( .A1(G559), .A2(n612), .ZN(n613) );
  XOR2_X1 U688 ( .A(KEYINPUT73), .B(n613), .Z(n615) );
  NOR2_X1 U689 ( .A1(G868), .A2(n913), .ZN(n614) );
  NOR2_X1 U690 ( .A1(n615), .A2(n614), .ZN(G282) );
  NAND2_X1 U691 ( .A1(G559), .A2(n928), .ZN(n616) );
  XNOR2_X1 U692 ( .A(n616), .B(n913), .ZN(n665) );
  NOR2_X1 U693 ( .A1(G860), .A2(n665), .ZN(n625) );
  NAND2_X1 U694 ( .A1(n652), .A2(G67), .ZN(n619) );
  NAND2_X1 U695 ( .A1(G80), .A2(n648), .ZN(n617) );
  XOR2_X1 U696 ( .A(KEYINPUT77), .B(n617), .Z(n618) );
  NAND2_X1 U697 ( .A1(n619), .A2(n618), .ZN(n623) );
  NAND2_X1 U698 ( .A1(G93), .A2(n649), .ZN(n621) );
  NAND2_X1 U699 ( .A1(G55), .A2(n653), .ZN(n620) );
  NAND2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U701 ( .A1(n623), .A2(n622), .ZN(n661) );
  XNOR2_X1 U702 ( .A(n661), .B(KEYINPUT76), .ZN(n624) );
  XNOR2_X1 U703 ( .A(n625), .B(n624), .ZN(G145) );
  NAND2_X1 U704 ( .A1(n649), .A2(G85), .ZN(n632) );
  NAND2_X1 U705 ( .A1(G60), .A2(n652), .ZN(n627) );
  NAND2_X1 U706 ( .A1(G47), .A2(n653), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U708 ( .A1(G72), .A2(n648), .ZN(n628) );
  XNOR2_X1 U709 ( .A(KEYINPUT65), .B(n628), .ZN(n629) );
  NOR2_X1 U710 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U711 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U712 ( .A(n633), .B(KEYINPUT66), .ZN(G290) );
  NAND2_X1 U713 ( .A1(G86), .A2(n649), .ZN(n635) );
  NAND2_X1 U714 ( .A1(G61), .A2(n652), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n648), .A2(G73), .ZN(n636) );
  XOR2_X1 U717 ( .A(KEYINPUT2), .B(n636), .Z(n637) );
  NOR2_X1 U718 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n653), .A2(G48), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n640), .A2(n639), .ZN(G305) );
  NAND2_X1 U721 ( .A1(G49), .A2(n653), .ZN(n642) );
  NAND2_X1 U722 ( .A1(G74), .A2(G651), .ZN(n641) );
  NAND2_X1 U723 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U724 ( .A1(n652), .A2(n643), .ZN(n644) );
  XNOR2_X1 U725 ( .A(n644), .B(KEYINPUT78), .ZN(n647) );
  NAND2_X1 U726 ( .A1(G87), .A2(n645), .ZN(n646) );
  NAND2_X1 U727 ( .A1(n647), .A2(n646), .ZN(G288) );
  NAND2_X1 U728 ( .A1(G75), .A2(n648), .ZN(n651) );
  NAND2_X1 U729 ( .A1(G88), .A2(n649), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n651), .A2(n650), .ZN(n657) );
  NAND2_X1 U731 ( .A1(G62), .A2(n652), .ZN(n655) );
  NAND2_X1 U732 ( .A1(G50), .A2(n653), .ZN(n654) );
  NAND2_X1 U733 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U734 ( .A1(n657), .A2(n656), .ZN(G166) );
  NOR2_X1 U735 ( .A1(G868), .A2(n661), .ZN(n658) );
  XNOR2_X1 U736 ( .A(n658), .B(KEYINPUT79), .ZN(n668) );
  XNOR2_X1 U737 ( .A(n916), .B(G305), .ZN(n659) );
  XNOR2_X1 U738 ( .A(n659), .B(G288), .ZN(n660) );
  XOR2_X1 U739 ( .A(n661), .B(n660), .Z(n663) );
  XNOR2_X1 U740 ( .A(G166), .B(KEYINPUT19), .ZN(n662) );
  XNOR2_X1 U741 ( .A(n663), .B(n662), .ZN(n664) );
  XOR2_X1 U742 ( .A(G290), .B(n664), .Z(n900) );
  XNOR2_X1 U743 ( .A(n900), .B(n665), .ZN(n666) );
  NAND2_X1 U744 ( .A1(G868), .A2(n666), .ZN(n667) );
  NAND2_X1 U745 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U746 ( .A1(G2078), .A2(G2084), .ZN(n669) );
  XOR2_X1 U747 ( .A(KEYINPUT20), .B(n669), .Z(n670) );
  NAND2_X1 U748 ( .A1(G2090), .A2(n670), .ZN(n671) );
  XNOR2_X1 U749 ( .A(KEYINPUT21), .B(n671), .ZN(n672) );
  NAND2_X1 U750 ( .A1(n672), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U751 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U752 ( .A1(G220), .A2(G219), .ZN(n673) );
  XOR2_X1 U753 ( .A(KEYINPUT22), .B(n673), .Z(n674) );
  NOR2_X1 U754 ( .A1(G218), .A2(n674), .ZN(n675) );
  XOR2_X1 U755 ( .A(KEYINPUT80), .B(n675), .Z(n676) );
  NOR2_X1 U756 ( .A1(G221), .A2(n676), .ZN(n677) );
  XNOR2_X1 U757 ( .A(KEYINPUT81), .B(n677), .ZN(n833) );
  NAND2_X1 U758 ( .A1(n833), .A2(G2106), .ZN(n682) );
  NAND2_X1 U759 ( .A1(G120), .A2(G69), .ZN(n678) );
  NOR2_X1 U760 ( .A1(G237), .A2(n678), .ZN(n679) );
  XNOR2_X1 U761 ( .A(KEYINPUT82), .B(n679), .ZN(n680) );
  NAND2_X1 U762 ( .A1(n680), .A2(G108), .ZN(n834) );
  NAND2_X1 U763 ( .A1(G567), .A2(n834), .ZN(n681) );
  NAND2_X1 U764 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U765 ( .A(n683), .B(KEYINPUT83), .ZN(G319) );
  INV_X1 U766 ( .A(G319), .ZN(n685) );
  NAND2_X1 U767 ( .A1(G661), .A2(G483), .ZN(n684) );
  NOR2_X1 U768 ( .A1(n685), .A2(n684), .ZN(n832) );
  NAND2_X1 U769 ( .A1(n832), .A2(G36), .ZN(G176) );
  INV_X1 U770 ( .A(G166), .ZN(G303) );
  INV_X1 U771 ( .A(n798), .ZN(n686) );
  NAND2_X1 U772 ( .A1(G160), .A2(G40), .ZN(n797) );
  NOR2_X2 U773 ( .A1(n686), .A2(n797), .ZN(n712) );
  AND2_X1 U774 ( .A1(n712), .A2(G1996), .ZN(n688) );
  XOR2_X1 U775 ( .A(KEYINPUT26), .B(KEYINPUT98), .Z(n687) );
  XNOR2_X1 U776 ( .A(n688), .B(n687), .ZN(n690) );
  NAND2_X1 U777 ( .A1(n731), .A2(G1341), .ZN(n689) );
  NAND2_X1 U778 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U779 ( .A(n692), .B(KEYINPUT99), .ZN(n699) );
  NAND2_X1 U780 ( .A1(n693), .A2(n928), .ZN(n697) );
  NOR2_X1 U781 ( .A1(n712), .A2(G1348), .ZN(n695) );
  NOR2_X1 U782 ( .A1(G2067), .A2(n731), .ZN(n694) );
  NOR2_X1 U783 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U784 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U785 ( .A1(n699), .A2(n698), .ZN(n704) );
  NAND2_X1 U786 ( .A1(n712), .A2(G2072), .ZN(n700) );
  XNOR2_X1 U787 ( .A(n700), .B(KEYINPUT27), .ZN(n702) );
  XNOR2_X1 U788 ( .A(G1956), .B(KEYINPUT97), .ZN(n937) );
  NOR2_X1 U789 ( .A1(n937), .A2(n712), .ZN(n701) );
  NOR2_X1 U790 ( .A1(n702), .A2(n701), .ZN(n705) );
  NAND2_X1 U791 ( .A1(n916), .A2(n705), .ZN(n703) );
  NAND2_X1 U792 ( .A1(n704), .A2(n703), .ZN(n708) );
  NOR2_X1 U793 ( .A1(n916), .A2(n705), .ZN(n706) );
  XOR2_X1 U794 ( .A(n706), .B(KEYINPUT28), .Z(n707) );
  NAND2_X1 U795 ( .A1(n708), .A2(n707), .ZN(n710) );
  NOR2_X1 U796 ( .A1(n712), .A2(G1961), .ZN(n711) );
  XOR2_X1 U797 ( .A(KEYINPUT96), .B(n711), .Z(n714) );
  XNOR2_X1 U798 ( .A(G2078), .B(KEYINPUT25), .ZN(n970) );
  NAND2_X1 U799 ( .A1(n712), .A2(n970), .ZN(n713) );
  NAND2_X1 U800 ( .A1(n714), .A2(n713), .ZN(n723) );
  NAND2_X1 U801 ( .A1(n723), .A2(G171), .ZN(n715) );
  NAND2_X1 U802 ( .A1(n716), .A2(n715), .ZN(n729) );
  INV_X1 U803 ( .A(G1966), .ZN(n717) );
  AND2_X1 U804 ( .A1(G8), .A2(n717), .ZN(n718) );
  AND2_X1 U805 ( .A1(n731), .A2(n718), .ZN(n743) );
  NOR2_X1 U806 ( .A1(G2084), .A2(n731), .ZN(n740) );
  NOR2_X1 U807 ( .A1(n743), .A2(n740), .ZN(n719) );
  NAND2_X1 U808 ( .A1(n719), .A2(G8), .ZN(n721) );
  NOR2_X1 U809 ( .A1(n722), .A2(G168), .ZN(n725) );
  NOR2_X1 U810 ( .A1(G171), .A2(n723), .ZN(n724) );
  NOR2_X1 U811 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U812 ( .A(n726), .B(KEYINPUT31), .ZN(n727) );
  XNOR2_X1 U813 ( .A(n727), .B(KEYINPUT101), .ZN(n728) );
  NAND2_X1 U814 ( .A1(n729), .A2(n728), .ZN(n742) );
  NAND2_X1 U815 ( .A1(n742), .A2(G286), .ZN(n730) );
  XNOR2_X1 U816 ( .A(n730), .B(KEYINPUT102), .ZN(n737) );
  NAND2_X1 U817 ( .A1(n731), .A2(G8), .ZN(n762) );
  NOR2_X1 U818 ( .A1(G1971), .A2(n762), .ZN(n733) );
  NOR2_X1 U819 ( .A1(G2090), .A2(n731), .ZN(n732) );
  NOR2_X1 U820 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U821 ( .A1(n734), .A2(G303), .ZN(n735) );
  XOR2_X1 U822 ( .A(KEYINPUT103), .B(n735), .Z(n736) );
  NAND2_X1 U823 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U824 ( .A1(n738), .A2(G8), .ZN(n739) );
  XNOR2_X1 U825 ( .A(n739), .B(KEYINPUT32), .ZN(n748) );
  NAND2_X1 U826 ( .A1(G8), .A2(n740), .ZN(n741) );
  XOR2_X1 U827 ( .A(KEYINPUT95), .B(n741), .Z(n746) );
  INV_X1 U828 ( .A(n742), .ZN(n744) );
  NOR2_X1 U829 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U830 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U831 ( .A1(n748), .A2(n747), .ZN(n760) );
  NOR2_X1 U832 ( .A1(G2090), .A2(G303), .ZN(n749) );
  NAND2_X1 U833 ( .A1(G8), .A2(n749), .ZN(n750) );
  NAND2_X1 U834 ( .A1(n760), .A2(n750), .ZN(n751) );
  XNOR2_X1 U835 ( .A(n751), .B(KEYINPUT106), .ZN(n752) );
  NAND2_X1 U836 ( .A1(n752), .A2(n762), .ZN(n753) );
  XNOR2_X1 U837 ( .A(KEYINPUT107), .B(n753), .ZN(n775) );
  XNOR2_X1 U838 ( .A(G1981), .B(G305), .ZN(n911) );
  INV_X1 U839 ( .A(KEYINPUT33), .ZN(n758) );
  INV_X1 U840 ( .A(n762), .ZN(n770) );
  NOR2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n757) );
  NAND2_X1 U842 ( .A1(n770), .A2(n757), .ZN(n754) );
  NOR2_X1 U843 ( .A1(n758), .A2(n754), .ZN(n755) );
  XNOR2_X1 U844 ( .A(n755), .B(KEYINPUT105), .ZN(n767) );
  NOR2_X1 U845 ( .A1(G1971), .A2(G303), .ZN(n756) );
  NOR2_X1 U846 ( .A1(n757), .A2(n756), .ZN(n922) );
  AND2_X1 U847 ( .A1(n922), .A2(n758), .ZN(n759) );
  NAND2_X1 U848 ( .A1(n760), .A2(n759), .ZN(n765) );
  NAND2_X1 U849 ( .A1(G288), .A2(G1976), .ZN(n761) );
  XOR2_X1 U850 ( .A(KEYINPUT104), .B(n761), .Z(n920) );
  NOR2_X1 U851 ( .A1(n762), .A2(n920), .ZN(n763) );
  OR2_X1 U852 ( .A1(KEYINPUT33), .A2(n763), .ZN(n764) );
  AND2_X1 U853 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U854 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U855 ( .A1(n911), .A2(n768), .ZN(n773) );
  NOR2_X1 U856 ( .A1(G1981), .A2(G305), .ZN(n769) );
  XNOR2_X1 U857 ( .A(n769), .B(KEYINPUT24), .ZN(n771) );
  AND2_X1 U858 ( .A1(n771), .A2(n770), .ZN(n772) );
  OR2_X1 U859 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U860 ( .A1(n775), .A2(n774), .ZN(n811) );
  NAND2_X1 U861 ( .A1(n882), .A2(G107), .ZN(n776) );
  XNOR2_X1 U862 ( .A(KEYINPUT88), .B(n776), .ZN(n779) );
  NAND2_X1 U863 ( .A1(n881), .A2(G119), .ZN(n777) );
  XOR2_X1 U864 ( .A(KEYINPUT87), .B(n777), .Z(n778) );
  NAND2_X1 U865 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U866 ( .A(KEYINPUT89), .B(n780), .ZN(n784) );
  NAND2_X1 U867 ( .A1(G131), .A2(n877), .ZN(n782) );
  NAND2_X1 U868 ( .A1(G95), .A2(n878), .ZN(n781) );
  AND2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U870 ( .A1(n784), .A2(n783), .ZN(n873) );
  XNOR2_X1 U871 ( .A(KEYINPUT90), .B(G1991), .ZN(n965) );
  NAND2_X1 U872 ( .A1(n873), .A2(n965), .ZN(n796) );
  NAND2_X1 U873 ( .A1(n878), .A2(G105), .ZN(n787) );
  XOR2_X1 U874 ( .A(KEYINPUT38), .B(KEYINPUT92), .Z(n785) );
  XNOR2_X1 U875 ( .A(KEYINPUT91), .B(n785), .ZN(n786) );
  XNOR2_X1 U876 ( .A(n787), .B(n786), .ZN(n794) );
  NAND2_X1 U877 ( .A1(G129), .A2(n881), .ZN(n789) );
  NAND2_X1 U878 ( .A1(G117), .A2(n882), .ZN(n788) );
  NAND2_X1 U879 ( .A1(n789), .A2(n788), .ZN(n792) );
  NAND2_X1 U880 ( .A1(G141), .A2(n877), .ZN(n790) );
  XNOR2_X1 U881 ( .A(KEYINPUT93), .B(n790), .ZN(n791) );
  NOR2_X1 U882 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U883 ( .A1(n794), .A2(n793), .ZN(n894) );
  NAND2_X1 U884 ( .A1(G1996), .A2(n894), .ZN(n795) );
  NAND2_X1 U885 ( .A1(n796), .A2(n795), .ZN(n996) );
  NOR2_X1 U886 ( .A1(n798), .A2(n797), .ZN(n824) );
  NAND2_X1 U887 ( .A1(n996), .A2(n824), .ZN(n799) );
  XOR2_X1 U888 ( .A(KEYINPUT94), .B(n799), .Z(n816) );
  INV_X1 U889 ( .A(n816), .ZN(n809) );
  XNOR2_X1 U890 ( .A(KEYINPUT37), .B(G2067), .ZN(n821) );
  NAND2_X1 U891 ( .A1(G140), .A2(n877), .ZN(n801) );
  NAND2_X1 U892 ( .A1(G104), .A2(n878), .ZN(n800) );
  NAND2_X1 U893 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U894 ( .A(KEYINPUT34), .B(n802), .ZN(n807) );
  NAND2_X1 U895 ( .A1(G128), .A2(n881), .ZN(n804) );
  NAND2_X1 U896 ( .A1(G116), .A2(n882), .ZN(n803) );
  NAND2_X1 U897 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U898 ( .A(KEYINPUT35), .B(n805), .Z(n806) );
  NOR2_X1 U899 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U900 ( .A(KEYINPUT36), .B(n808), .ZN(n889) );
  NOR2_X1 U901 ( .A1(n821), .A2(n889), .ZN(n990) );
  NAND2_X1 U902 ( .A1(n824), .A2(n990), .ZN(n819) );
  NAND2_X1 U903 ( .A1(n809), .A2(n819), .ZN(n810) );
  NOR2_X1 U904 ( .A1(n811), .A2(n810), .ZN(n813) );
  XNOR2_X1 U905 ( .A(G1986), .B(G290), .ZN(n924) );
  NAND2_X1 U906 ( .A1(n924), .A2(n824), .ZN(n812) );
  NAND2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n827) );
  NOR2_X1 U908 ( .A1(G1996), .A2(n894), .ZN(n1004) );
  NOR2_X1 U909 ( .A1(G1986), .A2(G290), .ZN(n814) );
  NOR2_X1 U910 ( .A1(n965), .A2(n873), .ZN(n992) );
  NOR2_X1 U911 ( .A1(n814), .A2(n992), .ZN(n815) );
  NOR2_X1 U912 ( .A1(n816), .A2(n815), .ZN(n817) );
  NOR2_X1 U913 ( .A1(n1004), .A2(n817), .ZN(n818) );
  XNOR2_X1 U914 ( .A(n818), .B(KEYINPUT39), .ZN(n820) );
  NAND2_X1 U915 ( .A1(n820), .A2(n819), .ZN(n822) );
  NAND2_X1 U916 ( .A1(n821), .A2(n889), .ZN(n988) );
  NAND2_X1 U917 ( .A1(n822), .A2(n988), .ZN(n823) );
  XNOR2_X1 U918 ( .A(KEYINPUT108), .B(n823), .ZN(n825) );
  NAND2_X1 U919 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U920 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U921 ( .A(n828), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n829), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n830) );
  NAND2_X1 U924 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U926 ( .A1(n832), .A2(n831), .ZN(G188) );
  INV_X1 U928 ( .A(G120), .ZN(G236) );
  INV_X1 U929 ( .A(G108), .ZN(G238) );
  INV_X1 U930 ( .A(G69), .ZN(G235) );
  NOR2_X1 U931 ( .A1(n834), .A2(n833), .ZN(n835) );
  XNOR2_X1 U932 ( .A(n835), .B(KEYINPUT109), .ZN(G261) );
  INV_X1 U933 ( .A(G261), .ZN(G325) );
  XOR2_X1 U934 ( .A(G1966), .B(G1981), .Z(n837) );
  XNOR2_X1 U935 ( .A(G1996), .B(G1991), .ZN(n836) );
  XNOR2_X1 U936 ( .A(n837), .B(n836), .ZN(n847) );
  XOR2_X1 U937 ( .A(KEYINPUT111), .B(KEYINPUT41), .Z(n839) );
  XNOR2_X1 U938 ( .A(G1956), .B(KEYINPUT113), .ZN(n838) );
  XNOR2_X1 U939 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U940 ( .A(G1961), .B(G1971), .Z(n841) );
  XNOR2_X1 U941 ( .A(G1986), .B(G1976), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U943 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U944 ( .A(KEYINPUT112), .B(G2474), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U946 ( .A(n847), .B(n846), .Z(G229) );
  XOR2_X1 U947 ( .A(G2096), .B(KEYINPUT43), .Z(n849) );
  XNOR2_X1 U948 ( .A(G2072), .B(KEYINPUT110), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U950 ( .A(n850), .B(G2678), .Z(n852) );
  XNOR2_X1 U951 ( .A(G2067), .B(G2090), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U953 ( .A(KEYINPUT42), .B(G2100), .Z(n854) );
  XNOR2_X1 U954 ( .A(G2078), .B(G2084), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(G227) );
  NAND2_X1 U957 ( .A1(G136), .A2(n877), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n857), .B(KEYINPUT114), .ZN(n864) );
  NAND2_X1 U959 ( .A1(G100), .A2(n878), .ZN(n859) );
  NAND2_X1 U960 ( .A1(G112), .A2(n882), .ZN(n858) );
  NAND2_X1 U961 ( .A1(n859), .A2(n858), .ZN(n862) );
  NAND2_X1 U962 ( .A1(n881), .A2(G124), .ZN(n860) );
  XOR2_X1 U963 ( .A(KEYINPUT44), .B(n860), .Z(n861) );
  NOR2_X1 U964 ( .A1(n862), .A2(n861), .ZN(n863) );
  NAND2_X1 U965 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U966 ( .A(KEYINPUT115), .B(n865), .ZN(G162) );
  NAND2_X1 U967 ( .A1(G130), .A2(n881), .ZN(n867) );
  NAND2_X1 U968 ( .A1(G118), .A2(n882), .ZN(n866) );
  NAND2_X1 U969 ( .A1(n867), .A2(n866), .ZN(n872) );
  NAND2_X1 U970 ( .A1(G142), .A2(n877), .ZN(n869) );
  NAND2_X1 U971 ( .A1(G106), .A2(n878), .ZN(n868) );
  NAND2_X1 U972 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U973 ( .A(n870), .B(KEYINPUT45), .Z(n871) );
  NOR2_X1 U974 ( .A1(n872), .A2(n871), .ZN(n874) );
  XNOR2_X1 U975 ( .A(n874), .B(n873), .ZN(n898) );
  XNOR2_X1 U976 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n876) );
  XNOR2_X1 U977 ( .A(n993), .B(KEYINPUT116), .ZN(n875) );
  XNOR2_X1 U978 ( .A(n876), .B(n875), .ZN(n893) );
  NAND2_X1 U979 ( .A1(G139), .A2(n877), .ZN(n880) );
  NAND2_X1 U980 ( .A1(G103), .A2(n878), .ZN(n879) );
  NAND2_X1 U981 ( .A1(n880), .A2(n879), .ZN(n888) );
  NAND2_X1 U982 ( .A1(G127), .A2(n881), .ZN(n884) );
  NAND2_X1 U983 ( .A1(G115), .A2(n882), .ZN(n883) );
  NAND2_X1 U984 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U985 ( .A(KEYINPUT47), .B(n885), .ZN(n886) );
  XNOR2_X1 U986 ( .A(KEYINPUT117), .B(n886), .ZN(n887) );
  NOR2_X1 U987 ( .A1(n888), .A2(n887), .ZN(n999) );
  XNOR2_X1 U988 ( .A(n889), .B(n999), .ZN(n891) );
  XNOR2_X1 U989 ( .A(G164), .B(G160), .ZN(n890) );
  XNOR2_X1 U990 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U991 ( .A(n893), .B(n892), .ZN(n896) );
  XNOR2_X1 U992 ( .A(n894), .B(G162), .ZN(n895) );
  XNOR2_X1 U993 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U994 ( .A(n898), .B(n897), .Z(n899) );
  NOR2_X1 U995 ( .A1(G37), .A2(n899), .ZN(G395) );
  XNOR2_X1 U996 ( .A(n913), .B(n900), .ZN(n902) );
  XNOR2_X1 U997 ( .A(G171), .B(n928), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U999 ( .A(n903), .B(G286), .Z(n904) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n904), .ZN(G397) );
  NOR2_X1 U1001 ( .A1(G229), .A2(G227), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(KEYINPUT49), .B(n905), .ZN(n906) );
  NOR2_X1 U1003 ( .A1(G401), .A2(n906), .ZN(n907) );
  AND2_X1 U1004 ( .A1(G319), .A2(n907), .ZN(n909) );
  NOR2_X1 U1005 ( .A1(G395), .A2(G397), .ZN(n908) );
  NAND2_X1 U1006 ( .A1(n909), .A2(n908), .ZN(G225) );
  INV_X1 U1007 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1008 ( .A(G1966), .B(G168), .Z(n910) );
  NOR2_X1 U1009 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1010 ( .A(KEYINPUT57), .B(n912), .ZN(n933) );
  XNOR2_X1 U1011 ( .A(G301), .B(G1961), .ZN(n915) );
  XNOR2_X1 U1012 ( .A(n913), .B(G1341), .ZN(n914) );
  NOR2_X1 U1013 ( .A1(n915), .A2(n914), .ZN(n927) );
  XNOR2_X1 U1014 ( .A(G1956), .B(n916), .ZN(n918) );
  NAND2_X1 U1015 ( .A1(G1971), .A2(G303), .ZN(n917) );
  NAND2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n919) );
  NOR2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1018 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1019 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1020 ( .A(n925), .B(KEYINPUT122), .ZN(n926) );
  NAND2_X1 U1021 ( .A1(n927), .A2(n926), .ZN(n930) );
  XOR2_X1 U1022 ( .A(G1348), .B(n928), .Z(n929) );
  NOR2_X1 U1023 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1024 ( .A(KEYINPUT123), .B(n931), .ZN(n932) );
  NOR2_X1 U1025 ( .A1(n933), .A2(n932), .ZN(n935) );
  XOR2_X1 U1026 ( .A(KEYINPUT56), .B(G16), .Z(n934) );
  NOR2_X1 U1027 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1028 ( .A(KEYINPUT124), .B(n936), .Z(n986) );
  XNOR2_X1 U1029 ( .A(G20), .B(n937), .ZN(n941) );
  XNOR2_X1 U1030 ( .A(G1981), .B(G6), .ZN(n939) );
  XNOR2_X1 U1031 ( .A(G1341), .B(G19), .ZN(n938) );
  NOR2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1033 ( .A1(n941), .A2(n940), .ZN(n944) );
  XOR2_X1 U1034 ( .A(KEYINPUT59), .B(G1348), .Z(n942) );
  XNOR2_X1 U1035 ( .A(G4), .B(n942), .ZN(n943) );
  NOR2_X1 U1036 ( .A1(n944), .A2(n943), .ZN(n946) );
  XOR2_X1 U1037 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n945) );
  XNOR2_X1 U1038 ( .A(n946), .B(n945), .ZN(n950) );
  XNOR2_X1 U1039 ( .A(G1966), .B(G21), .ZN(n948) );
  XNOR2_X1 U1040 ( .A(G1961), .B(G5), .ZN(n947) );
  NOR2_X1 U1041 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1042 ( .A1(n950), .A2(n949), .ZN(n958) );
  XNOR2_X1 U1043 ( .A(G1986), .B(G24), .ZN(n952) );
  XNOR2_X1 U1044 ( .A(G1971), .B(G22), .ZN(n951) );
  NOR2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n955) );
  XOR2_X1 U1046 ( .A(G1976), .B(KEYINPUT126), .Z(n953) );
  XNOR2_X1 U1047 ( .A(G23), .B(n953), .ZN(n954) );
  NAND2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(KEYINPUT58), .B(n956), .ZN(n957) );
  NOR2_X1 U1050 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1051 ( .A(KEYINPUT61), .B(n959), .Z(n960) );
  NOR2_X1 U1052 ( .A1(G16), .A2(n960), .ZN(n984) );
  XNOR2_X1 U1053 ( .A(G2084), .B(G34), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(n961), .B(KEYINPUT54), .ZN(n978) );
  XNOR2_X1 U1055 ( .A(G2090), .B(G35), .ZN(n975) );
  XNOR2_X1 U1056 ( .A(G1996), .B(G32), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(G33), .B(G2072), .ZN(n962) );
  NOR2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n969) );
  XOR2_X1 U1059 ( .A(G2067), .B(G26), .Z(n964) );
  NAND2_X1 U1060 ( .A1(n964), .A2(G28), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(G25), .B(n965), .ZN(n966) );
  NOR2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n972) );
  XOR2_X1 U1064 ( .A(G27), .B(n970), .Z(n971) );
  NOR2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1066 ( .A(KEYINPUT53), .B(n973), .ZN(n974) );
  NOR2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1068 ( .A(KEYINPUT120), .B(n976), .Z(n977) );
  NOR2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1070 ( .A(n979), .B(KEYINPUT55), .ZN(n981) );
  XNOR2_X1 U1071 ( .A(G29), .B(KEYINPUT121), .ZN(n980) );
  NAND2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1073 ( .A1(G11), .A2(n982), .ZN(n983) );
  NOR2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1076 ( .A(n987), .B(KEYINPUT127), .ZN(n1016) );
  INV_X1 U1077 ( .A(n988), .ZN(n989) );
  NOR2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n998) );
  XOR2_X1 U1079 ( .A(G2084), .B(G160), .Z(n991) );
  NOR2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n994) );
  NAND2_X1 U1081 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1082 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1083 ( .A1(n998), .A2(n997), .ZN(n1010) );
  XOR2_X1 U1084 ( .A(G2072), .B(n999), .Z(n1001) );
  XOR2_X1 U1085 ( .A(G164), .B(G2078), .Z(n1000) );
  NOR2_X1 U1086 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1087 ( .A(KEYINPUT50), .B(n1002), .ZN(n1008) );
  XOR2_X1 U1088 ( .A(G2090), .B(G162), .Z(n1003) );
  NOR2_X1 U1089 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1090 ( .A(KEYINPUT51), .B(n1005), .Z(n1006) );
  XNOR2_X1 U1091 ( .A(KEYINPUT118), .B(n1006), .ZN(n1007) );
  NAND2_X1 U1092 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1093 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1094 ( .A(KEYINPUT52), .B(n1011), .Z(n1012) );
  NOR2_X1 U1095 ( .A1(KEYINPUT55), .A2(n1012), .ZN(n1013) );
  XNOR2_X1 U1096 ( .A(KEYINPUT119), .B(n1013), .ZN(n1014) );
  NAND2_X1 U1097 ( .A1(n1014), .A2(G29), .ZN(n1015) );
  NAND2_X1 U1098 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1099 ( .A(KEYINPUT62), .B(n1017), .Z(G311) );
  INV_X1 U1100 ( .A(G311), .ZN(G150) );
endmodule

