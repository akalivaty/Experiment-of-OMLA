//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 1 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 1 1 1 0 1 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT27), .B(G183gat), .ZN(new_n203));
  INV_X1    g002(.A(G190gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NOR2_X1   g004(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n205), .B(new_n206), .Z(new_n207));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT69), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  AOI22_X1  g009(.A1(new_n210), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n211));
  AND2_X1   g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n212), .A2(KEYINPUT26), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n211), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n207), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G169gat), .ZN(new_n216));
  INV_X1    g015(.A(G176gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AND2_X1   g017(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n219));
  NOR2_X1   g018(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n212), .B1(KEYINPUT23), .B2(new_n208), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n218), .B(new_n224), .C1(new_n219), .C2(new_n220), .ZN(new_n225));
  AND3_X1   g024(.A1(new_n222), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT67), .ZN(new_n227));
  AND3_X1   g026(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230));
  NOR3_X1   g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n226), .A2(new_n227), .A3(KEYINPUT25), .A4(new_n232), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n222), .A2(KEYINPUT25), .A3(new_n223), .A4(new_n225), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT67), .B1(new_n234), .B2(new_n231), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT25), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n222), .A2(new_n223), .A3(new_n225), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT66), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n222), .A2(new_n241), .A3(new_n223), .A4(new_n225), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(new_n232), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n237), .B1(new_n240), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n215), .B1(new_n236), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n202), .B1(new_n245), .B2(KEYINPUT29), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT74), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n247), .B1(new_n245), .B2(new_n202), .ZN(new_n248));
  XNOR2_X1  g047(.A(G197gat), .B(G204gat), .ZN(new_n249));
  INV_X1    g048(.A(G211gat), .ZN(new_n250));
  INV_X1    g049(.A(G218gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n249), .B1(KEYINPUT22), .B2(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(G211gat), .B(G218gat), .Z(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  OR2_X1    g054(.A1(new_n207), .A2(new_n214), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n242), .A2(new_n232), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT25), .B1(new_n257), .B2(new_n239), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n233), .A2(new_n235), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n256), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n202), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(KEYINPUT74), .A3(new_n261), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n246), .A2(new_n248), .A3(new_n255), .A4(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT75), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n246), .B1(new_n202), .B2(new_n245), .ZN(new_n266));
  INV_X1    g065(.A(new_n255), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT76), .B(G64gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(G92gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(G8gat), .B(G36gat), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n270), .B(new_n271), .Z(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n265), .A2(KEYINPUT30), .A3(new_n268), .A4(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n262), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT74), .B1(new_n260), .B2(new_n261), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n277), .A2(new_n264), .A3(new_n255), .A4(new_n246), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT75), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(new_n279), .A3(new_n268), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(new_n272), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n278), .A2(new_n279), .A3(new_n268), .A4(new_n273), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT30), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n274), .A2(new_n281), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n286));
  INV_X1    g085(.A(G120gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(G113gat), .ZN(new_n288));
  INV_X1    g087(.A(G113gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G120gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G127gat), .B(G134gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT1), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n292), .B1(new_n293), .B2(new_n291), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n286), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n291), .A2(new_n293), .ZN(new_n297));
  INV_X1    g096(.A(new_n292), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(KEYINPUT70), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n296), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G148gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G141gat), .ZN(new_n304));
  INV_X1    g103(.A(G141gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G148gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G155gat), .ZN(new_n308));
  INV_X1    g107(.A(G162gat), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT2), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT77), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n305), .A2(G148gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n303), .A2(G141gat), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G155gat), .B(G162gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n311), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n307), .B(new_n310), .C1(new_n316), .C2(new_n312), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT4), .B1(new_n302), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT3), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n318), .A2(new_n322), .A3(new_n319), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT78), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT78), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n318), .A2(new_n325), .A3(new_n322), .A4(new_n319), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n318), .A2(new_n319), .ZN(new_n327));
  AOI22_X1  g126(.A1(new_n324), .A2(new_n326), .B1(KEYINPUT3), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n299), .A2(new_n300), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n321), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n320), .A2(KEYINPUT80), .A3(new_n300), .A4(new_n299), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT80), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n332), .B1(new_n327), .B2(new_n329), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(KEYINPUT4), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G225gat), .A2(G233gat), .ZN(new_n336));
  XOR2_X1   g135(.A(new_n336), .B(KEYINPUT79), .Z(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  OR2_X1    g137(.A1(new_n338), .A2(KEYINPUT39), .ZN(new_n339));
  XNOR2_X1  g138(.A(G1gat), .B(G29gat), .ZN(new_n340));
  INV_X1    g139(.A(G85gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT0), .B(G57gat), .ZN(new_n343));
  XOR2_X1   g142(.A(new_n342), .B(new_n343), .Z(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n331), .A2(new_n333), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n327), .A2(new_n329), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT81), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n327), .A2(KEYINPUT81), .A3(new_n329), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n337), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n346), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n338), .A2(new_n353), .A3(KEYINPUT39), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n339), .A2(new_n345), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT40), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n324), .A2(new_n326), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n327), .A2(KEYINPUT3), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n358), .A2(new_n329), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT4), .ZN(new_n361));
  AND2_X1   g160(.A1(new_n296), .A2(new_n301), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n361), .B1(new_n362), .B2(new_n327), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n337), .A2(KEYINPUT5), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n360), .A2(new_n334), .A3(new_n363), .A4(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT82), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT82), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n330), .A2(new_n367), .A3(new_n334), .A4(new_n364), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n349), .A2(new_n337), .A3(new_n350), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n352), .A2(KEYINPUT4), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n370), .A2(new_n346), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n327), .B1(new_n296), .B2(new_n301), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT4), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n337), .B1(new_n360), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT5), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n369), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(new_n344), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n339), .A2(KEYINPUT40), .A3(new_n345), .A4(new_n354), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n357), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n285), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT29), .B1(new_n324), .B2(new_n326), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT29), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT3), .B1(new_n255), .B2(new_n384), .ZN(new_n385));
  OAI22_X1  g184(.A1(new_n383), .A2(new_n255), .B1(new_n320), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT85), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(G22gat), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n388), .A2(G22gat), .ZN(new_n391));
  OAI211_X1 g190(.A(G228gat), .B(G233gat), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  OR2_X1    g191(.A1(new_n388), .A2(G22gat), .ZN(new_n393));
  INV_X1    g192(.A(G228gat), .ZN(new_n394));
  INV_X1    g193(.A(G233gat), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n393), .B(new_n389), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(G78gat), .B(G106gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT31), .B(G50gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n397), .B(new_n398), .ZN(new_n399));
  XOR2_X1   g198(.A(new_n399), .B(KEYINPUT86), .Z(new_n400));
  AND3_X1   g199(.A1(new_n392), .A2(new_n396), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(KEYINPUT86), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n402), .B1(new_n392), .B2(new_n396), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT87), .B(KEYINPUT38), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT37), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n280), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n278), .A2(new_n279), .A3(KEYINPUT37), .A4(new_n268), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n405), .B1(new_n409), .B2(new_n272), .ZN(new_n410));
  XOR2_X1   g209(.A(KEYINPUT83), .B(KEYINPUT6), .Z(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n369), .A2(new_n345), .A3(new_n377), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n379), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n378), .A2(new_n344), .A3(new_n411), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n282), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n246), .A2(new_n248), .A3(new_n262), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n267), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n246), .B(new_n255), .C1(new_n202), .C2(new_n245), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n418), .A2(KEYINPUT37), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n420), .B1(new_n406), .B2(new_n280), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n272), .A2(new_n405), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n416), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n382), .B(new_n404), .C1(new_n410), .C2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  OR2_X1    g224(.A1(new_n401), .A2(new_n403), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n411), .B1(new_n378), .B2(new_n344), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT84), .B1(new_n427), .B2(new_n413), .ZN(new_n428));
  AOI22_X1  g227(.A1(new_n328), .A2(new_n329), .B1(KEYINPUT4), .B2(new_n374), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n372), .B1(new_n429), .B2(new_n337), .ZN(new_n430));
  AOI22_X1  g229(.A1(new_n366), .A2(new_n368), .B1(new_n430), .B2(KEYINPUT5), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n412), .B1(new_n431), .B2(new_n345), .ZN(new_n432));
  INV_X1    g231(.A(new_n413), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n415), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n428), .B1(KEYINPUT84), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n426), .B1(new_n285), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT36), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT34), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n260), .A2(new_n362), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n302), .B(new_n256), .C1(new_n258), .C2(new_n259), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G227gat), .A2(G233gat), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n438), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n439), .A2(KEYINPUT34), .A3(new_n442), .A4(new_n440), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT73), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT71), .ZN(new_n449));
  XNOR2_X1  g248(.A(G15gat), .B(G43gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(G71gat), .B(G99gat), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n450), .B(new_n451), .Z(new_n452));
  AOI21_X1  g251(.A(new_n442), .B1(new_n439), .B2(new_n440), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n452), .B1(new_n453), .B2(KEYINPUT33), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT32), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n455), .B1(new_n441), .B2(new_n443), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n449), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n244), .A2(new_n235), .A3(new_n233), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n302), .B1(new_n458), .B2(new_n256), .ZN(new_n459));
  INV_X1    g258(.A(new_n440), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n443), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT32), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT33), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n462), .A2(new_n464), .A3(KEYINPUT71), .A4(new_n452), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n457), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n444), .A2(KEYINPUT73), .A3(new_n445), .ZN(new_n467));
  INV_X1    g266(.A(new_n452), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n463), .B1(new_n468), .B2(KEYINPUT72), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n469), .B1(KEYINPUT72), .B2(new_n468), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n456), .A2(new_n470), .ZN(new_n471));
  AND4_X1   g270(.A1(new_n448), .A2(new_n466), .A3(new_n467), .A4(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n471), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n473), .B1(new_n457), .B2(new_n465), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n448), .B1(new_n474), .B2(new_n467), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n437), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n468), .B1(new_n461), .B2(new_n463), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT71), .B1(new_n477), .B2(new_n462), .ZN(new_n478));
  NOR3_X1   g277(.A1(new_n454), .A2(new_n449), .A3(new_n456), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n471), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n480), .A2(new_n447), .A3(new_n446), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n474), .A2(new_n448), .A3(new_n467), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(KEYINPUT36), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n436), .A2(new_n476), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n285), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n481), .A2(new_n482), .ZN(new_n486));
  AOI211_X1 g285(.A(new_n345), .B(new_n412), .C1(new_n369), .C2(new_n377), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n487), .B1(new_n427), .B2(new_n413), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n488), .A2(KEYINPUT35), .ZN(new_n489));
  AND4_X1   g288(.A1(new_n485), .A2(new_n486), .A3(new_n404), .A4(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT35), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n426), .B1(new_n481), .B2(new_n482), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n285), .A2(new_n435), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI22_X1  g293(.A1(new_n425), .A2(new_n484), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  XOR2_X1   g294(.A(G15gat), .B(G22gat), .Z(new_n496));
  INV_X1    g295(.A(G1gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(G8gat), .B1(new_n498), .B2(KEYINPUT90), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n497), .A2(KEYINPUT16), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n498), .B1(new_n500), .B2(new_n496), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n499), .B(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT21), .ZN(new_n503));
  NAND2_X1  g302(.A1(G71gat), .A2(G78gat), .ZN(new_n504));
  OR2_X1    g303(.A1(G71gat), .A2(G78gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(G57gat), .B(G64gat), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT9), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n504), .B(new_n505), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  OR2_X1    g307(.A1(new_n508), .A2(KEYINPUT93), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n505), .A2(new_n507), .ZN(new_n510));
  INV_X1    g309(.A(new_n504), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OR2_X1    g311(.A1(new_n512), .A2(new_n506), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n508), .A2(KEYINPUT93), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n509), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n502), .B1(new_n503), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(G183gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n515), .A2(new_n503), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(G211gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n519), .B(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G127gat), .B(G155gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(G231gat), .A2(G233gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n522), .A2(new_n526), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OR3_X1    g328(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n531));
  AOI22_X1  g330(.A1(new_n530), .A2(new_n531), .B1(G29gat), .B2(G36gat), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT15), .ZN(new_n533));
  XOR2_X1   g332(.A(G43gat), .B(G50gat), .Z(new_n534));
  OR3_X1    g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n534), .A2(new_n533), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n533), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n536), .A2(new_n537), .A3(new_n532), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(KEYINPUT89), .A2(KEYINPUT17), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(KEYINPUT89), .A2(KEYINPUT17), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(G85gat), .A2(G92gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT7), .ZN(new_n545));
  INV_X1    g344(.A(G99gat), .ZN(new_n546));
  INV_X1    g345(.A(G106gat), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT8), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n545), .B(new_n548), .C1(G85gat), .C2(G92gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT94), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(G99gat), .B(G106gat), .Z(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OR2_X1    g352(.A1(new_n551), .A2(new_n552), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n543), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n553), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n539), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G190gat), .B(G218gat), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(G134gat), .B(G162gat), .Z(new_n562));
  AOI21_X1  g361(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT95), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n559), .A2(new_n560), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(new_n565), .ZN(new_n568));
  INV_X1    g367(.A(new_n564), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n568), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n566), .B1(new_n570), .B2(new_n561), .ZN(new_n571));
  NAND2_X1  g370(.A1(G230gat), .A2(G233gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n515), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT10), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n554), .A2(new_n515), .A3(new_n553), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n557), .A2(KEYINPUT10), .A3(new_n574), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n573), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n575), .A2(new_n577), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n580), .B1(new_n581), .B2(new_n573), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT96), .B(G176gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(G204gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(G120gat), .B(G148gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n584), .B(new_n585), .Z(new_n586));
  OR2_X1    g385(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n578), .A2(new_n579), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(new_n572), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n581), .A2(new_n573), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n589), .A2(new_n590), .A3(new_n586), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n529), .A2(new_n571), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n539), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n502), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n596), .B1(new_n543), .B2(new_n502), .ZN(new_n597));
  NAND2_X1  g396(.A1(G229gat), .A2(G233gat), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OR2_X1    g398(.A1(new_n599), .A2(KEYINPUT18), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n502), .A2(new_n595), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT92), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n502), .A2(new_n595), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(new_n598), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n599), .A2(KEYINPUT18), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n600), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G169gat), .B(G197gat), .Z(new_n611));
  XNOR2_X1  g410(.A(G113gat), .B(G141gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n615), .B(KEYINPUT12), .Z(new_n616));
  NAND2_X1  g415(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n616), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n600), .A2(new_n608), .A3(new_n609), .A4(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n594), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n495), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT84), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n414), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n625), .B1(new_n488), .B2(new_n624), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT97), .B(G1gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(G1324gat));
  INV_X1    g428(.A(new_n623), .ZN(new_n630));
  XOR2_X1   g429(.A(KEYINPUT16), .B(G8gat), .Z(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(new_n285), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT42), .ZN(new_n633));
  OAI21_X1  g432(.A(G8gat), .B1(new_n623), .B2(new_n485), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(G1325gat));
  NAND2_X1  g434(.A1(new_n476), .A2(new_n483), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n637), .A2(KEYINPUT98), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(KEYINPUT98), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n630), .A2(G15gat), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n486), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n623), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n641), .B1(G15gat), .B2(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n644), .B(KEYINPUT99), .Z(G1326gat));
  NOR2_X1   g444(.A1(new_n623), .A2(new_n404), .ZN(new_n646));
  XOR2_X1   g445(.A(KEYINPUT43), .B(G22gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(G1327gat));
  AND3_X1   g447(.A1(new_n436), .A2(new_n476), .A3(new_n483), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n404), .B1(new_n472), .B2(new_n475), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n626), .A2(new_n281), .A3(new_n274), .A4(new_n284), .ZN(new_n651));
  OAI21_X1  g450(.A(KEYINPUT35), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n492), .A2(new_n485), .A3(new_n489), .ZN(new_n653));
  AOI22_X1  g452(.A1(new_n649), .A2(new_n424), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(new_n571), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n527), .A2(new_n528), .ZN(new_n656));
  AND4_X1   g455(.A1(new_n620), .A2(new_n655), .A3(new_n656), .A4(new_n593), .ZN(new_n657));
  INV_X1    g456(.A(G29gat), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(new_n658), .A3(new_n435), .ZN(new_n659));
  XNOR2_X1  g458(.A(KEYINPUT100), .B(KEYINPUT45), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT44), .B1(new_n654), .B2(new_n571), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663));
  INV_X1    g462(.A(new_n571), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n495), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n592), .B(KEYINPUT101), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n667), .A2(new_n620), .A3(new_n656), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n658), .B1(new_n671), .B2(new_n435), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n661), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT102), .ZN(G1328gat));
  INV_X1    g473(.A(G36gat), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n657), .A2(new_n675), .A3(new_n285), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n676), .B(KEYINPUT46), .Z(new_n677));
  OAI21_X1  g476(.A(G36gat), .B1(new_n670), .B2(new_n485), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(G1329gat));
  OAI21_X1  g478(.A(G43gat), .B1(new_n670), .B2(new_n637), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n642), .A2(G43gat), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n657), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n680), .A2(KEYINPUT47), .A3(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n640), .ZN(new_n684));
  OAI21_X1  g483(.A(G43gat), .B1(new_n670), .B2(new_n684), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n685), .A2(new_n682), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT103), .B(KEYINPUT47), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n683), .B1(new_n686), .B2(new_n687), .ZN(G1330gat));
  INV_X1    g487(.A(G50gat), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n657), .A2(new_n689), .A3(new_n426), .ZN(new_n690));
  AOI211_X1 g489(.A(new_n404), .B(new_n668), .C1(new_n662), .C2(new_n665), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n690), .B(KEYINPUT48), .C1(new_n689), .C2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT105), .B1(new_n691), .B2(new_n689), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n666), .A2(new_n426), .A3(new_n669), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(new_n695), .A3(G50gat), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n693), .A2(new_n690), .A3(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT106), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT104), .B(KEYINPUT48), .Z(new_n699));
  AND3_X1   g498(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n698), .B1(new_n697), .B2(new_n699), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n692), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI211_X1 g503(.A(KEYINPUT107), .B(new_n692), .C1(new_n700), .C2(new_n701), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(G1331gat));
  NOR2_X1   g505(.A1(new_n656), .A2(new_n664), .ZN(new_n707));
  INV_X1    g506(.A(new_n667), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n495), .A2(new_n621), .A3(new_n707), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT108), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n435), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g511(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n710), .A2(new_n285), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT109), .ZN(new_n715));
  NOR2_X1   g514(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1333gat));
  AOI21_X1  g516(.A(G71gat), .B1(new_n710), .B2(new_n486), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n640), .A2(G71gat), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n718), .B1(new_n710), .B2(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g520(.A1(new_n710), .A2(new_n426), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT110), .B(G78gat), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1335gat));
  AOI21_X1  g523(.A(new_n593), .B1(new_n662), .B2(new_n665), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n529), .A2(new_n620), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(KEYINPUT111), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n729), .B1(new_n725), .B2(new_n726), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(G85gat), .B1(new_n731), .B2(new_n626), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n655), .A2(KEYINPUT51), .A3(new_n726), .ZN(new_n733));
  AOI21_X1  g532(.A(KEYINPUT51), .B1(new_n655), .B2(new_n726), .ZN(new_n734));
  OR2_X1    g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n592), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n435), .A2(new_n341), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n732), .B1(new_n736), .B2(new_n737), .ZN(G1336gat));
  OR3_X1    g537(.A1(new_n727), .A2(KEYINPUT112), .A3(new_n485), .ZN(new_n739));
  OAI21_X1  g538(.A(KEYINPUT112), .B1(new_n727), .B2(new_n485), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n739), .A2(G92gat), .A3(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT52), .ZN(new_n742));
  INV_X1    g541(.A(G92gat), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n735), .A2(new_n743), .A3(new_n285), .A4(new_n708), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(G92gat), .B1(new_n731), .B2(new_n485), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n746), .A2(new_n744), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n747), .B2(new_n742), .ZN(G1337gat));
  OAI21_X1  g547(.A(G99gat), .B1(new_n731), .B2(new_n684), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n486), .A2(new_n546), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n736), .B2(new_n750), .ZN(G1338gat));
  OAI21_X1  g550(.A(G106gat), .B1(new_n727), .B2(new_n404), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT53), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n547), .B(new_n708), .C1(new_n733), .C2(new_n734), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n752), .B(new_n753), .C1(new_n754), .C2(new_n404), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n754), .A2(new_n404), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n426), .B1(new_n728), .B2(new_n730), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n756), .B1(new_n757), .B2(G106gat), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n755), .B1(new_n758), .B2(new_n753), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT113), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OAI211_X1 g560(.A(KEYINPUT113), .B(new_n755), .C1(new_n758), .C2(new_n753), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(G1339gat));
  NAND3_X1  g562(.A1(new_n578), .A2(new_n579), .A3(new_n573), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n589), .A2(KEYINPUT54), .A3(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT54), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n586), .B1(new_n580), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT55), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n605), .A2(new_n607), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n597), .A2(new_n598), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n615), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n619), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n765), .A2(KEYINPUT55), .A3(new_n767), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n775), .A2(new_n591), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n770), .A2(new_n664), .A3(new_n774), .A4(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n770), .A2(new_n620), .A3(new_n776), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n592), .A2(new_n774), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n777), .B1(new_n780), .B2(new_n664), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n656), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n594), .A2(new_n620), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n285), .A2(new_n626), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n787), .A2(new_n492), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n620), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(G113gat), .ZN(G1340gat));
  NAND3_X1  g589(.A1(new_n788), .A2(new_n287), .A3(new_n592), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n788), .A2(new_n708), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n792), .A2(KEYINPUT115), .A3(G120gat), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT115), .B1(new_n792), .B2(G120gat), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n791), .B1(new_n793), .B2(new_n794), .ZN(G1341gat));
  NAND2_X1  g594(.A1(new_n788), .A2(new_n529), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g596(.A1(new_n788), .A2(new_n664), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT56), .ZN(new_n799));
  INV_X1    g598(.A(G134gat), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT116), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n798), .A2(KEYINPUT56), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n799), .A2(new_n804), .A3(new_n800), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n802), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n804), .B1(new_n799), .B2(new_n800), .ZN(new_n807));
  AOI211_X1 g606(.A(KEYINPUT116), .B(G134gat), .C1(new_n798), .C2(KEYINPUT56), .ZN(new_n808));
  OAI22_X1  g607(.A1(new_n807), .A2(new_n808), .B1(KEYINPUT56), .B2(new_n798), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n806), .A2(new_n809), .ZN(G1343gat));
  INV_X1    g609(.A(KEYINPUT58), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n404), .B1(new_n782), .B2(new_n784), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n636), .A2(new_n626), .A3(new_n285), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n765), .A2(new_n767), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n620), .A2(new_n776), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n664), .B1(new_n819), .B2(new_n779), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n820), .A2(KEYINPUT117), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n777), .B1(new_n820), .B2(KEYINPUT117), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n656), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n404), .B1(new_n823), .B2(new_n784), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n814), .B(new_n815), .C1(new_n824), .C2(new_n813), .ZN(new_n825));
  OAI21_X1  g624(.A(G141gat), .B1(new_n825), .B2(new_n621), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n811), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n812), .A2(new_n684), .A3(new_n786), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n621), .A2(G141gat), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n826), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n828), .B(new_n832), .ZN(G1344gat));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n769), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n768), .A2(KEYINPUT114), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n834), .A2(new_n664), .A3(new_n776), .A4(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT121), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n770), .A2(KEYINPUT121), .A3(new_n664), .A4(new_n776), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n838), .A2(new_n839), .A3(new_n774), .ZN(new_n840));
  INV_X1    g639(.A(new_n820), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n529), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n707), .A2(KEYINPUT120), .A3(new_n621), .A4(new_n593), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT120), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n844), .B1(new_n594), .B2(new_n620), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n426), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n813), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT122), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n812), .A2(KEYINPUT57), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n847), .A2(KEYINPUT122), .A3(new_n813), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(new_n592), .A3(new_n815), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT123), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n853), .A2(KEYINPUT123), .A3(new_n592), .A4(new_n815), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n856), .A2(G148gat), .A3(new_n857), .ZN(new_n858));
  XNOR2_X1  g657(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n861), .B(G148gat), .C1(new_n825), .C2(new_n593), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  OR3_X1    g662(.A1(new_n829), .A2(G148gat), .A3(new_n593), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(G1345gat));
  NOR3_X1   g664(.A1(new_n825), .A2(new_n308), .A3(new_n656), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n829), .A2(new_n656), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n866), .B1(new_n308), .B2(new_n867), .ZN(G1346gat));
  NOR3_X1   g667(.A1(new_n825), .A2(new_n309), .A3(new_n571), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n829), .A2(new_n571), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n869), .B1(new_n309), .B2(new_n870), .ZN(G1347gat));
  NOR2_X1   g670(.A1(new_n485), .A2(new_n435), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  AOI211_X1 g672(.A(new_n650), .B(new_n873), .C1(new_n782), .C2(new_n784), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n620), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(G169gat), .ZN(G1348gat));
  AOI21_X1  g675(.A(G176gat), .B1(new_n874), .B2(new_n592), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n874), .A2(G176gat), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n708), .B2(new_n878), .ZN(G1349gat));
  NAND2_X1  g678(.A1(new_n874), .A2(new_n529), .ZN(new_n880));
  MUX2_X1   g679(.A(new_n203), .B(G183gat), .S(new_n880), .Z(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g681(.A1(new_n874), .A2(new_n664), .ZN(new_n883));
  NAND2_X1  g682(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n883), .A2(G190gat), .A3(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n886));
  XOR2_X1   g685(.A(new_n885), .B(new_n886), .Z(new_n887));
  OAI21_X1  g686(.A(new_n887), .B1(G190gat), .B2(new_n883), .ZN(G1351gat));
  NOR2_X1   g687(.A1(new_n640), .A2(new_n873), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n853), .A2(new_n620), .A3(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT126), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(G197gat), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n812), .A2(new_n889), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT125), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n895), .B(new_n896), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n621), .A2(G197gat), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(G1352gat));
  NOR3_X1   g698(.A1(new_n895), .A2(G204gat), .A3(new_n593), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT62), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n853), .A2(new_n889), .ZN(new_n902));
  OAI21_X1  g701(.A(G204gat), .B1(new_n902), .B2(new_n667), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(G1353gat));
  NAND3_X1  g703(.A1(new_n853), .A2(new_n529), .A3(new_n889), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n905), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT63), .B1(new_n905), .B2(G211gat), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n529), .A2(new_n250), .ZN(new_n908));
  OAI22_X1  g707(.A1(new_n906), .A2(new_n907), .B1(new_n897), .B2(new_n908), .ZN(G1354gat));
  NOR3_X1   g708(.A1(new_n902), .A2(new_n251), .A3(new_n571), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n251), .B1(new_n897), .B2(new_n571), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n911), .A2(KEYINPUT127), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(KEYINPUT127), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(G1355gat));
endmodule


