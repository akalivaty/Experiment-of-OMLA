//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087, new_n1088, new_n1089, new_n1090, new_n1091,
    new_n1092, new_n1093, new_n1094;
  XNOR2_X1  g000(.A(G110), .B(G122), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OR2_X1    g002(.A1(KEYINPUT71), .A2(G119), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT5), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT71), .A2(G119), .ZN(new_n191));
  NAND4_X1  g005(.A1(new_n189), .A2(new_n190), .A3(G116), .A4(new_n191), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n192), .A2(G113), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n189), .A2(G116), .A3(new_n191), .ZN(new_n194));
  INV_X1    g008(.A(G116), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G119), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(KEYINPUT5), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n196), .ZN(new_n198));
  AND2_X1   g012(.A1(KEYINPUT71), .A2(G119), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT71), .A2(G119), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n198), .B1(new_n201), .B2(G116), .ZN(new_n202));
  XOR2_X1   g016(.A(KEYINPUT2), .B(G113), .Z(new_n203));
  AOI22_X1  g017(.A1(new_n193), .A2(new_n197), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G101), .ZN(new_n205));
  INV_X1    g019(.A(G107), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G104), .ZN(new_n207));
  INV_X1    g021(.A(G104), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G107), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n205), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT3), .B1(new_n208), .B2(G107), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(new_n206), .A3(G104), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n211), .A2(new_n213), .A3(new_n209), .ZN(new_n214));
  AND2_X1   g028(.A1(KEYINPUT81), .A2(G101), .ZN(new_n215));
  NOR2_X1   g029(.A1(KEYINPUT81), .A2(G101), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n210), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(KEYINPUT84), .B1(new_n204), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n197), .A2(G113), .A3(new_n192), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n202), .A2(new_n203), .ZN(new_n221));
  AND4_X1   g035(.A1(KEYINPUT84), .A2(new_n220), .A3(new_n218), .A4(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n211), .A2(new_n213), .A3(new_n209), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT4), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(new_n225), .A3(G101), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n202), .A2(new_n203), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n203), .A2(new_n194), .A3(new_n196), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n225), .B1(new_n214), .B2(new_n217), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT82), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n224), .A2(G101), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n217), .A2(new_n211), .A3(new_n213), .A4(new_n209), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT4), .ZN(new_n235));
  INV_X1    g049(.A(new_n232), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT82), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n229), .B1(new_n233), .B2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n188), .B1(new_n223), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n227), .A2(new_n228), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n231), .B1(new_n230), .B2(new_n232), .ZN(new_n242));
  AND4_X1   g056(.A1(new_n231), .A2(new_n232), .A3(KEYINPUT4), .A4(new_n234), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n241), .B(new_n226), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT84), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n220), .A2(new_n221), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n207), .A2(new_n209), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G101), .ZN(new_n248));
  OR2_X1    g062(.A1(new_n215), .A2(new_n216), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n248), .B1(new_n224), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n245), .B1(new_n246), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n204), .A2(KEYINPUT84), .A3(new_n218), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n244), .A2(new_n253), .A3(new_n187), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n239), .A2(KEYINPUT6), .A3(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(G143), .B(G146), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT64), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XOR2_X1   g072(.A(KEYINPUT0), .B(G128), .Z(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI211_X1 g074(.A(KEYINPUT0), .B(G128), .C1(new_n256), .C2(new_n257), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G125), .ZN(new_n263));
  INV_X1    g077(.A(G143), .ZN(new_n264));
  INV_X1    g078(.A(G128), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n264), .B(G146), .C1(new_n265), .C2(KEYINPUT1), .ZN(new_n266));
  INV_X1    g080(.A(G146), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n265), .A2(new_n267), .A3(G143), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n266), .A2(KEYINPUT70), .A3(new_n268), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT69), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n265), .A2(KEYINPUT1), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n273), .B1(new_n256), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n267), .A2(G143), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n264), .A2(G146), .ZN(new_n277));
  AND4_X1   g091(.A1(new_n273), .A2(new_n274), .A3(new_n276), .A4(new_n277), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n271), .B(new_n272), .C1(new_n275), .C2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n263), .B1(G125), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G224), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n282), .A2(G953), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n283), .B(KEYINPUT85), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n281), .B(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT6), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n286), .B(new_n188), .C1(new_n223), .C2(new_n238), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n255), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT7), .B1(new_n282), .B2(G953), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n281), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n289), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n263), .B(new_n291), .C1(G125), .C2(new_n280), .ZN(new_n292));
  OR2_X1    g106(.A1(new_n250), .A2(KEYINPUT86), .ZN(new_n293));
  OR2_X1    g107(.A1(new_n293), .A2(new_n204), .ZN(new_n294));
  XOR2_X1   g108(.A(new_n187), .B(KEYINPUT8), .Z(new_n295));
  AOI21_X1  g109(.A(new_n295), .B1(new_n293), .B2(new_n204), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n290), .A2(new_n292), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(G902), .B1(new_n297), .B2(new_n254), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n288), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G210), .B1(G237), .B2(G902), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n288), .A2(new_n298), .A3(new_n300), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G214), .B1(G237), .B2(G902), .ZN(new_n305));
  INV_X1    g119(.A(G902), .ZN(new_n306));
  INV_X1    g120(.A(G237), .ZN(new_n307));
  INV_X1    g121(.A(G953), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n308), .A3(G214), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT87), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n309), .B1(new_n310), .B2(new_n264), .ZN(new_n311));
  NOR2_X1   g125(.A1(G237), .A2(G953), .ZN(new_n312));
  AND2_X1   g126(.A1(KEYINPUT87), .A2(G143), .ZN(new_n313));
  NOR2_X1   g127(.A1(KEYINPUT87), .A2(G143), .ZN(new_n314));
  OAI211_X1 g128(.A(G214), .B(new_n312), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  XOR2_X1   g130(.A(KEYINPUT66), .B(G131), .Z(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT17), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n311), .A2(new_n315), .A3(new_n317), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G140), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G125), .ZN(new_n324));
  INV_X1    g138(.A(G125), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G140), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT16), .ZN(new_n327));
  OR3_X1    g141(.A1(new_n325), .A2(KEYINPUT16), .A3(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n267), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n327), .A2(new_n328), .A3(G146), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n316), .A2(KEYINPUT17), .A3(new_n318), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n322), .A2(new_n330), .A3(new_n331), .A4(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(G113), .B(G122), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(new_n208), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT18), .ZN(new_n336));
  INV_X1    g150(.A(G131), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n316), .A2(new_n338), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n324), .A2(new_n326), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n267), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n324), .A2(new_n326), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G146), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n311), .B(new_n315), .C1(new_n336), .C2(new_n337), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n339), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(KEYINPUT88), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT88), .ZN(new_n348));
  AOI22_X1  g162(.A1(new_n316), .A2(new_n338), .B1(new_n341), .B2(new_n343), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n348), .B1(new_n349), .B2(new_n345), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n333), .B(new_n335), .C1(new_n347), .C2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n346), .A2(KEYINPUT88), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n349), .A2(new_n348), .A3(new_n345), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n335), .B1(new_n355), .B2(new_n333), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n306), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G475), .ZN(new_n358));
  INV_X1    g172(.A(new_n331), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n340), .B(KEYINPUT19), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n359), .B1(new_n360), .B2(new_n267), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n319), .A2(new_n321), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n353), .A2(new_n354), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n351), .B1(new_n363), .B2(new_n335), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT20), .ZN(new_n365));
  NOR2_X1   g179(.A1(G475), .A2(G902), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n365), .B1(new_n364), .B2(new_n366), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n358), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  XOR2_X1   g183(.A(G116), .B(G122), .Z(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G107), .ZN(new_n371));
  XNOR2_X1  g185(.A(G116), .B(G122), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n206), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT13), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(new_n264), .A3(G128), .ZN(new_n376));
  XOR2_X1   g190(.A(G128), .B(G143), .Z(new_n377));
  OAI211_X1 g191(.A(G134), .B(new_n376), .C1(new_n377), .C2(new_n375), .ZN(new_n378));
  XNOR2_X1  g192(.A(G128), .B(G143), .ZN(new_n379));
  INV_X1    g193(.A(G134), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT89), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT89), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n379), .A2(new_n383), .A3(new_n380), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n374), .A2(new_n378), .A3(new_n382), .A4(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n377), .A2(G134), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n381), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n195), .A2(KEYINPUT14), .A3(G122), .ZN(new_n388));
  OAI211_X1 g202(.A(G107), .B(new_n388), .C1(new_n370), .C2(KEYINPUT14), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n387), .A2(new_n389), .A3(new_n373), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT9), .B(G234), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(KEYINPUT80), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n308), .A2(G217), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n385), .A2(new_n390), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n394), .B1(new_n385), .B2(new_n390), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n306), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G478), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(KEYINPUT15), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n385), .A2(new_n390), .ZN(new_n401));
  INV_X1    g215(.A(new_n394), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n385), .A2(new_n394), .A3(new_n390), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n399), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n306), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n400), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT90), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G952), .ZN(new_n411));
  AOI211_X1 g225(.A(G953), .B(new_n411), .C1(G234), .C2(G237), .ZN(new_n412));
  AOI211_X1 g226(.A(new_n306), .B(new_n308), .C1(G234), .C2(G237), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT21), .B(G898), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n400), .A2(new_n407), .A3(KEYINPUT90), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n410), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n369), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n304), .A2(new_n305), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G469), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n260), .A2(new_n226), .A3(new_n261), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n423), .B1(new_n242), .B2(new_n243), .ZN(new_n424));
  INV_X1    g238(.A(new_n269), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n425), .B1(new_n275), .B2(new_n278), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT10), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n427), .A3(new_n218), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n266), .A2(KEYINPUT70), .A3(new_n268), .ZN(new_n429));
  AOI21_X1  g243(.A(KEYINPUT70), .B1(new_n266), .B2(new_n268), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n274), .A2(new_n276), .A3(new_n277), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT69), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n256), .A2(new_n273), .A3(new_n274), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n250), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n428), .B1(new_n436), .B2(new_n427), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT65), .B1(new_n380), .B2(G137), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT11), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT11), .ZN(new_n440));
  OAI211_X1 g254(.A(KEYINPUT65), .B(new_n440), .C1(new_n380), .C2(G137), .ZN(new_n441));
  INV_X1    g255(.A(G137), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(G134), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n439), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT67), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n446), .A3(G131), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n443), .B1(new_n438), .B2(KEYINPUT11), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(new_n441), .A3(new_n317), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n337), .B1(new_n448), .B2(new_n441), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n451), .A2(new_n446), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n424), .A2(new_n437), .A3(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G110), .B(G140), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n308), .A2(G227), .ZN(new_n456));
  XOR2_X1   g270(.A(new_n455), .B(new_n456), .Z(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n426), .A2(new_n218), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n431), .A2(new_n435), .A3(new_n250), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n439), .A2(new_n441), .A3(new_n444), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT67), .B1(new_n463), .B2(new_n337), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(new_n449), .A3(new_n447), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT12), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n462), .A2(new_n465), .A3(KEYINPUT12), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n466), .B1(KEYINPUT83), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT83), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n462), .A2(new_n465), .A3(new_n469), .A4(KEYINPUT12), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n459), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n427), .B1(new_n279), .B2(new_n218), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n269), .B1(new_n433), .B2(new_n434), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n473), .A2(KEYINPUT10), .A3(new_n250), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n422), .B1(new_n237), .B2(new_n233), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n465), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n458), .B1(new_n477), .B2(new_n454), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n421), .B(new_n306), .C1(new_n471), .C2(new_n478), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n454), .A2(new_n458), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n477), .ZN(new_n481));
  INV_X1    g295(.A(new_n454), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n482), .B1(new_n468), .B2(new_n470), .ZN(new_n483));
  OAI211_X1 g297(.A(G469), .B(new_n481), .C1(new_n483), .C2(new_n458), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n421), .A2(new_n306), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n479), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G221), .ZN(new_n488));
  INV_X1    g302(.A(new_n392), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n488), .B1(new_n489), .B2(new_n306), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n420), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G217), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n494), .B1(G234), .B2(new_n306), .ZN(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT22), .B(G137), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n308), .A2(G221), .A3(G234), .ZN(new_n497));
  XOR2_X1   g311(.A(new_n496), .B(new_n497), .Z(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT79), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n265), .A2(KEYINPUT23), .A3(G119), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n501), .B1(new_n201), .B2(G128), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n265), .B1(new_n199), .B2(new_n200), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT23), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(G110), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n502), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n189), .A2(G128), .A3(new_n191), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n265), .A2(G119), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n506), .A2(KEYINPUT24), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT24), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G110), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n510), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n507), .A2(new_n514), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n331), .A2(new_n341), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT78), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n189), .A2(new_n191), .ZN(new_n518));
  AOI21_X1  g332(.A(KEYINPUT23), .B1(new_n518), .B2(new_n265), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n265), .A2(KEYINPUT23), .A3(G119), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n508), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n517), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n502), .A2(new_n505), .A3(KEYINPUT78), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(G110), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n511), .A2(new_n513), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n508), .A2(new_n509), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT77), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT77), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n508), .A2(new_n525), .A3(new_n528), .A4(new_n509), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n527), .A2(new_n529), .B1(new_n330), .B2(new_n331), .ZN(new_n530));
  AOI221_X4 g344(.A(new_n500), .B1(new_n515), .B2(new_n516), .C1(new_n524), .C2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n524), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n515), .A2(new_n516), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT79), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n499), .B1(new_n531), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n532), .A2(new_n533), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n498), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT25), .B1(new_n538), .B2(new_n306), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT25), .ZN(new_n540));
  AOI211_X1 g354(.A(new_n540), .B(G902), .C1(new_n535), .C2(new_n537), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n495), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n495), .A2(G902), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  AND2_X1   g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(G472), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n262), .B1(new_n450), .B2(new_n452), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n442), .A2(KEYINPUT68), .A3(G134), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT68), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n380), .B2(G137), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n444), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(G131), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n279), .A2(new_n449), .A3(new_n552), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n547), .A2(new_n240), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n240), .B1(new_n547), .B2(new_n553), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT28), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT76), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n312), .A2(G210), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(KEYINPUT27), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT26), .B(G101), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n559), .B(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n547), .A2(new_n240), .A3(new_n553), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT28), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT76), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n566), .B(KEYINPUT28), .C1(new_n554), .C2(new_n555), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n557), .A2(KEYINPUT29), .A3(new_n565), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n306), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n260), .A2(new_n261), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n446), .A2(new_n451), .B1(new_n463), .B2(new_n317), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n570), .B1(new_n571), .B2(new_n464), .ZN(new_n572));
  INV_X1    g386(.A(new_n553), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT30), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT30), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n547), .A2(new_n575), .A3(new_n553), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n554), .B1(new_n577), .B2(new_n241), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT74), .B1(new_n578), .B2(new_n561), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n556), .A2(new_n565), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT29), .B1(new_n580), .B2(KEYINPUT73), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT74), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n240), .B1(new_n574), .B2(new_n576), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n582), .B(new_n562), .C1(new_n583), .C2(new_n554), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT73), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n556), .A2(new_n585), .A3(new_n565), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n579), .A2(new_n581), .A3(new_n584), .A4(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n569), .B1(new_n587), .B2(KEYINPUT75), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n241), .B1(new_n572), .B2(new_n573), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n564), .B1(new_n589), .B2(new_n563), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n563), .A2(new_n564), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n561), .ZN(new_n592));
  OAI21_X1  g406(.A(KEYINPUT73), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT29), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n593), .A2(new_n594), .A3(new_n586), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT75), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n595), .A2(new_n596), .A3(new_n584), .A4(new_n579), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n546), .B1(new_n588), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT31), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n563), .A2(new_n561), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n599), .B1(new_n583), .B2(new_n600), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n547), .A2(new_n575), .A3(new_n553), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n575), .B1(new_n547), .B2(new_n553), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n241), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n600), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(KEYINPUT31), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n556), .A2(new_n591), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n601), .A2(new_n606), .B1(new_n607), .B2(new_n562), .ZN(new_n608));
  NOR2_X1   g422(.A1(G472), .A2(G902), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT72), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n591), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n562), .B1(new_n590), .B2(new_n612), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n583), .A2(new_n599), .A3(new_n600), .ZN(new_n614));
  AOI21_X1  g428(.A(KEYINPUT31), .B1(new_n604), .B2(new_n605), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT72), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n616), .A2(new_n617), .A3(new_n609), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT32), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n611), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n608), .A2(new_n610), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(KEYINPUT32), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n493), .B(new_n545), .C1(new_n598), .C2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(new_n249), .ZN(G3));
  OAI21_X1  g439(.A(G472), .B1(new_n608), .B2(G902), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n611), .A2(new_n626), .A3(new_n618), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n487), .A2(new_n542), .A3(new_n544), .A4(new_n491), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT91), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n302), .A2(new_n631), .A3(new_n303), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n288), .A2(KEYINPUT91), .A3(new_n298), .A4(new_n300), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n633), .A2(new_n305), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n398), .A2(G902), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT92), .ZN(new_n637));
  AOI21_X1  g451(.A(KEYINPUT33), .B1(new_n405), .B2(new_n637), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n637), .B(KEYINPUT33), .C1(new_n395), .C2(new_n396), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n636), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n397), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n641), .B1(G478), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n364), .A2(new_n366), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(KEYINPUT20), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n647));
  AOI22_X1  g461(.A1(new_n646), .A2(new_n647), .B1(G475), .B2(new_n357), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n635), .A2(new_n416), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n630), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT34), .B(G104), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  AND2_X1   g467(.A1(new_n410), .A2(new_n417), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n369), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n635), .A2(new_n416), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n630), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT35), .B(G107), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  INV_X1    g473(.A(new_n627), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n536), .A2(new_n500), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n532), .A2(KEYINPUT79), .A3(new_n533), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n499), .A2(KEYINPUT36), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n661), .B(new_n662), .C1(KEYINPUT36), .C2(new_n499), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n543), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n542), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n493), .A2(new_n660), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT93), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT37), .B(G110), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G12));
  INV_X1    g487(.A(G900), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n412), .B1(new_n413), .B2(new_n674), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n654), .A2(new_n369), .A3(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n676), .A2(new_n632), .A3(new_n634), .ZN(new_n677));
  INV_X1    g491(.A(new_n495), .ZN(new_n678));
  INV_X1    g492(.A(new_n537), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n679), .B1(new_n663), .B2(new_n499), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n540), .B1(new_n680), .B2(G902), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n538), .A2(KEYINPUT25), .A3(new_n306), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n678), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n668), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n487), .B(new_n491), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n677), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n686), .B1(new_n598), .B2(new_n623), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G128), .ZN(G30));
  AND3_X1   g502(.A1(new_n288), .A2(new_n298), .A3(new_n300), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n300), .B1(new_n288), .B2(new_n298), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g505(.A1(new_n691), .A2(KEYINPUT38), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(KEYINPUT38), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n669), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n648), .A2(new_n654), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n695), .A2(new_n305), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(new_n675), .B(KEYINPUT39), .Z(new_n699));
  NAND3_X1  g513(.A1(new_n487), .A2(new_n491), .A3(new_n699), .ZN(new_n700));
  OR2_X1    g514(.A1(new_n700), .A2(KEYINPUT40), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(KEYINPUT40), .ZN(new_n702));
  INV_X1    g516(.A(new_n578), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n561), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n554), .A2(new_n555), .ZN(new_n705));
  AOI21_X1  g519(.A(G902), .B1(new_n705), .B2(new_n562), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n546), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n707), .B1(new_n621), .B2(KEYINPUT32), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n620), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n698), .A2(new_n701), .A3(new_n702), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G143), .ZN(G45));
  INV_X1    g525(.A(new_n675), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n369), .A2(new_n643), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n632), .A2(new_n713), .A3(new_n634), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n714), .A2(new_n685), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n715), .B1(new_n598), .B2(new_n623), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G146), .ZN(G48));
  INV_X1    g531(.A(new_n623), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n587), .A2(KEYINPUT75), .ZN(new_n719));
  INV_X1    g533(.A(new_n569), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n719), .A2(new_n597), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(G472), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n650), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n467), .A2(KEYINPUT83), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n462), .A2(new_n465), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT12), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n725), .A2(new_n470), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n477), .A2(new_n454), .ZN(new_n730));
  AOI22_X1  g544(.A1(new_n729), .A2(new_n480), .B1(new_n730), .B2(new_n457), .ZN(new_n731));
  OAI21_X1  g545(.A(G469), .B1(new_n731), .B2(G902), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n732), .A2(new_n491), .A3(new_n479), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n723), .A2(new_n724), .A3(new_n545), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT41), .B(G113), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G15));
  OAI211_X1 g550(.A(new_n545), .B(new_n733), .C1(new_n598), .C2(new_n623), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n656), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n195), .ZN(G18));
  AND4_X1   g553(.A1(new_n632), .A2(new_n733), .A3(new_n634), .A4(new_n669), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n740), .B(new_n419), .C1(new_n598), .C2(new_n623), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G119), .ZN(G21));
  NAND3_X1  g556(.A1(new_n557), .A2(new_n591), .A3(new_n567), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n562), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n601), .A2(new_n606), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT94), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n747), .A3(new_n609), .ZN(new_n748));
  AOI22_X1  g562(.A1(new_n743), .A2(new_n562), .B1(new_n601), .B2(new_n606), .ZN(new_n749));
  OAI21_X1  g563(.A(KEYINPUT94), .B1(new_n749), .B2(new_n610), .ZN(new_n750));
  XNOR2_X1  g564(.A(KEYINPUT95), .B(G472), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n608), .B2(G902), .ZN(new_n752));
  AND4_X1   g566(.A1(new_n545), .A2(new_n748), .A3(new_n750), .A4(new_n752), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n632), .A2(new_n634), .A3(new_n696), .ZN(new_n754));
  INV_X1    g568(.A(new_n733), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n415), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n753), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G122), .ZN(G24));
  AND3_X1   g572(.A1(new_n748), .A2(new_n750), .A3(new_n752), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n740), .A2(new_n759), .A3(new_n713), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G125), .ZN(G27));
  AOI21_X1  g575(.A(KEYINPUT97), .B1(new_n691), .B2(new_n305), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n479), .B(new_n486), .C1(new_n484), .C2(KEYINPUT96), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n484), .A2(KEYINPUT96), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n491), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT97), .ZN(new_n766));
  INV_X1    g580(.A(new_n305), .ZN(new_n767));
  NOR4_X1   g581(.A1(new_n689), .A2(new_n690), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n762), .A2(new_n765), .A3(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n723), .A2(new_n545), .A3(new_n713), .A4(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT42), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n479), .A2(new_n486), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n458), .B1(new_n729), .B2(new_n454), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n453), .B1(new_n424), .B2(new_n437), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n459), .A2(new_n774), .ZN(new_n775));
  NOR4_X1   g589(.A1(new_n773), .A2(new_n775), .A3(KEYINPUT96), .A4(new_n421), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n484), .A2(KEYINPUT96), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n490), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n766), .B1(new_n304), .B2(new_n767), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n691), .A2(KEYINPUT97), .A3(new_n305), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n779), .A2(new_n713), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n771), .ZN(new_n783));
  INV_X1    g597(.A(new_n545), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n621), .B(new_n619), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n784), .B1(new_n722), .B2(new_n785), .ZN(new_n786));
  AOI22_X1  g600(.A1(new_n770), .A2(new_n771), .B1(new_n783), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(new_n337), .ZN(G33));
  NAND4_X1  g602(.A1(new_n723), .A2(new_n545), .A3(new_n676), .A4(new_n769), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G134), .ZN(G36));
  NAND2_X1  g604(.A1(new_n780), .A2(new_n781), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n648), .A2(KEYINPUT43), .A3(new_n643), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT99), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n643), .A2(new_n794), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n641), .B(KEYINPUT99), .C1(G478), .C2(new_n642), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n648), .A3(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT43), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n797), .A2(KEYINPUT100), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT100), .B1(new_n797), .B2(new_n798), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n793), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n627), .A3(new_n669), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT44), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n792), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n805), .A2(KEYINPUT101), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(KEYINPUT101), .ZN(new_n807));
  AOI22_X1  g621(.A1(new_n806), .A2(new_n807), .B1(new_n804), .B2(new_n803), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT46), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT45), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n810), .B1(new_n773), .B2(new_n775), .ZN(new_n811));
  OAI211_X1 g625(.A(KEYINPUT45), .B(new_n481), .C1(new_n483), .C2(new_n458), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(new_n812), .A3(G469), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n809), .B1(new_n814), .B2(new_n485), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(KEYINPUT46), .A3(new_n486), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n479), .A3(new_n816), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n817), .A2(new_n491), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n818), .A2(KEYINPUT98), .A3(new_n699), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT98), .B1(new_n818), .B2(new_n699), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n808), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(G137), .ZN(G39));
  INV_X1    g638(.A(new_n713), .ZN(new_n825));
  NOR4_X1   g639(.A1(new_n723), .A2(new_n545), .A3(new_n825), .A4(new_n791), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT102), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n826), .B(new_n827), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n817), .A2(KEYINPUT47), .A3(new_n491), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT47), .B1(new_n817), .B2(new_n491), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(G140), .ZN(G42));
  AND2_X1   g648(.A1(new_n732), .A2(new_n479), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n836), .A2(KEYINPUT49), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(KEYINPUT49), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n648), .A2(new_n491), .A3(new_n305), .A4(new_n643), .ZN(new_n839));
  NOR4_X1   g653(.A1(new_n837), .A2(new_n838), .A3(new_n784), .A4(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n709), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n840), .A2(new_n694), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n545), .B1(new_n598), .B2(new_n623), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n648), .A2(new_n400), .A3(new_n407), .A4(new_n712), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n791), .A2(new_n685), .A3(new_n846), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n845), .A2(new_n676), .B1(new_n723), .B2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT104), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n748), .A2(new_n750), .A3(new_n669), .A4(new_n752), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n769), .A2(new_n849), .A3(new_n713), .A4(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(KEYINPUT104), .B1(new_n782), .B2(new_n850), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n420), .A2(new_n695), .A3(new_n492), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n358), .B(new_n408), .C1(new_n367), .C2(new_n368), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n856), .B1(new_n644), .B2(new_n648), .ZN(new_n857));
  AND4_X1   g671(.A1(new_n305), .A2(new_n857), .A3(new_n304), .A4(new_n416), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n855), .A2(new_n660), .B1(new_n858), .B2(new_n629), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n859), .A2(KEYINPUT103), .A3(new_n624), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT103), .B1(new_n859), .B2(new_n624), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n848), .B(new_n854), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n741), .B(new_n757), .C1(new_n737), .C2(new_n650), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(new_n738), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n783), .A2(new_n786), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n843), .A2(new_n825), .A3(new_n844), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n865), .B1(new_n866), .B2(KEYINPUT42), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n862), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n542), .A2(new_n668), .A3(new_n712), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT105), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT105), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n542), .A2(new_n668), .A3(new_n872), .A4(new_n712), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n709), .A3(new_n754), .A4(new_n779), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n716), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n733), .A2(new_n632), .A3(new_n669), .A4(new_n634), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n877), .A2(new_n825), .ZN(new_n878));
  AOI22_X1  g692(.A1(new_n723), .A2(new_n686), .B1(new_n878), .B2(new_n759), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT52), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n876), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n687), .A2(new_n716), .A3(new_n875), .A4(new_n760), .ZN(new_n882));
  XOR2_X1   g696(.A(KEYINPUT106), .B(KEYINPUT52), .Z(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n881), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n869), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n847), .A2(new_n723), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n854), .A2(new_n789), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT103), .ZN(new_n891));
  INV_X1    g705(.A(new_n624), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n858), .A2(new_n629), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n670), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n891), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n859), .A2(KEYINPUT103), .A3(new_n624), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n890), .A2(new_n897), .A3(new_n867), .A4(new_n864), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n880), .B1(new_n876), .B2(new_n879), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n882), .A2(KEYINPUT52), .ZN(new_n900));
  OAI21_X1  g714(.A(KEYINPUT107), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n882), .A2(KEYINPUT52), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT107), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n881), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n898), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  OAI211_X1 g719(.A(KEYINPUT54), .B(new_n888), .C1(new_n905), .C2(new_n886), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n854), .A2(new_n789), .A3(new_n889), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n908), .B1(new_n895), .B2(new_n896), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n881), .A2(new_n885), .A3(KEYINPUT53), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT108), .ZN(new_n911));
  INV_X1    g725(.A(new_n656), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n723), .A2(new_n912), .A3(new_n545), .A4(new_n733), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n734), .A2(new_n913), .A3(new_n741), .A4(new_n757), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n911), .B1(new_n914), .B2(new_n787), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n864), .A2(new_n867), .A3(KEYINPUT108), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n909), .A2(new_n910), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n907), .B(new_n917), .C1(new_n905), .C2(KEYINPUT53), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n906), .A2(new_n918), .A3(KEYINPUT109), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT109), .B1(new_n906), .B2(new_n918), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AND4_X1   g735(.A1(new_n412), .A2(new_n802), .A3(new_n733), .A4(new_n792), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n786), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT48), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n802), .A2(new_n412), .A3(new_n753), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n925), .A2(new_n635), .A3(new_n733), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n926), .A2(G952), .A3(new_n308), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n841), .A2(new_n545), .A3(new_n412), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n928), .A2(new_n755), .A3(new_n791), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n927), .B1(new_n649), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT114), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n836), .A2(new_n491), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n832), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n925), .A2(new_n792), .ZN(new_n934));
  INV_X1    g748(.A(new_n932), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT114), .B1(new_n831), .B2(new_n935), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n933), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n644), .A2(new_n648), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  AOI22_X1  g753(.A1(new_n929), .A2(new_n939), .B1(new_n922), .B2(new_n851), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n733), .A2(new_n767), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n692), .B2(new_n693), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n802), .A2(new_n412), .A3(new_n942), .A4(new_n753), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT50), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT111), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n944), .A2(KEYINPUT111), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n943), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n925), .A2(KEYINPUT111), .A3(new_n944), .A4(new_n942), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n940), .A2(KEYINPUT51), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n924), .B(new_n930), .C1(new_n937), .C2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT51), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n948), .A2(new_n947), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(KEYINPUT112), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT112), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n948), .A2(new_n954), .A3(new_n947), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n953), .A2(new_n955), .A3(new_n940), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n831), .A2(KEYINPUT110), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n932), .B1(new_n831), .B2(KEYINPUT110), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n934), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n951), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(KEYINPUT113), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT113), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n962), .B(new_n951), .C1(new_n956), .C2(new_n959), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n950), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(KEYINPUT115), .B1(new_n921), .B2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT109), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n901), .A2(new_n904), .ZN(new_n967));
  AOI21_X1  g781(.A(KEYINPUT53), .B1(new_n967), .B2(new_n869), .ZN(new_n968));
  AND4_X1   g782(.A1(new_n909), .A2(new_n910), .A3(new_n915), .A4(new_n916), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n968), .A2(new_n969), .A3(KEYINPUT54), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n886), .B1(new_n967), .B2(new_n869), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n881), .A2(new_n885), .A3(new_n886), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n898), .A2(new_n972), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n971), .A2(new_n907), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n966), .B1(new_n970), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n906), .A2(new_n918), .A3(KEYINPUT109), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n975), .A2(KEYINPUT115), .A3(new_n976), .A4(new_n964), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n411), .A2(new_n308), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n842), .B1(new_n965), .B2(new_n979), .ZN(G75));
  NOR2_X1   g794(.A1(new_n308), .A2(G952), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n968), .A2(new_n969), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n982), .A2(new_n306), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(G210), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT56), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n255), .A2(new_n287), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(new_n285), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT55), .Z(new_n989));
  AOI21_X1  g803(.A(new_n981), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n984), .A2(KEYINPUT116), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT116), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n983), .A2(new_n992), .A3(G210), .ZN(new_n993));
  XNOR2_X1  g807(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n989), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n991), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n990), .A2(new_n996), .ZN(G51));
  INV_X1    g811(.A(new_n981), .ZN(new_n998));
  OAI21_X1  g812(.A(KEYINPUT54), .B1(new_n968), .B2(new_n969), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n918), .ZN(new_n1000));
  XNOR2_X1  g814(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(new_n485), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n731), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n917), .B1(new_n905), .B2(KEYINPUT53), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1004), .A2(G902), .A3(new_n814), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n998), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT119), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g823(.A(KEYINPUT119), .B(new_n998), .C1(new_n1003), .C2(new_n1006), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1009), .A2(new_n1010), .ZN(G54));
  NAND3_X1  g825(.A1(new_n983), .A2(KEYINPUT58), .A3(G475), .ZN(new_n1012));
  INV_X1    g826(.A(new_n364), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1015));
  NOR3_X1   g829(.A1(new_n1014), .A2(new_n1015), .A3(new_n981), .ZN(G60));
  OR2_X1    g830(.A1(new_n638), .A2(new_n640), .ZN(new_n1017));
  XOR2_X1   g831(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1018));
  NOR2_X1   g832(.A1(new_n398), .A2(new_n306), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1018), .B(new_n1019), .ZN(new_n1020));
  AND3_X1   g834(.A1(new_n1000), .A2(new_n1017), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1020), .B1(new_n919), .B2(new_n920), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1017), .ZN(new_n1023));
  AOI211_X1 g837(.A(new_n981), .B(new_n1021), .C1(new_n1022), .C2(new_n1023), .ZN(G63));
  NAND2_X1  g838(.A1(G217), .A2(G902), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1025), .B(KEYINPUT60), .ZN(new_n1026));
  INV_X1    g840(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1004), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n981), .B1(new_n1028), .B2(new_n680), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n982), .A2(new_n1026), .ZN(new_n1030));
  XNOR2_X1  g844(.A(new_n667), .B(KEYINPUT121), .ZN(new_n1031));
  AOI21_X1  g845(.A(KEYINPUT122), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AND4_X1   g846(.A1(KEYINPUT122), .A2(new_n1004), .A3(new_n1027), .A4(new_n1031), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1029), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g848(.A(KEYINPUT61), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  OAI211_X1 g850(.A(new_n1029), .B(KEYINPUT61), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1036), .A2(new_n1037), .ZN(G66));
  OAI21_X1  g852(.A(G953), .B1(new_n414), .B2(new_n282), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n914), .B1(new_n895), .B2(new_n896), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n1039), .B1(new_n1040), .B2(G953), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n987), .B1(G898), .B2(new_n308), .ZN(new_n1042));
  XNOR2_X1  g856(.A(new_n1041), .B(new_n1042), .ZN(G69));
  NAND2_X1  g857(.A1(new_n803), .A2(new_n804), .ZN(new_n1044));
  INV_X1    g858(.A(new_n807), .ZN(new_n1045));
  NOR2_X1   g859(.A1(new_n805), .A2(KEYINPUT101), .ZN(new_n1046));
  OAI21_X1  g860(.A(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n833), .B1(new_n1047), .B2(new_n821), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n879), .A2(new_n716), .ZN(new_n1049));
  OR2_X1    g863(.A1(new_n1049), .A2(KEYINPUT123), .ZN(new_n1050));
  OAI211_X1 g864(.A(new_n754), .B(new_n786), .C1(new_n819), .C2(new_n820), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1049), .A2(KEYINPUT123), .ZN(new_n1052));
  AND3_X1   g866(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n867), .A2(new_n789), .ZN(new_n1054));
  INV_X1    g868(.A(new_n1054), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g870(.A1(new_n1048), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n1057), .A2(new_n308), .ZN(new_n1058));
  XOR2_X1   g872(.A(new_n577), .B(new_n360), .Z(new_n1059));
  AOI21_X1  g873(.A(new_n1059), .B1(G900), .B2(G953), .ZN(new_n1060));
  AOI21_X1  g874(.A(KEYINPUT124), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g875(.A(new_n308), .B1(G227), .B2(G900), .ZN(new_n1062));
  NOR2_X1   g876(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI22_X1  g877(.A1(new_n808), .A2(new_n822), .B1(new_n832), .B2(new_n828), .ZN(new_n1064));
  NAND3_X1  g878(.A1(new_n1050), .A2(new_n710), .A3(new_n1052), .ZN(new_n1065));
  OR2_X1    g879(.A1(new_n1065), .A2(KEYINPUT62), .ZN(new_n1066));
  NAND2_X1  g880(.A1(new_n1065), .A2(KEYINPUT62), .ZN(new_n1067));
  INV_X1    g881(.A(new_n857), .ZN(new_n1068));
  OR4_X1    g882(.A1(new_n843), .A2(new_n700), .A3(new_n791), .A4(new_n1068), .ZN(new_n1069));
  NAND4_X1  g883(.A1(new_n1064), .A2(new_n1066), .A3(new_n1067), .A4(new_n1069), .ZN(new_n1070));
  NAND2_X1  g884(.A1(new_n1070), .A2(new_n308), .ZN(new_n1071));
  AOI22_X1  g885(.A1(new_n1071), .A2(new_n1059), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1072));
  XNOR2_X1  g886(.A(new_n1063), .B(new_n1072), .ZN(G72));
  NAND2_X1  g887(.A1(new_n578), .A2(new_n562), .ZN(new_n1074));
  NAND4_X1  g888(.A1(new_n1064), .A2(new_n1040), .A3(new_n1055), .A4(new_n1053), .ZN(new_n1075));
  NAND2_X1  g889(.A1(G472), .A2(G902), .ZN(new_n1076));
  XOR2_X1   g890(.A(new_n1076), .B(KEYINPUT63), .Z(new_n1077));
  AOI21_X1  g891(.A(new_n1074), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g892(.A(KEYINPUT126), .B1(new_n1078), .B2(new_n981), .ZN(new_n1079));
  INV_X1    g893(.A(KEYINPUT126), .ZN(new_n1080));
  INV_X1    g894(.A(new_n1077), .ZN(new_n1081));
  AOI21_X1  g895(.A(new_n1081), .B1(new_n1057), .B2(new_n1040), .ZN(new_n1082));
  OAI211_X1 g896(.A(new_n1080), .B(new_n998), .C1(new_n1082), .C2(new_n1074), .ZN(new_n1083));
  NAND2_X1  g897(.A1(new_n1079), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g898(.A(new_n1040), .ZN(new_n1085));
  OAI21_X1  g899(.A(new_n1077), .B1(new_n1070), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g900(.A(KEYINPUT125), .ZN(new_n1087));
  NAND2_X1  g901(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g902(.A(KEYINPUT125), .B(new_n1077), .C1(new_n1070), .C2(new_n1085), .ZN(new_n1089));
  NAND4_X1  g903(.A1(new_n1088), .A2(new_n561), .A3(new_n703), .A4(new_n1089), .ZN(new_n1090));
  OAI211_X1 g904(.A(new_n579), .B(new_n584), .C1(new_n583), .C2(new_n600), .ZN(new_n1091));
  NAND2_X1  g905(.A1(new_n1091), .A2(new_n1077), .ZN(new_n1092));
  XNOR2_X1  g906(.A(new_n1092), .B(KEYINPUT127), .ZN(new_n1093));
  OAI211_X1 g907(.A(new_n888), .B(new_n1093), .C1(new_n905), .C2(new_n886), .ZN(new_n1094));
  AND3_X1   g908(.A1(new_n1084), .A2(new_n1090), .A3(new_n1094), .ZN(G57));
endmodule


