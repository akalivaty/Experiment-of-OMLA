//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 0 1 0 0 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 0 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n435, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n558, new_n559, new_n560, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n574, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n609, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1168, new_n1169, new_n1170, new_n1171;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(new_n435));
  INV_X1    g010(.A(new_n435), .ZN(G219));
  XNOR2_X1  g011(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G69), .Z(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G218), .A3(G221), .A4(G220), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n462), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT67), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(new_n462), .A3(G137), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n471), .B1(new_n472), .B2(G2105), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n464), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n473), .A2(G101), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n469), .A2(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n472), .A2(KEYINPUT3), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT3), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(new_n468), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  OAI221_X1 g058(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n468), .C2(G112), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n481), .A2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND3_X1  g063(.A1(new_n464), .A2(G102), .A3(G2104), .ZN(new_n489));
  NAND2_X1  g064(.A1(G114), .A2(G2104), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(new_n462), .B2(G126), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n489), .B1(new_n492), .B2(new_n464), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n468), .A2(new_n462), .A3(G138), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n468), .A2(new_n462), .A3(new_n496), .A4(G138), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n493), .B1(new_n495), .B2(new_n497), .ZN(G164));
  XNOR2_X1  g073(.A(KEYINPUT69), .B(KEYINPUT6), .ZN(new_n499));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT70), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT70), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n505), .A2(KEYINPUT69), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n502), .B(G651), .C1(new_n504), .C2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n500), .A2(KEYINPUT6), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n501), .A2(G543), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT71), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g086(.A(G651), .B1(new_n504), .B2(new_n506), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(KEYINPUT70), .B1(KEYINPUT6), .B2(new_n500), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT72), .B1(new_n514), .B2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT5), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n516), .A2(new_n517), .A3(G543), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n515), .A2(new_n518), .B1(KEYINPUT5), .B2(new_n514), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n513), .A2(G88), .A3(new_n507), .A4(new_n519), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n519), .A2(G62), .ZN(new_n521));
  NAND2_X1  g096(.A1(G75), .A2(G543), .ZN(new_n522));
  XOR2_X1   g097(.A(new_n522), .B(KEYINPUT73), .Z(new_n523));
  OAI21_X1  g098(.A(G651), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n511), .A2(new_n520), .A3(new_n524), .ZN(new_n525));
  NOR3_X1   g100(.A1(new_n509), .A2(KEYINPUT71), .A3(new_n510), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XOR2_X1   g103(.A(new_n528), .B(KEYINPUT7), .Z(new_n529));
  AND2_X1   g104(.A1(G63), .A2(G651), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n529), .B1(new_n519), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G51), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n513), .A2(new_n507), .A3(new_n519), .ZN(new_n533));
  INV_X1    g108(.A(G89), .ZN(new_n534));
  OAI221_X1 g109(.A(new_n531), .B1(new_n532), .B2(new_n509), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT74), .ZN(new_n536));
  INV_X1    g111(.A(new_n533), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G89), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT74), .ZN(new_n539));
  INV_X1    g114(.A(new_n509), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G51), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n538), .A2(new_n539), .A3(new_n541), .A4(new_n531), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n536), .A2(new_n542), .ZN(G168));
  AND2_X1   g118(.A1(new_n537), .A2(G90), .ZN(new_n544));
  INV_X1    g119(.A(G52), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n509), .A2(new_n545), .B1(new_n546), .B2(new_n500), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(G171));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n533), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n519), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n509), .A2(new_n551), .B1(new_n552), .B2(new_n500), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT75), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(G188));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(KEYINPUT76), .A2(G53), .ZN(new_n563));
  NOR3_X1   g138(.A1(new_n509), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n562), .B1(new_n509), .B2(new_n563), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n513), .A2(G91), .A3(new_n507), .A4(new_n519), .ZN(new_n567));
  AND2_X1   g142(.A1(new_n519), .A2(G65), .ZN(new_n568));
  AND2_X1   g143(.A1(G78), .A2(G543), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n565), .A2(new_n566), .A3(new_n567), .A4(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  AND2_X1   g147(.A1(new_n536), .A2(new_n542), .ZN(G286));
  INV_X1    g148(.A(new_n526), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n574), .A2(new_n511), .A3(new_n520), .A4(new_n524), .ZN(G303));
  NAND4_X1  g150(.A1(new_n513), .A2(G87), .A3(new_n507), .A4(new_n519), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n577));
  INV_X1    g152(.A(G49), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n576), .B(new_n577), .C1(new_n578), .C2(new_n509), .ZN(G288));
  NAND2_X1  g154(.A1(new_n537), .A2(G86), .ZN(new_n580));
  INV_X1    g155(.A(G48), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n509), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n519), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(new_n500), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n580), .A2(new_n583), .A3(new_n585), .ZN(G305));
  AOI22_X1  g161(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(new_n500), .ZN(new_n588));
  INV_X1    g163(.A(G47), .ZN(new_n589));
  XNOR2_X1  g164(.A(KEYINPUT77), .B(G85), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  OAI221_X1 g166(.A(new_n588), .B1(new_n589), .B2(new_n509), .C1(new_n533), .C2(new_n591), .ZN(G290));
  XNOR2_X1  g167(.A(KEYINPUT78), .B(G66), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n519), .A2(new_n593), .B1(G79), .B2(G543), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(new_n500), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(new_n540), .B2(G54), .ZN(new_n596));
  AOI21_X1  g171(.A(KEYINPUT10), .B1(new_n537), .B2(G92), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  NOR3_X1   g174(.A1(new_n533), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n596), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(new_n602), .B2(G171), .ZN(G284));
  OAI21_X1  g179(.A(new_n603), .B1(new_n602), .B2(G171), .ZN(G321));
  NAND2_X1  g180(.A1(G299), .A2(new_n602), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G168), .B2(new_n602), .ZN(G297));
  OAI21_X1  g182(.A(new_n606), .B1(G168), .B2(new_n602), .ZN(G280));
  INV_X1    g183(.A(new_n601), .ZN(new_n609));
  XNOR2_X1  g184(.A(KEYINPUT79), .B(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(G860), .B2(new_n610), .ZN(G148));
  NAND2_X1  g186(.A1(new_n609), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g190(.A1(new_n473), .A2(new_n474), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(new_n462), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT12), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT13), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n619), .A2(G2100), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(G2100), .ZN(new_n621));
  AOI22_X1  g196(.A1(G123), .A2(new_n482), .B1(new_n485), .B2(G135), .ZN(new_n622));
  OAI221_X1 g197(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n468), .C2(G111), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(G2096), .Z(new_n625));
  NAND3_X1  g200(.A1(new_n620), .A2(new_n621), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT80), .Z(G156));
  XNOR2_X1  g202(.A(KEYINPUT15), .B(G2430), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2435), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2427), .B(G2438), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n631), .A2(KEYINPUT14), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n634));
  XNOR2_X1  g209(.A(G2451), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n633), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2443), .B(G2446), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(G14), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(new_n639), .B2(new_n640), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(G401));
  XNOR2_X1  g220(.A(G2072), .B(G2078), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT82), .B(KEYINPUT17), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2067), .B(G2678), .Z(new_n649));
  NOR2_X1   g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n649), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n652), .B1(new_n653), .B2(new_n646), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT83), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n653), .A2(new_n646), .A3(new_n651), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT18), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n653), .A2(new_n652), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n658), .B1(new_n648), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2096), .B(G2100), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XNOR2_X1  g238(.A(G1971), .B(G1976), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n665), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n665), .A2(new_n669), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n672));
  OAI221_X1 g247(.A(new_n670), .B1(new_n665), .B2(new_n668), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n672), .B2(new_n671), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT84), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT85), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1991), .B(G1996), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1981), .B(G1986), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n679), .B(new_n680), .Z(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n676), .A2(new_n677), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n676), .A2(new_n677), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n684), .A2(new_n681), .A3(new_n685), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n683), .A2(new_n686), .ZN(G229));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G6), .ZN(new_n689));
  INV_X1    g264(.A(G305), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n689), .B1(new_n690), .B2(new_n688), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT32), .B(G1981), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(G16), .A2(G23), .ZN(new_n694));
  INV_X1    g269(.A(G288), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n694), .B1(new_n695), .B2(G16), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT33), .B(G1976), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n688), .A2(G22), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G166), .B2(new_n688), .ZN(new_n700));
  INV_X1    g275(.A(G1971), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n693), .A2(new_n698), .A3(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT34), .Z(new_n704));
  NAND2_X1  g279(.A1(new_n482), .A2(G119), .ZN(new_n705));
  OAI221_X1 g280(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n468), .C2(G107), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n485), .A2(G131), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  MUX2_X1   g283(.A(G25), .B(new_n708), .S(G29), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT87), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT35), .B(G1991), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT86), .Z(new_n712));
  XOR2_X1   g287(.A(new_n710), .B(new_n712), .Z(new_n713));
  NAND2_X1  g288(.A1(new_n688), .A2(G24), .ZN(new_n714));
  INV_X1    g289(.A(G290), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n688), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n716), .A2(G1986), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(G1986), .ZN(new_n718));
  NOR4_X1   g293(.A1(new_n713), .A2(new_n717), .A3(KEYINPUT88), .A4(new_n718), .ZN(new_n719));
  AND3_X1   g294(.A1(new_n704), .A2(KEYINPUT36), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(KEYINPUT36), .B1(new_n704), .B2(new_n719), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n688), .A2(G19), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT89), .Z(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(new_n554), .B2(new_n688), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(G1341), .Z(new_n725));
  NOR2_X1   g300(.A1(G4), .A2(G16), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n609), .B2(G16), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n725), .B1(G1348), .B2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT28), .ZN(new_n729));
  INV_X1    g304(.A(G29), .ZN(new_n730));
  AND3_X1   g305(.A1(new_n729), .A2(new_n730), .A3(G26), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT91), .ZN(new_n732));
  INV_X1    g307(.A(G128), .ZN(new_n733));
  NOR3_X1   g308(.A1(new_n481), .A2(new_n468), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT90), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n468), .A2(G116), .ZN(new_n736));
  OAI21_X1  g311(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n736), .A2(new_n738), .B1(new_n485), .B2(G140), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n732), .B1(new_n735), .B2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n735), .A2(new_n732), .A3(new_n739), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G29), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n729), .B1(G26), .B2(new_n730), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n731), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT92), .B(G2067), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  AOI211_X1 g323(.A(new_n728), .B(new_n748), .C1(G1348), .C2(new_n727), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT97), .B(KEYINPUT23), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n688), .A2(G20), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G299), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(new_n688), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT98), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G1956), .ZN(new_n756));
  NOR2_X1   g331(.A1(G16), .A2(G21), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G168), .B2(G16), .ZN(new_n758));
  INV_X1    g333(.A(G1966), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n730), .A2(G35), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G162), .B2(new_n730), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT29), .Z(new_n763));
  INV_X1    g338(.A(G2090), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(G29), .A2(G32), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n616), .A2(G105), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT96), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n482), .A2(G129), .ZN(new_n769));
  NAND3_X1  g344(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT26), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G141), .B2(new_n485), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n768), .A2(new_n769), .A3(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n766), .B1(new_n774), .B2(G29), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT27), .B(G1996), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT30), .B(G28), .ZN(new_n778));
  OR2_X1    g353(.A1(KEYINPUT31), .A2(G11), .ZN(new_n779));
  NAND2_X1  g354(.A1(KEYINPUT31), .A2(G11), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n778), .A2(new_n730), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AND2_X1   g356(.A1(KEYINPUT24), .A2(G34), .ZN(new_n782));
  NOR2_X1   g357(.A1(KEYINPUT24), .A2(G34), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n730), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT94), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G160), .B2(G29), .ZN(new_n787));
  OAI221_X1 g362(.A(new_n781), .B1(new_n730), .B2(new_n624), .C1(new_n787), .C2(G2084), .ZN(new_n788));
  INV_X1    g363(.A(G2078), .ZN(new_n789));
  NOR2_X1   g364(.A1(G27), .A2(G29), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G164), .B2(G29), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n788), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n763), .A2(new_n764), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n765), .A2(new_n777), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n730), .A2(G33), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT25), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G139), .B2(new_n485), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(new_n468), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT93), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n796), .B1(new_n804), .B2(new_n730), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G2072), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n787), .A2(G2084), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(KEYINPUT95), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(KEYINPUT95), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n808), .B(new_n809), .C1(new_n789), .C2(new_n792), .ZN(new_n810));
  NOR2_X1   g385(.A1(G5), .A2(G16), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G171), .B2(G16), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1961), .ZN(new_n813));
  NOR4_X1   g388(.A1(new_n795), .A2(new_n806), .A3(new_n810), .A4(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n749), .A2(new_n756), .A3(new_n760), .A4(new_n814), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n720), .A2(new_n721), .A3(new_n815), .ZN(G311));
  INV_X1    g391(.A(G311), .ZN(G150));
  OR2_X1    g392(.A1(new_n550), .A2(new_n553), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n513), .A2(G93), .A3(new_n507), .A4(new_n519), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(G55), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  OAI22_X1  g397(.A1(new_n509), .A2(new_n821), .B1(new_n822), .B2(new_n500), .ZN(new_n823));
  OAI21_X1  g398(.A(KEYINPUT99), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n540), .A2(G55), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n822), .A2(new_n500), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT99), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n825), .A2(new_n826), .A3(new_n827), .A4(new_n819), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n818), .A2(new_n824), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n820), .A2(new_n823), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n554), .A2(new_n830), .A3(new_n827), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT38), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n609), .A2(G559), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n833), .B(new_n834), .Z(new_n835));
  AOI21_X1  g410(.A(G860), .B1(new_n835), .B2(KEYINPUT39), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(KEYINPUT39), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n836), .B1(new_n837), .B2(KEYINPUT100), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n837), .A2(KEYINPUT100), .ZN(new_n839));
  INV_X1    g414(.A(new_n830), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n840), .A2(KEYINPUT37), .A3(G860), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(KEYINPUT37), .B1(new_n840), .B2(G860), .ZN(new_n843));
  OAI22_X1  g418(.A1(new_n838), .A2(new_n839), .B1(new_n842), .B2(new_n843), .ZN(G145));
  AOI22_X1  g419(.A1(G130), .A2(new_n482), .B1(new_n485), .B2(G142), .ZN(new_n845));
  OAI221_X1 g420(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n468), .C2(G118), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n708), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT101), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n618), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n741), .A2(new_n774), .A3(new_n742), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n774), .B1(new_n741), .B2(new_n742), .ZN(new_n854));
  OAI21_X1  g429(.A(G164), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n854), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n495), .A2(new_n497), .ZN(new_n857));
  INV_X1    g432(.A(new_n489), .ZN(new_n858));
  INV_X1    g433(.A(G126), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n490), .B1(new_n481), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n858), .B1(new_n860), .B2(G2105), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n856), .A2(new_n852), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n855), .A2(new_n863), .A3(new_n804), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n804), .B1(new_n855), .B2(new_n863), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n851), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n855), .A2(new_n863), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(new_n803), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n869), .A2(new_n850), .A3(new_n864), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n867), .A2(KEYINPUT102), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n864), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT102), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(new_n873), .A3(new_n851), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n624), .B(G160), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(G162), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n871), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n876), .B1(new_n872), .B2(new_n851), .ZN(new_n878));
  AOI21_X1  g453(.A(G37), .B1(new_n878), .B2(new_n870), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT103), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n877), .A2(new_n879), .A3(KEYINPUT103), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n877), .A2(new_n879), .A3(KEYINPUT103), .ZN(new_n885));
  OAI21_X1  g460(.A(KEYINPUT40), .B1(new_n885), .B2(new_n880), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(G395));
  XNOR2_X1  g462(.A(new_n612), .B(new_n832), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n609), .A2(G299), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n753), .A2(new_n601), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n889), .A2(KEYINPUT41), .A3(new_n890), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n888), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  XOR2_X1   g470(.A(new_n895), .B(KEYINPUT105), .Z(new_n896));
  NAND2_X1  g471(.A1(new_n888), .A2(new_n891), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n897), .B(KEYINPUT104), .Z(new_n898));
  NAND2_X1  g473(.A1(new_n715), .A2(new_n695), .ZN(new_n899));
  NAND2_X1  g474(.A1(G290), .A2(G288), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n899), .A2(new_n900), .A3(G303), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(G303), .B1(new_n899), .B2(new_n900), .ZN(new_n903));
  OAI21_X1  g478(.A(G305), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n899), .A2(new_n900), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(G166), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n906), .A2(new_n690), .A3(new_n901), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT42), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n896), .A2(new_n898), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n909), .B1(new_n896), .B2(new_n898), .ZN(new_n911));
  OAI21_X1  g486(.A(G868), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n912), .B1(G868), .B2(new_n830), .ZN(G295));
  OAI21_X1  g488(.A(new_n912), .B1(G868), .B2(new_n830), .ZN(G331));
  NAND2_X1  g489(.A1(new_n904), .A2(new_n907), .ZN(new_n915));
  NAND3_X1  g490(.A1(G168), .A2(new_n829), .A3(new_n831), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(G168), .B1(new_n831), .B2(new_n829), .ZN(new_n918));
  OAI21_X1  g493(.A(G301), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n832), .A2(G286), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n920), .A2(G171), .A3(new_n916), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n919), .A2(new_n891), .A3(new_n921), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n915), .A2(new_n922), .A3(KEYINPUT106), .ZN(new_n923));
  INV_X1    g498(.A(new_n922), .ZN(new_n924));
  AOI22_X1  g499(.A1(new_n919), .A2(new_n921), .B1(new_n893), .B2(new_n894), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n915), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n919), .A2(new_n921), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n893), .A2(new_n894), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n929), .A2(new_n908), .A3(new_n922), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n923), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  AND4_X1   g506(.A1(KEYINPUT106), .A2(new_n929), .A3(new_n915), .A4(new_n922), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n933));
  NOR4_X1   g508(.A1(new_n931), .A2(new_n932), .A3(new_n933), .A4(G37), .ZN(new_n934));
  INV_X1    g509(.A(G37), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n926), .A2(new_n930), .A3(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n936), .A2(new_n933), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT44), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n939));
  NOR4_X1   g514(.A1(new_n931), .A2(new_n932), .A3(KEYINPUT43), .A4(G37), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n938), .A2(new_n942), .ZN(G397));
  INV_X1    g518(.A(KEYINPUT45), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n944), .B1(G164), .B2(G1384), .ZN(new_n945));
  INV_X1    g520(.A(G40), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n469), .A2(new_n476), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(G1384), .B1(new_n857), .B2(new_n861), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT45), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n945), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n950), .A2(KEYINPUT116), .A3(new_n759), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT50), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n947), .B1(new_n948), .B2(new_n952), .ZN(new_n953));
  AOI211_X1 g528(.A(KEYINPUT50), .B(G1384), .C1(new_n857), .C2(new_n861), .ZN(new_n954));
  OR3_X1    g529(.A1(new_n953), .A2(G2084), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT116), .B1(new_n950), .B2(new_n759), .ZN(new_n957));
  OR2_X1    g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n958), .A2(G8), .A3(G168), .ZN(new_n959));
  INV_X1    g534(.A(G1976), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT52), .B1(G288), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(G8), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n962), .B1(new_n948), .B2(new_n947), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n961), .B(new_n963), .C1(new_n960), .C2(G288), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n963), .B1(new_n960), .B2(G288), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT52), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT113), .ZN(new_n968));
  INV_X1    g543(.A(G86), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n585), .B1(new_n969), .B2(new_n533), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT49), .B1(new_n970), .B2(new_n582), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT49), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n580), .A2(new_n972), .A3(new_n583), .A4(new_n585), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT114), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n585), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(G1981), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n971), .A2(G1981), .A3(new_n973), .A4(new_n976), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(new_n963), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT113), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n964), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n968), .A2(new_n980), .A3(KEYINPUT63), .A4(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n959), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n950), .A2(KEYINPUT110), .ZN(new_n985));
  INV_X1    g560(.A(G1384), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT45), .B1(new_n862), .B2(new_n986), .ZN(new_n987));
  AOI211_X1 g562(.A(new_n944), .B(G1384), .C1(new_n857), .C2(new_n861), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n989), .A2(new_n990), .A3(new_n947), .ZN(new_n991));
  AOI21_X1  g566(.A(G1971), .B1(new_n985), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n948), .A2(new_n952), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n993), .A2(new_n947), .A3(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n995), .A2(G2090), .ZN(new_n996));
  OAI21_X1  g571(.A(G8), .B1(new_n992), .B2(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(KEYINPUT55), .B(G8), .C1(new_n525), .C2(new_n526), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT111), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n1000), .B1(G166), .B2(new_n962), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT111), .ZN(new_n1002));
  NAND4_X1  g577(.A1(G303), .A2(new_n1002), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n997), .A2(new_n999), .A3(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n999), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT112), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n999), .A2(new_n1001), .A3(new_n1003), .A4(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n990), .B1(new_n989), .B2(new_n947), .ZN(new_n1011));
  INV_X1    g586(.A(new_n947), .ZN(new_n1012));
  NOR4_X1   g587(.A1(new_n987), .A2(new_n988), .A3(KEYINPUT110), .A4(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n701), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n996), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n962), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1010), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n984), .A2(new_n1005), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT117), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT117), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n984), .A2(new_n1020), .A3(new_n1005), .A4(new_n1017), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1022), .B1(new_n1017), .B2(new_n1005), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n968), .A2(new_n980), .A3(new_n982), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1006), .B1(new_n1025), .B2(G8), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1024), .B1(new_n1026), .B2(KEYINPUT115), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1023), .A2(new_n1027), .A3(new_n959), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1019), .B(new_n1021), .C1(new_n1028), .C2(KEYINPUT63), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT51), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1030), .B(G8), .C1(new_n956), .C2(new_n957), .ZN(new_n1031));
  NOR2_X1   g606(.A1(G168), .A2(new_n962), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1032), .B1(KEYINPUT124), .B2(KEYINPUT51), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(G8), .B1(new_n956), .B2(new_n957), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT123), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g612(.A(KEYINPUT123), .B(G8), .C1(new_n956), .C2(new_n957), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1032), .A2(KEYINPUT124), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1034), .B1(new_n1040), .B2(KEYINPUT51), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n958), .A2(new_n1032), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT62), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT62), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n1035), .A2(new_n1036), .B1(KEYINPUT124), .B2(new_n1032), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1030), .B1(new_n1046), .B2(new_n1038), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1045), .B(new_n1042), .C1(new_n1047), .C2(new_n1034), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n985), .A2(new_n991), .A3(new_n789), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n1050));
  INV_X1    g625(.A(G1961), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1049), .A2(new_n1050), .B1(new_n1051), .B2(new_n995), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n989), .A2(KEYINPUT53), .A3(new_n789), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1052), .B1(new_n1012), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(G171), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n1023), .A2(new_n1027), .A3(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1044), .A2(new_n1048), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1348), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(new_n953), .B2(new_n954), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n1060));
  INV_X1    g635(.A(G2067), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n948), .A2(new_n1061), .A3(new_n947), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1059), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1060), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1064));
  OR3_X1    g639(.A1(new_n1063), .A2(new_n1064), .A3(KEYINPUT60), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT121), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1059), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n601), .B1(new_n1069), .B2(KEYINPUT60), .ZN(new_n1070));
  OAI211_X1 g645(.A(KEYINPUT60), .B(new_n601), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1065), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT56), .B(G2072), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n945), .A2(new_n947), .A3(new_n949), .A4(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT120), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n989), .A2(new_n1077), .A3(new_n947), .A4(new_n1074), .ZN(new_n1078));
  INV_X1    g653(.A(G1956), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n995), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1076), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n566), .A2(new_n567), .A3(new_n570), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1082), .B1(new_n1083), .B2(new_n564), .ZN(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(G299), .A2(new_n1082), .A3(new_n1085), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1081), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1091));
  AOI22_X1  g666(.A1(KEYINPUT120), .A2(new_n1075), .B1(new_n995), .B2(new_n1079), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1091), .B1(new_n1092), .B2(new_n1078), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT61), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1081), .A2(new_n1089), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT61), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1092), .A2(new_n1078), .A3(new_n1091), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT58), .B(G1341), .Z(new_n1100));
  INV_X1    g675(.A(new_n948), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1100), .B1(new_n1101), .B2(new_n1012), .ZN(new_n1102));
  OR2_X1    g677(.A1(new_n1102), .A2(KEYINPUT122), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(KEYINPUT122), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1103), .B(new_n1104), .C1(G1996), .C2(new_n950), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1105), .A2(KEYINPUT59), .A3(new_n554), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT59), .B1(new_n1105), .B2(new_n554), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1073), .A2(new_n1099), .A3(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1069), .A2(new_n601), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1093), .B1(new_n1110), .B2(new_n1097), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1023), .A2(new_n1027), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1042), .B1(new_n1047), .B2(new_n1034), .ZN(new_n1114));
  XOR2_X1   g689(.A(G171), .B(KEYINPUT54), .Z(new_n1115));
  INV_X1    g690(.A(new_n1053), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n476), .A2(KEYINPUT125), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n476), .A2(KEYINPUT125), .ZN(new_n1118));
  NOR4_X1   g693(.A1(new_n1117), .A2(new_n1118), .A3(new_n946), .A4(new_n469), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1115), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1054), .A2(new_n1115), .B1(new_n1120), .B2(new_n1052), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .A4(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1017), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n980), .A2(new_n960), .A3(new_n695), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(G1981), .B2(G305), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1123), .A2(new_n1024), .B1(new_n1125), .B2(new_n963), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1029), .A2(new_n1057), .A3(new_n1122), .A4(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n945), .A2(new_n1012), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1128), .A2(G1996), .A3(new_n773), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1129), .B(KEYINPUT107), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n743), .B(new_n1061), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n1131), .A2(KEYINPUT108), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(KEYINPUT108), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1132), .B(new_n1133), .C1(G1996), .C2(new_n773), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1130), .B1(new_n1134), .B2(new_n1128), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n708), .A2(new_n712), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n708), .A2(new_n712), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1128), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(G290), .B(G1986), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(new_n1128), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1135), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1141), .B(KEYINPUT109), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1127), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1128), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1144), .A2(G1996), .ZN(new_n1145));
  NAND2_X1  g720(.A1(KEYINPUT126), .A2(KEYINPUT46), .ZN(new_n1146));
  XOR2_X1   g721(.A(new_n1145), .B(new_n1146), .Z(new_n1147));
  NOR2_X1   g722(.A1(KEYINPUT126), .A2(KEYINPUT46), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  XOR2_X1   g724(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n1150));
  AND2_X1   g725(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1151), .A2(new_n774), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1149), .B(new_n1150), .C1(new_n1152), .C2(new_n1144), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1150), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1144), .B1(new_n1151), .B2(new_n774), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1149), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1154), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1144), .A2(G1986), .A3(G290), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT48), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1153), .B(new_n1157), .C1(new_n1158), .C2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n741), .A2(new_n1061), .A3(new_n742), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1144), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1143), .A2(new_n1165), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g741(.A1(new_n940), .A2(new_n941), .ZN(new_n1168));
  OR3_X1    g742(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1169));
  AOI21_X1  g743(.A(new_n1169), .B1(new_n683), .B2(new_n686), .ZN(new_n1170));
  OAI21_X1  g744(.A(new_n1170), .B1(new_n885), .B2(new_n880), .ZN(new_n1171));
  NOR2_X1   g745(.A1(new_n1168), .A2(new_n1171), .ZN(G308));
  OAI221_X1 g746(.A(new_n1170), .B1(new_n885), .B2(new_n880), .C1(new_n940), .C2(new_n941), .ZN(G225));
endmodule


