

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732;

  BUF_X1 U369 ( .A(n672), .Z(n347) );
  XNOR2_X1 U370 ( .A(n377), .B(n376), .ZN(n594) );
  OR2_X1 U371 ( .A1(n516), .A2(KEYINPUT64), .ZN(n517) );
  NOR2_X1 U372 ( .A1(n577), .A2(n404), .ZN(n403) );
  AND2_X1 U373 ( .A1(n506), .A2(n617), .ZN(n665) );
  XNOR2_X1 U374 ( .A(n529), .B(KEYINPUT99), .ZN(n530) );
  INV_X1 U375 ( .A(n568), .ZN(n536) );
  XNOR2_X1 U376 ( .A(G122), .B(n418), .ZN(n481) );
  NAND2_X1 U377 ( .A1(n594), .A2(n398), .ZN(n717) );
  INV_X1 U378 ( .A(n566), .ZN(n567) );
  NAND2_X1 U379 ( .A1(n617), .A2(n549), .ZN(n566) );
  XNOR2_X2 U380 ( .A(KEYINPUT75), .B(KEYINPUT74), .ZN(n373) );
  NAND2_X1 U381 ( .A1(n607), .A2(n598), .ZN(n426) );
  XNOR2_X1 U382 ( .A(n408), .B(n407), .ZN(n607) );
  AND2_X2 U383 ( .A1(n519), .A2(n513), .ZN(n514) );
  OR2_X2 U384 ( .A1(n601), .A2(G902), .ZN(n392) );
  XNOR2_X1 U385 ( .A(n419), .B(n481), .ZN(n701) );
  XNOR2_X1 U386 ( .A(KEYINPUT10), .B(G125), .ZN(n382) );
  INV_X1 U387 ( .A(G953), .ZN(n718) );
  OR2_X2 U388 ( .A1(n695), .A2(n396), .ZN(n612) );
  XNOR2_X2 U389 ( .A(KEYINPUT31), .B(n530), .ZN(n676) );
  NOR2_X2 U390 ( .A1(n527), .A2(n536), .ZN(n472) );
  NOR2_X1 U391 ( .A1(n572), .A2(n571), .ZN(n679) );
  XNOR2_X1 U392 ( .A(n370), .B(G478), .ZN(n531) );
  XNOR2_X1 U393 ( .A(n455), .B(n454), .ZN(n617) );
  XNOR2_X1 U394 ( .A(n711), .B(n462), .ZN(n601) );
  XNOR2_X1 U395 ( .A(n383), .B(n411), .ZN(n711) );
  INV_X1 U396 ( .A(n457), .ZN(n411) );
  XNOR2_X1 U397 ( .A(n460), .B(n702), .ZN(n470) );
  NOR2_X1 U398 ( .A1(G953), .A2(G237), .ZN(n474) );
  XNOR2_X1 U399 ( .A(G101), .B(n712), .ZN(n460) );
  XNOR2_X1 U400 ( .A(n391), .B(G469), .ZN(n390) );
  INV_X1 U401 ( .A(KEYINPUT71), .ZN(n391) );
  XNOR2_X1 U402 ( .A(G119), .B(KEYINPUT3), .ZN(n425) );
  XNOR2_X1 U403 ( .A(n583), .B(n415), .ZN(n595) );
  INV_X1 U404 ( .A(KEYINPUT39), .ZN(n415) );
  AND2_X1 U405 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U406 ( .A1(n364), .A2(n573), .ZN(n404) );
  AND2_X1 U407 ( .A1(n539), .A2(n540), .ZN(n368) );
  XOR2_X1 U408 ( .A(KEYINPUT18), .B(KEYINPUT82), .Z(n423) );
  NOR2_X1 U409 ( .A1(n730), .A2(n729), .ZN(n585) );
  XNOR2_X1 U410 ( .A(n400), .B(n379), .ZN(n378) );
  INV_X1 U411 ( .A(KEYINPUT70), .ZN(n379) );
  NAND2_X1 U412 ( .A1(n403), .A2(n401), .ZN(n400) );
  XNOR2_X1 U413 ( .A(KEYINPUT4), .B(G146), .ZN(n712) );
  XOR2_X1 U414 ( .A(G116), .B(G107), .Z(n491) );
  XNOR2_X1 U415 ( .A(G104), .B(G107), .ZN(n387) );
  XNOR2_X1 U416 ( .A(G140), .B(KEYINPUT93), .ZN(n388) );
  XNOR2_X1 U417 ( .A(n459), .B(n458), .ZN(n389) );
  XNOR2_X1 U418 ( .A(G137), .B(KEYINPUT5), .ZN(n466) );
  INV_X1 U419 ( .A(G113), .ZN(n465) );
  XOR2_X1 U420 ( .A(KEYINPUT79), .B(G116), .Z(n464) );
  XNOR2_X1 U421 ( .A(n470), .B(n350), .ZN(n407) );
  XNOR2_X1 U422 ( .A(n701), .B(n409), .ZN(n408) );
  XNOR2_X1 U423 ( .A(n550), .B(KEYINPUT6), .ZN(n568) );
  NOR2_X1 U424 ( .A1(n688), .A2(G902), .ZN(n370) );
  XNOR2_X1 U425 ( .A(n524), .B(n363), .ZN(n582) );
  INV_X1 U426 ( .A(KEYINPUT98), .ZN(n363) );
  XNOR2_X1 U427 ( .A(n504), .B(n503), .ZN(n507) );
  XNOR2_X1 U428 ( .A(n382), .B(n381), .ZN(n715) );
  INV_X1 U429 ( .A(G140), .ZN(n381) );
  XNOR2_X1 U430 ( .A(G131), .B(G143), .ZN(n478) );
  XOR2_X1 U431 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n476) );
  XNOR2_X1 U432 ( .A(n424), .B(n410), .ZN(n409) );
  XNOR2_X1 U433 ( .A(n421), .B(KEYINPUT17), .ZN(n410) );
  XOR2_X1 U434 ( .A(KEYINPUT89), .B(G125), .Z(n421) );
  AND2_X1 U435 ( .A1(n727), .A2(n593), .ZN(n398) );
  INV_X1 U436 ( .A(KEYINPUT48), .ZN(n376) );
  XNOR2_X1 U437 ( .A(G902), .B(KEYINPUT15), .ZN(n598) );
  XNOR2_X1 U438 ( .A(n374), .B(n491), .ZN(n419) );
  XNOR2_X1 U439 ( .A(n373), .B(n372), .ZN(n374) );
  INV_X1 U440 ( .A(KEYINPUT16), .ZN(n372) );
  INV_X1 U441 ( .A(KEYINPUT45), .ZN(n399) );
  XNOR2_X1 U442 ( .A(n715), .B(n380), .ZN(n483) );
  INV_X1 U443 ( .A(G146), .ZN(n380) );
  XNOR2_X1 U444 ( .A(G110), .B(KEYINPUT23), .ZN(n443) );
  XNOR2_X1 U445 ( .A(G128), .B(G119), .ZN(n441) );
  XOR2_X1 U446 ( .A(G137), .B(KEYINPUT69), .Z(n457) );
  XNOR2_X1 U447 ( .A(n439), .B(n365), .ZN(n487) );
  XNOR2_X1 U448 ( .A(n440), .B(KEYINPUT86), .ZN(n365) );
  XOR2_X1 U449 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n440) );
  XNOR2_X1 U450 ( .A(G122), .B(KEYINPUT101), .ZN(n488) );
  XOR2_X1 U451 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n489) );
  XNOR2_X1 U452 ( .A(n492), .B(n369), .ZN(n493) );
  INV_X1 U453 ( .A(n491), .ZN(n369) );
  XNOR2_X1 U454 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U455 ( .A(n389), .B(n386), .ZN(n461) );
  XNOR2_X1 U456 ( .A(n388), .B(n387), .ZN(n386) );
  NAND2_X1 U457 ( .A1(G234), .A2(G237), .ZN(n430) );
  NAND2_X1 U458 ( .A1(n394), .A2(n568), .ZN(n587) );
  AND2_X1 U459 ( .A1(n567), .A2(n349), .ZN(n394) );
  XNOR2_X1 U460 ( .A(n565), .B(n428), .ZN(n555) );
  XNOR2_X1 U461 ( .A(n470), .B(n469), .ZN(n393) );
  INV_X1 U462 ( .A(n608), .ZN(n610) );
  XNOR2_X1 U463 ( .A(n414), .B(n412), .ZN(n729) );
  XNOR2_X1 U464 ( .A(n584), .B(n413), .ZN(n412) );
  INV_X1 U465 ( .A(KEYINPUT107), .ZN(n413) );
  XNOR2_X1 U466 ( .A(n499), .B(n500), .ZN(n384) );
  XNOR2_X1 U467 ( .A(n512), .B(n511), .ZN(n731) );
  OR2_X1 U468 ( .A1(n563), .A2(n564), .ZN(n364) );
  NOR2_X1 U469 ( .A1(n375), .A2(n555), .ZN(n672) );
  OR2_X1 U470 ( .A1(n623), .A2(n621), .ZN(n405) );
  NOR2_X1 U471 ( .A1(n507), .A2(n623), .ZN(n406) );
  XNOR2_X1 U472 ( .A(n687), .B(n366), .ZN(n689) );
  XNOR2_X1 U473 ( .A(n688), .B(KEYINPUT120), .ZN(n366) );
  INV_X1 U474 ( .A(KEYINPUT60), .ZN(n361) );
  XNOR2_X1 U475 ( .A(n471), .B(G472), .ZN(n550) );
  XOR2_X1 U476 ( .A(n613), .B(KEYINPUT84), .Z(n348) );
  AND2_X1 U477 ( .A1(n531), .A2(n395), .ZN(n349) );
  XOR2_X1 U478 ( .A(n456), .B(n458), .Z(n350) );
  AND2_X1 U479 ( .A1(n427), .A2(G210), .ZN(n351) );
  AND2_X1 U480 ( .A1(n541), .A2(n368), .ZN(n352) );
  NOR2_X1 U481 ( .A1(n634), .A2(n375), .ZN(n353) );
  XNOR2_X1 U482 ( .A(n682), .B(KEYINPUT59), .ZN(n354) );
  XOR2_X1 U483 ( .A(n657), .B(KEYINPUT62), .Z(n355) );
  XOR2_X1 U484 ( .A(n610), .B(n609), .Z(n356) );
  NOR2_X1 U485 ( .A1(G952), .A2(n718), .ZN(n694) );
  INV_X1 U486 ( .A(n694), .ZN(n684) );
  XOR2_X1 U487 ( .A(KEYINPUT56), .B(KEYINPUT118), .Z(n357) );
  BUF_X2 U488 ( .A(n686), .Z(n690) );
  XNOR2_X1 U489 ( .A(n358), .B(n357), .ZN(G51) );
  NAND2_X1 U490 ( .A1(n360), .A2(n684), .ZN(n358) );
  XNOR2_X1 U491 ( .A(n359), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U492 ( .A1(n367), .A2(n684), .ZN(n359) );
  NOR2_X2 U493 ( .A1(n665), .A2(n731), .ZN(n519) );
  NOR2_X1 U494 ( .A1(n526), .A2(n502), .ZN(n504) );
  XNOR2_X1 U495 ( .A(n611), .B(n356), .ZN(n360) );
  XNOR2_X1 U496 ( .A(n362), .B(n361), .ZN(G60) );
  NAND2_X1 U497 ( .A1(n685), .A2(n684), .ZN(n362) );
  XNOR2_X1 U498 ( .A(n658), .B(n355), .ZN(n367) );
  NAND2_X1 U499 ( .A1(n378), .A2(n586), .ZN(n377) );
  INV_X1 U500 ( .A(n364), .ZN(n670) );
  XNOR2_X1 U501 ( .A(n505), .B(KEYINPUT66), .ZN(n506) );
  OR2_X2 U502 ( .A1(n543), .A2(n544), .ZN(n371) );
  XNOR2_X2 U503 ( .A(n456), .B(G134), .ZN(n492) );
  XNOR2_X2 U504 ( .A(n371), .B(n399), .ZN(n695) );
  OR2_X1 U505 ( .A1(n728), .A2(n513), .ZN(n541) );
  NAND2_X1 U506 ( .A1(n498), .A2(n497), .ZN(n385) );
  NOR2_X1 U507 ( .A1(n507), .A2(n405), .ZN(n505) );
  NOR2_X2 U508 ( .A1(n555), .A2(n433), .ZN(n435) );
  NAND2_X1 U509 ( .A1(n553), .A2(n554), .ZN(n375) );
  XNOR2_X1 U510 ( .A(n383), .B(n393), .ZN(n657) );
  XNOR2_X2 U511 ( .A(n492), .B(G131), .ZN(n383) );
  XNOR2_X2 U512 ( .A(n385), .B(n384), .ZN(n728) );
  XNOR2_X2 U513 ( .A(n554), .B(KEYINPUT1), .ZN(n623) );
  XNOR2_X2 U514 ( .A(n392), .B(n390), .ZN(n554) );
  INV_X1 U515 ( .A(n531), .ZN(n532) );
  INV_X1 U516 ( .A(n533), .ZN(n395) );
  NOR2_X1 U517 ( .A1(n695), .A2(n717), .ZN(n597) );
  NAND2_X1 U518 ( .A1(n594), .A2(n397), .ZN(n396) );
  AND2_X1 U519 ( .A1(n398), .A2(KEYINPUT2), .ZN(n397) );
  XNOR2_X1 U520 ( .A(n679), .B(n402), .ZN(n401) );
  INV_X1 U521 ( .A(KEYINPUT88), .ZN(n402) );
  NAND2_X1 U522 ( .A1(n406), .A2(n536), .ZN(n537) );
  NAND2_X1 U523 ( .A1(n592), .A2(n635), .ZN(n565) );
  XNOR2_X2 U524 ( .A(n426), .B(n351), .ZN(n592) );
  NAND2_X1 U525 ( .A1(n595), .A2(n349), .ZN(n414) );
  XNOR2_X1 U526 ( .A(n605), .B(n604), .ZN(n606) );
  NOR2_X2 U527 ( .A1(n613), .A2(n600), .ZN(n686) );
  AND2_X1 U528 ( .A1(n606), .A2(n684), .ZN(G54) );
  INV_X1 U529 ( .A(KEYINPUT11), .ZN(n477) );
  XNOR2_X1 U530 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U531 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U532 ( .A(n480), .B(n479), .ZN(n482) );
  XNOR2_X1 U533 ( .A(n468), .B(n467), .ZN(n469) );
  INV_X1 U534 ( .A(n681), .ZN(n593) );
  INV_X1 U535 ( .A(KEYINPUT22), .ZN(n503) );
  XNOR2_X1 U536 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U537 ( .A(n683), .B(n354), .ZN(n685) );
  XNOR2_X1 U538 ( .A(KEYINPUT32), .B(KEYINPUT65), .ZN(n511) );
  XNOR2_X1 U539 ( .A(n450), .B(n449), .ZN(n692) );
  XNOR2_X1 U540 ( .A(n656), .B(n655), .ZN(G75) );
  NOR2_X1 U541 ( .A1(G237), .A2(G902), .ZN(n417) );
  XOR2_X1 U542 ( .A(KEYINPUT78), .B(n417), .Z(n427) );
  XOR2_X1 U543 ( .A(G113), .B(G104), .Z(n418) );
  XNOR2_X2 U544 ( .A(G128), .B(KEYINPUT83), .ZN(n420) );
  XNOR2_X2 U545 ( .A(n420), .B(G143), .ZN(n456) );
  XOR2_X1 U546 ( .A(KEYINPUT73), .B(G110), .Z(n458) );
  NAND2_X1 U547 ( .A1(G224), .A2(n718), .ZN(n422) );
  XNOR2_X1 U548 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U549 ( .A(n425), .B(KEYINPUT72), .ZN(n702) );
  NAND2_X1 U550 ( .A1(n427), .A2(G214), .ZN(n635) );
  XOR2_X1 U551 ( .A(KEYINPUT80), .B(KEYINPUT19), .Z(n428) );
  XOR2_X1 U552 ( .A(G898), .B(KEYINPUT91), .Z(n697) );
  NOR2_X1 U553 ( .A1(n697), .A2(n718), .ZN(n706) );
  NAND2_X1 U554 ( .A1(n706), .A2(G902), .ZN(n429) );
  NAND2_X1 U555 ( .A1(G952), .A2(n718), .ZN(n546) );
  NAND2_X1 U556 ( .A1(n429), .A2(n546), .ZN(n432) );
  XOR2_X1 U557 ( .A(KEYINPUT77), .B(KEYINPUT14), .Z(n431) );
  XNOR2_X1 U558 ( .A(n431), .B(n430), .ZN(n648) );
  NAND2_X1 U559 ( .A1(n432), .A2(n648), .ZN(n433) );
  INV_X1 U560 ( .A(KEYINPUT0), .ZN(n434) );
  XNOR2_X2 U561 ( .A(n435), .B(n434), .ZN(n526) );
  XNOR2_X1 U562 ( .A(n526), .B(KEYINPUT92), .ZN(n523) );
  XOR2_X1 U563 ( .A(KEYINPUT21), .B(KEYINPUT97), .Z(n438) );
  NAND2_X1 U564 ( .A1(G234), .A2(n598), .ZN(n436) );
  XNOR2_X1 U565 ( .A(KEYINPUT20), .B(n436), .ZN(n451) );
  NAND2_X1 U566 ( .A1(n451), .A2(G221), .ZN(n437) );
  XNOR2_X1 U567 ( .A(n438), .B(n437), .ZN(n618) );
  XOR2_X1 U568 ( .A(n457), .B(n483), .Z(n450) );
  NAND2_X1 U569 ( .A1(G234), .A2(n718), .ZN(n439) );
  NAND2_X1 U570 ( .A1(n487), .A2(G221), .ZN(n448) );
  XOR2_X1 U571 ( .A(KEYINPUT95), .B(KEYINPUT24), .Z(n442) );
  XNOR2_X1 U572 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U573 ( .A(KEYINPUT94), .B(KEYINPUT81), .Z(n444) );
  XNOR2_X1 U574 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U575 ( .A(n446), .B(n445), .Z(n447) );
  NOR2_X1 U576 ( .A1(n692), .A2(G902), .ZN(n455) );
  XOR2_X1 U577 ( .A(KEYINPUT25), .B(KEYINPUT96), .Z(n453) );
  NAND2_X1 U578 ( .A1(G217), .A2(n451), .ZN(n452) );
  XNOR2_X1 U579 ( .A(n453), .B(n452), .ZN(n454) );
  NOR2_X1 U580 ( .A1(n618), .A2(n617), .ZN(n624) );
  NAND2_X1 U581 ( .A1(G227), .A2(n718), .ZN(n459) );
  NAND2_X1 U582 ( .A1(n624), .A2(n623), .ZN(n527) );
  NAND2_X1 U583 ( .A1(n474), .A2(G210), .ZN(n463) );
  XNOR2_X1 U584 ( .A(n464), .B(n463), .ZN(n468) );
  NOR2_X1 U585 ( .A1(n657), .A2(G902), .ZN(n471) );
  XNOR2_X1 U586 ( .A(n472), .B(KEYINPUT33), .ZN(n614) );
  NOR2_X1 U587 ( .A1(n523), .A2(n614), .ZN(n473) );
  XNOR2_X1 U588 ( .A(n473), .B(KEYINPUT34), .ZN(n498) );
  XNOR2_X1 U589 ( .A(KEYINPUT13), .B(G475), .ZN(n486) );
  NAND2_X1 U590 ( .A1(G214), .A2(n474), .ZN(n475) );
  XNOR2_X1 U591 ( .A(n476), .B(n475), .ZN(n480) );
  XNOR2_X1 U592 ( .A(n482), .B(n481), .ZN(n484) );
  XNOR2_X1 U593 ( .A(n483), .B(n484), .ZN(n682) );
  NOR2_X1 U594 ( .A1(G902), .A2(n682), .ZN(n485) );
  XOR2_X1 U595 ( .A(n486), .B(n485), .Z(n533) );
  NAND2_X1 U596 ( .A1(n487), .A2(G217), .ZN(n496) );
  XNOR2_X1 U597 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U598 ( .A(n490), .B(KEYINPUT102), .Z(n494) );
  XNOR2_X1 U599 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U600 ( .A(n496), .B(n495), .ZN(n688) );
  OR2_X1 U601 ( .A1(n533), .A2(n531), .ZN(n564) );
  INV_X1 U602 ( .A(n564), .ZN(n497) );
  INV_X1 U603 ( .A(KEYINPUT87), .ZN(n499) );
  INV_X1 U604 ( .A(KEYINPUT35), .ZN(n500) );
  INV_X1 U605 ( .A(KEYINPUT67), .ZN(n520) );
  XNOR2_X1 U606 ( .A(n728), .B(n520), .ZN(n515) );
  INV_X1 U607 ( .A(KEYINPUT44), .ZN(n513) );
  NAND2_X1 U608 ( .A1(n533), .A2(n531), .ZN(n638) );
  NOR2_X1 U609 ( .A1(n618), .A2(n638), .ZN(n501) );
  XNOR2_X1 U610 ( .A(n501), .B(KEYINPUT103), .ZN(n502) );
  INV_X1 U611 ( .A(n617), .ZN(n508) );
  NOR2_X1 U612 ( .A1(n508), .A2(n507), .ZN(n510) );
  XOR2_X1 U613 ( .A(n623), .B(KEYINPUT90), .Z(n572) );
  NOR2_X1 U614 ( .A1(n572), .A2(n568), .ZN(n509) );
  NAND2_X1 U615 ( .A1(n510), .A2(n509), .ZN(n512) );
  NAND2_X1 U616 ( .A1(n515), .A2(n514), .ZN(n518) );
  INV_X1 U617 ( .A(n519), .ZN(n516) );
  NAND2_X1 U618 ( .A1(n518), .A2(n517), .ZN(n544) );
  NAND2_X1 U619 ( .A1(n520), .A2(n519), .ZN(n522) );
  AND2_X1 U620 ( .A1(KEYINPUT64), .A2(KEYINPUT44), .ZN(n521) );
  NAND2_X1 U621 ( .A1(n522), .A2(n521), .ZN(n542) );
  INV_X1 U622 ( .A(n550), .ZN(n621) );
  NOR2_X1 U623 ( .A1(n621), .A2(n523), .ZN(n525) );
  NAND2_X1 U624 ( .A1(n624), .A2(n554), .ZN(n524) );
  NAND2_X1 U625 ( .A1(n525), .A2(n582), .ZN(n661) );
  INV_X1 U626 ( .A(n526), .ZN(n528) );
  NOR2_X1 U627 ( .A1(n550), .A2(n527), .ZN(n630) );
  NAND2_X1 U628 ( .A1(n528), .A2(n630), .ZN(n529) );
  NAND2_X1 U629 ( .A1(n661), .A2(n676), .ZN(n535) );
  NAND2_X1 U630 ( .A1(n532), .A2(n533), .ZN(n677) );
  INV_X1 U631 ( .A(n349), .ZN(n674) );
  NAND2_X1 U632 ( .A1(n677), .A2(n674), .ZN(n556) );
  INV_X1 U633 ( .A(n556), .ZN(n640) );
  XOR2_X1 U634 ( .A(n640), .B(KEYINPUT85), .Z(n574) );
  INV_X1 U635 ( .A(n574), .ZN(n534) );
  NAND2_X1 U636 ( .A1(n535), .A2(n534), .ZN(n540) );
  NOR2_X1 U637 ( .A1(n617), .A2(n537), .ZN(n659) );
  NOR2_X1 U638 ( .A1(KEYINPUT64), .A2(KEYINPUT44), .ZN(n538) );
  NOR2_X1 U639 ( .A1(n659), .A2(n538), .ZN(n539) );
  NAND2_X1 U640 ( .A1(n542), .A2(n352), .ZN(n543) );
  NOR2_X1 U641 ( .A1(G900), .A2(n718), .ZN(n545) );
  NAND2_X1 U642 ( .A1(n545), .A2(G902), .ZN(n547) );
  NAND2_X1 U643 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U644 ( .A1(n548), .A2(n648), .ZN(n560) );
  NOR2_X1 U645 ( .A1(n618), .A2(n560), .ZN(n549) );
  NOR2_X1 U646 ( .A1(n550), .A2(n566), .ZN(n552) );
  XNOR2_X1 U647 ( .A(KEYINPUT28), .B(KEYINPUT106), .ZN(n551) );
  XNOR2_X1 U648 ( .A(n552), .B(n551), .ZN(n553) );
  NAND2_X1 U649 ( .A1(n556), .A2(n672), .ZN(n557) );
  NAND2_X1 U650 ( .A1(n557), .A2(KEYINPUT47), .ZN(n573) );
  INV_X1 U651 ( .A(n592), .ZN(n578) );
  NAND2_X1 U652 ( .A1(n621), .A2(n635), .ZN(n558) );
  XNOR2_X1 U653 ( .A(KEYINPUT30), .B(n558), .ZN(n559) );
  NOR2_X1 U654 ( .A1(n560), .A2(n559), .ZN(n580) );
  NAND2_X1 U655 ( .A1(n582), .A2(n580), .ZN(n561) );
  NOR2_X1 U656 ( .A1(n578), .A2(n561), .ZN(n562) );
  XNOR2_X1 U657 ( .A(n562), .B(KEYINPUT105), .ZN(n563) );
  XNOR2_X1 U658 ( .A(KEYINPUT108), .B(n587), .ZN(n569) );
  NOR2_X1 U659 ( .A1(n565), .A2(n569), .ZN(n570) );
  XOR2_X1 U660 ( .A(KEYINPUT36), .B(n570), .Z(n571) );
  NOR2_X1 U661 ( .A1(KEYINPUT47), .A2(n574), .ZN(n575) );
  NAND2_X1 U662 ( .A1(n672), .A2(n575), .ZN(n576) );
  XOR2_X1 U663 ( .A(KEYINPUT76), .B(n576), .Z(n577) );
  XNOR2_X1 U664 ( .A(KEYINPUT38), .B(n578), .ZN(n636) );
  NAND2_X1 U665 ( .A1(n636), .A2(n635), .ZN(n639) );
  NOR2_X1 U666 ( .A1(n639), .A2(n638), .ZN(n579) );
  XNOR2_X1 U667 ( .A(n579), .B(KEYINPUT41), .ZN(n634) );
  XNOR2_X1 U668 ( .A(n353), .B(KEYINPUT42), .ZN(n730) );
  INV_X1 U669 ( .A(KEYINPUT40), .ZN(n584) );
  AND2_X1 U670 ( .A1(n580), .A2(n636), .ZN(n581) );
  XNOR2_X1 U671 ( .A(n585), .B(KEYINPUT46), .ZN(n586) );
  XOR2_X1 U672 ( .A(KEYINPUT104), .B(KEYINPUT43), .Z(n590) );
  NOR2_X1 U673 ( .A1(n623), .A2(n587), .ZN(n588) );
  NAND2_X1 U674 ( .A1(n588), .A2(n635), .ZN(n589) );
  XNOR2_X1 U675 ( .A(n590), .B(n589), .ZN(n591) );
  NOR2_X1 U676 ( .A1(n592), .A2(n591), .ZN(n681) );
  INV_X1 U677 ( .A(n677), .ZN(n666) );
  NAND2_X1 U678 ( .A1(n666), .A2(n595), .ZN(n596) );
  XOR2_X1 U679 ( .A(KEYINPUT109), .B(n596), .Z(n727) );
  NOR2_X1 U680 ( .A1(n597), .A2(KEYINPUT2), .ZN(n613) );
  INV_X1 U681 ( .A(n598), .ZN(n599) );
  NAND2_X1 U682 ( .A1(n612), .A2(n599), .ZN(n600) );
  NAND2_X1 U683 ( .A1(n690), .A2(G469), .ZN(n605) );
  XOR2_X1 U684 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n603) );
  XNOR2_X1 U685 ( .A(n601), .B(KEYINPUT119), .ZN(n602) );
  XNOR2_X1 U686 ( .A(n603), .B(n602), .ZN(n604) );
  NAND2_X1 U687 ( .A1(n686), .A2(G210), .ZN(n611) );
  BUF_X1 U688 ( .A(n607), .Z(n608) );
  XOR2_X1 U689 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n609) );
  NAND2_X1 U690 ( .A1(n612), .A2(n348), .ZN(n654) );
  NOR2_X1 U691 ( .A1(n634), .A2(n614), .ZN(n615) );
  XOR2_X1 U692 ( .A(KEYINPUT116), .B(n615), .Z(n616) );
  NAND2_X1 U693 ( .A1(n718), .A2(n616), .ZN(n652) );
  NAND2_X1 U694 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U695 ( .A(KEYINPUT49), .B(n619), .ZN(n620) );
  NOR2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U697 ( .A(KEYINPUT112), .B(n622), .Z(n628) );
  NOR2_X1 U698 ( .A1(n624), .A2(n623), .ZN(n625) );
  XOR2_X1 U699 ( .A(KEYINPUT113), .B(n625), .Z(n626) );
  XNOR2_X1 U700 ( .A(KEYINPUT50), .B(n626), .ZN(n627) );
  NOR2_X1 U701 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U702 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U703 ( .A(KEYINPUT114), .B(n631), .Z(n632) );
  XNOR2_X1 U704 ( .A(n632), .B(KEYINPUT51), .ZN(n633) );
  NOR2_X1 U705 ( .A1(n634), .A2(n633), .ZN(n646) );
  NOR2_X1 U706 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U707 ( .A1(n638), .A2(n637), .ZN(n642) );
  NOR2_X1 U708 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U709 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U710 ( .A1(n643), .A2(n614), .ZN(n644) );
  XOR2_X1 U711 ( .A(KEYINPUT115), .B(n644), .Z(n645) );
  NOR2_X1 U712 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U713 ( .A(KEYINPUT52), .B(n647), .ZN(n650) );
  NAND2_X1 U714 ( .A1(n648), .A2(G952), .ZN(n649) );
  NOR2_X1 U715 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U716 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U717 ( .A1(n654), .A2(n653), .ZN(n656) );
  XNOR2_X1 U718 ( .A(KEYINPUT117), .B(KEYINPUT53), .ZN(n655) );
  NAND2_X1 U719 ( .A1(n686), .A2(G472), .ZN(n658) );
  XOR2_X1 U720 ( .A(G101), .B(n659), .Z(G3) );
  NOR2_X1 U721 ( .A1(n674), .A2(n661), .ZN(n660) );
  XOR2_X1 U722 ( .A(G104), .B(n660), .Z(G6) );
  NOR2_X1 U723 ( .A1(n677), .A2(n661), .ZN(n663) );
  XNOR2_X1 U724 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n662) );
  XNOR2_X1 U725 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U726 ( .A(G107), .B(n664), .ZN(G9) );
  XOR2_X1 U727 ( .A(n665), .B(G110), .Z(G12) );
  XOR2_X1 U728 ( .A(KEYINPUT29), .B(KEYINPUT110), .Z(n668) );
  NAND2_X1 U729 ( .A1(n347), .A2(n666), .ZN(n667) );
  XNOR2_X1 U730 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U731 ( .A(G128), .B(n669), .ZN(G30) );
  XNOR2_X1 U732 ( .A(G143), .B(n670), .ZN(n671) );
  XNOR2_X1 U733 ( .A(n671), .B(KEYINPUT111), .ZN(G45) );
  NAND2_X1 U734 ( .A1(n349), .A2(n347), .ZN(n673) );
  XNOR2_X1 U735 ( .A(G146), .B(n673), .ZN(G48) );
  NOR2_X1 U736 ( .A1(n674), .A2(n676), .ZN(n675) );
  XOR2_X1 U737 ( .A(G113), .B(n675), .Z(G15) );
  NOR2_X1 U738 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U739 ( .A(G116), .B(n678), .Z(G18) );
  XNOR2_X1 U740 ( .A(G125), .B(n679), .ZN(n680) );
  XNOR2_X1 U741 ( .A(n680), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U742 ( .A(G140), .B(n681), .Z(G42) );
  NAND2_X1 U743 ( .A1(n686), .A2(G475), .ZN(n683) );
  NAND2_X1 U744 ( .A1(n690), .A2(G478), .ZN(n687) );
  NOR2_X1 U745 ( .A1(n694), .A2(n689), .ZN(G63) );
  NAND2_X1 U746 ( .A1(G217), .A2(n690), .ZN(n691) );
  XNOR2_X1 U747 ( .A(n692), .B(n691), .ZN(n693) );
  NOR2_X1 U748 ( .A1(n694), .A2(n693), .ZN(G66) );
  OR2_X1 U749 ( .A1(G953), .A2(n695), .ZN(n700) );
  NAND2_X1 U750 ( .A1(G953), .A2(G224), .ZN(n696) );
  XNOR2_X1 U751 ( .A(KEYINPUT61), .B(n696), .ZN(n698) );
  NAND2_X1 U752 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U753 ( .A1(n700), .A2(n699), .ZN(n708) );
  XNOR2_X1 U754 ( .A(n701), .B(n702), .ZN(n703) );
  XNOR2_X1 U755 ( .A(n703), .B(G110), .ZN(n704) );
  XNOR2_X1 U756 ( .A(n704), .B(G101), .ZN(n705) );
  NOR2_X1 U757 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U758 ( .A(n708), .B(n707), .ZN(n710) );
  XOR2_X1 U759 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n709) );
  XNOR2_X1 U760 ( .A(n710), .B(n709), .ZN(G69) );
  XNOR2_X1 U761 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n714) );
  XNOR2_X1 U762 ( .A(n712), .B(n711), .ZN(n713) );
  XNOR2_X1 U763 ( .A(n714), .B(n713), .ZN(n716) );
  XNOR2_X1 U764 ( .A(n715), .B(n716), .ZN(n720) );
  XOR2_X1 U765 ( .A(n720), .B(n717), .Z(n719) );
  NAND2_X1 U766 ( .A1(n719), .A2(n718), .ZN(n726) );
  XNOR2_X1 U767 ( .A(G227), .B(n720), .ZN(n721) );
  XNOR2_X1 U768 ( .A(n721), .B(KEYINPUT125), .ZN(n722) );
  NAND2_X1 U769 ( .A1(G900), .A2(n722), .ZN(n723) );
  XNOR2_X1 U770 ( .A(KEYINPUT126), .B(n723), .ZN(n724) );
  NAND2_X1 U771 ( .A1(n724), .A2(G953), .ZN(n725) );
  NAND2_X1 U772 ( .A1(n726), .A2(n725), .ZN(G72) );
  XNOR2_X1 U773 ( .A(G134), .B(n727), .ZN(G36) );
  XNOR2_X1 U774 ( .A(n728), .B(G122), .ZN(G24) );
  XOR2_X1 U775 ( .A(n729), .B(G131), .Z(G33) );
  XOR2_X1 U776 ( .A(G137), .B(n730), .Z(G39) );
  BUF_X1 U777 ( .A(n731), .Z(n732) );
  XOR2_X1 U778 ( .A(G119), .B(n732), .Z(G21) );
endmodule

