//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 1 0 0 0 1 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 0 0 0 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n794, new_n795, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982, new_n983;
  INV_X1    g000(.A(G50gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(G43gat), .ZN(new_n203));
  INV_X1    g002(.A(G43gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n204), .A2(G50gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT15), .ZN(new_n206));
  NOR3_X1   g005(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  OR3_X1    g007(.A1(new_n202), .A2(KEYINPUT85), .A3(G43gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT85), .B1(new_n204), .B2(G50gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n209), .B(new_n206), .C1(new_n203), .C2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT83), .B1(G29gat), .B2(G36gat), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n213), .A2(KEYINPUT14), .ZN(new_n214));
  NAND2_X1  g013(.A1(G29gat), .A2(G36gat), .ZN(new_n215));
  NOR3_X1   g014(.A1(KEYINPUT83), .A2(G29gat), .A3(G36gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(KEYINPUT14), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n214), .B(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n212), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n207), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n220), .A2(KEYINPUT84), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n220), .A2(KEYINPUT84), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n219), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n223), .B(KEYINPUT17), .ZN(new_n224));
  XNOR2_X1  g023(.A(G15gat), .B(G22gat), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n225), .A2(G1gat), .ZN(new_n226));
  AOI21_X1  g025(.A(G8gat), .B1(new_n226), .B2(KEYINPUT86), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT16), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n225), .B1(new_n228), .B2(G1gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n227), .B(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n224), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G229gat), .A2(G233gat), .ZN(new_n233));
  INV_X1    g032(.A(new_n231), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(new_n223), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n232), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT18), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n232), .A2(KEYINPUT18), .A3(new_n233), .A4(new_n235), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n234), .B(new_n223), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n233), .B(KEYINPUT13), .Z(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n238), .A2(new_n239), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G113gat), .B(G141gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(G169gat), .B(G197gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n248), .B(KEYINPUT12), .Z(new_n249));
  NAND2_X1  g048(.A1(new_n243), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n249), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n238), .A2(new_n239), .A3(new_n242), .A4(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT80), .ZN(new_n255));
  INV_X1    g054(.A(G155gat), .ZN(new_n256));
  INV_X1    g055(.A(G162gat), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT74), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G141gat), .B(G148gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT2), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n260), .B1(G155gat), .B2(G162gat), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n258), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(G155gat), .B(G162gat), .Z(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT29), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OR2_X1    g065(.A1(new_n266), .A2(KEYINPUT78), .ZN(new_n267));
  NAND2_X1  g066(.A1(G211gat), .A2(G218gat), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT22), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G197gat), .ZN(new_n271));
  INV_X1    g070(.A(G204gat), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(G197gat), .A2(G204gat), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n270), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n275), .A2(KEYINPUT70), .ZN(new_n276));
  XOR2_X1   g075(.A(G211gat), .B(G218gat), .Z(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  OR2_X1    g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n276), .A2(new_n278), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT78), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n267), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G228gat), .A2(G233gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT3), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n285), .B1(new_n281), .B2(KEYINPUT29), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n262), .A2(new_n263), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n262), .A2(new_n263), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT75), .ZN(new_n289));
  OR3_X1    g088(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n264), .A2(new_n289), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n284), .B1(new_n286), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n283), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n265), .ZN(new_n295));
  OR2_X1    g094(.A1(new_n278), .A2(new_n275), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT29), .B1(new_n278), .B2(new_n275), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OR3_X1    g097(.A1(new_n298), .A2(new_n264), .A3(KEYINPUT77), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT77), .B1(new_n298), .B2(new_n264), .ZN(new_n300));
  INV_X1    g099(.A(new_n281), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n299), .B(new_n300), .C1(new_n301), .C2(new_n266), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(new_n284), .ZN(new_n303));
  INV_X1    g102(.A(G22gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n294), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT79), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n304), .B1(new_n294), .B2(new_n303), .ZN(new_n308));
  OR3_X1    g107(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n307), .B1(new_n306), .B2(new_n308), .ZN(new_n310));
  XNOR2_X1  g109(.A(G78gat), .B(G106gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n311), .B(KEYINPUT31), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n312), .B(G50gat), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n309), .A2(new_n310), .A3(new_n314), .ZN(new_n315));
  OR2_X1    g114(.A1(new_n310), .A2(new_n314), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  XOR2_X1   g117(.A(G113gat), .B(G120gat), .Z(new_n319));
  INV_X1    g118(.A(KEYINPUT1), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n321), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n322));
  INV_X1    g121(.A(G134gat), .ZN(new_n323));
  INV_X1    g122(.A(G127gat), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n319), .A2(new_n320), .A3(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n322), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n323), .B1(new_n322), .B2(new_n325), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n264), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT4), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n328), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(new_n326), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n333), .A2(KEYINPUT4), .A3(new_n264), .ZN(new_n334));
  AND2_X1   g133(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n285), .B1(new_n290), .B2(new_n291), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n264), .A2(new_n265), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n337), .A2(new_n332), .A3(new_n326), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G225gat), .A2(G233gat), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n335), .A2(new_n340), .A3(KEYINPUT5), .A4(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n331), .A2(new_n334), .ZN(new_n343));
  INV_X1    g142(.A(new_n341), .ZN(new_n344));
  NOR3_X1   g143(.A1(new_n343), .A2(new_n339), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT5), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n327), .A2(new_n328), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n292), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(new_n329), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n346), .B1(new_n349), .B2(new_n344), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n342), .B1(new_n345), .B2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G1gat), .B(G29gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT0), .ZN(new_n353));
  XNOR2_X1  g152(.A(G57gat), .B(G85gat), .ZN(new_n354));
  XOR2_X1   g153(.A(new_n353), .B(new_n354), .Z(new_n355));
  NAND2_X1  g154(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT6), .ZN(new_n357));
  INV_X1    g156(.A(new_n355), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n342), .B(new_n358), .C1(new_n345), .C2(new_n350), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n356), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  OR3_X1    g159(.A1(new_n351), .A2(new_n357), .A3(new_n355), .ZN(new_n361));
  AND2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT30), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT29), .ZN(new_n364));
  AND2_X1   g163(.A1(G169gat), .A2(G176gat), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT26), .ZN(new_n366));
  NOR2_X1   g165(.A1(G169gat), .A2(G176gat), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n368), .A2(new_n369), .B1(G183gat), .B2(G190gat), .ZN(new_n370));
  INV_X1    g169(.A(G183gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT27), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT27), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(G183gat), .ZN(new_n374));
  INV_X1    g173(.A(G190gat), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n372), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT28), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT65), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n376), .A2(KEYINPUT65), .A3(new_n377), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n373), .A2(G183gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n371), .A2(KEYINPUT27), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT66), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT66), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n372), .A2(new_n374), .A3(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n377), .A2(G190gat), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n385), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT67), .B1(new_n382), .B2(new_n389), .ZN(new_n390));
  AND3_X1   g189(.A1(new_n376), .A2(KEYINPUT65), .A3(new_n377), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT65), .B1(new_n376), .B2(new_n377), .ZN(new_n392));
  OAI211_X1 g191(.A(KEYINPUT67), .B(new_n389), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  OAI211_X1 g193(.A(KEYINPUT68), .B(new_n370), .C1(new_n390), .C2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n396), .B1(new_n371), .B2(new_n375), .ZN(new_n397));
  NAND3_X1  g196(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT23), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n367), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n365), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT25), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT64), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n399), .A2(new_n403), .A3(KEYINPUT25), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n407), .B1(new_n406), .B2(new_n408), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n370), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n389), .B1(new_n391), .B2(new_n392), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT67), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n413), .B1(new_n416), .B2(new_n393), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n417), .A2(KEYINPUT68), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n364), .B1(new_n412), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G226gat), .A2(G233gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n370), .B1(new_n390), .B2(new_n394), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n408), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(KEYINPUT71), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT71), .ZN(new_n425));
  INV_X1    g224(.A(new_n423), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n425), .B1(new_n417), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n420), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n424), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT72), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT72), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n424), .A2(new_n427), .A3(new_n431), .A4(new_n428), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n421), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n281), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT73), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT73), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n433), .A2(new_n436), .A3(new_n281), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT68), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n439), .A2(new_n428), .A3(new_n395), .A4(new_n411), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n427), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n420), .A2(new_n364), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n301), .ZN(new_n444));
  XNOR2_X1  g243(.A(G8gat), .B(G36gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(G64gat), .B(G92gat), .ZN(new_n446));
  XOR2_X1   g245(.A(new_n445), .B(new_n446), .Z(new_n447));
  NAND4_X1  g246(.A1(new_n435), .A2(new_n437), .A3(new_n444), .A4(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n362), .B1(new_n363), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n447), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n420), .A2(new_n419), .B1(new_n429), .B2(KEYINPUT72), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n301), .B1(new_n451), .B2(new_n432), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n444), .B1(new_n452), .B2(new_n436), .ZN(new_n453));
  INV_X1    g252(.A(new_n437), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n450), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n434), .A2(KEYINPUT73), .B1(new_n301), .B2(new_n443), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n456), .A2(KEYINPUT30), .A3(new_n437), .A4(new_n447), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n318), .B1(new_n449), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT36), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n333), .B1(new_n412), .B2(new_n418), .ZN(new_n461));
  INV_X1    g260(.A(G227gat), .ZN(new_n462));
  INV_X1    g261(.A(G233gat), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n439), .A2(new_n347), .A3(new_n395), .A4(new_n411), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n461), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT33), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  XOR2_X1   g267(.A(G15gat), .B(G43gat), .Z(new_n469));
  XNOR2_X1  g268(.A(G71gat), .B(G99gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  AOI211_X1 g271(.A(KEYINPUT34), .B(new_n464), .C1(new_n461), .C2(new_n465), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n461), .A2(new_n465), .ZN(new_n475));
  INV_X1    g274(.A(new_n464), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT34), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n472), .A2(new_n474), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n466), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT32), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n471), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n483), .B1(new_n466), .B2(new_n467), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT34), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n485), .B1(new_n475), .B2(new_n476), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n484), .B1(new_n486), .B2(new_n473), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n479), .A2(new_n482), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n482), .B1(new_n479), .B2(new_n487), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n460), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n487), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n484), .A2(new_n486), .A3(new_n473), .ZN(new_n492));
  OAI22_X1  g291(.A1(new_n491), .A2(new_n492), .B1(new_n481), .B2(new_n480), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n479), .A2(new_n482), .A3(new_n487), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(KEYINPUT36), .A3(new_n494), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n255), .B1(new_n459), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n448), .A2(new_n363), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n360), .A2(new_n361), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n498), .A2(new_n499), .A3(new_n455), .A4(new_n457), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n317), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n490), .A2(new_n495), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(KEYINPUT80), .A3(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(KEYINPUT81), .B(KEYINPUT37), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n435), .A2(new_n437), .A3(new_n444), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n450), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT37), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n507), .B1(new_n456), .B2(new_n437), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT38), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n433), .A2(new_n301), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n507), .B1(new_n443), .B2(new_n281), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT38), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n505), .A2(new_n450), .A3(new_n512), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n509), .A2(new_n513), .A3(new_n362), .A4(new_n448), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n455), .A3(new_n457), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n344), .B1(new_n343), .B2(new_n339), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n516), .B(KEYINPUT39), .C1(new_n344), .C2(new_n349), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n517), .B(new_n355), .C1(KEYINPUT39), .C2(new_n516), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT40), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n519), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n520), .A2(new_n359), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n317), .B1(new_n515), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n514), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n497), .A2(new_n503), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT35), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n488), .A2(new_n489), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n318), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n526), .B1(new_n528), .B2(new_n500), .ZN(new_n529));
  NOR3_X1   g328(.A1(new_n317), .A2(new_n488), .A3(new_n489), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n530), .A2(new_n449), .A3(new_n458), .A4(KEYINPUT35), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n254), .B1(new_n525), .B2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G231gat), .A2(G233gat), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(G71gat), .A2(G78gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(G71gat), .A2(G78gat), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n543), .B1(KEYINPUT87), .B2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G57gat), .B(G64gat), .ZN(new_n546));
  NOR2_X1   g345(.A1(KEYINPUT87), .A2(KEYINPUT9), .ZN(new_n547));
  OAI221_X1 g346(.A(new_n545), .B1(KEYINPUT87), .B2(new_n544), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(KEYINPUT89), .A2(G57gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT88), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n549), .A2(new_n550), .A3(G64gat), .ZN(new_n551));
  INV_X1    g350(.A(G64gat), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT88), .B1(new_n552), .B2(G57gat), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n551), .B(new_n553), .C1(G64gat), .C2(new_n549), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT90), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n543), .A2(KEYINPUT9), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(new_n544), .ZN(new_n557));
  AND3_X1   g356(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n555), .B1(new_n554), .B2(new_n557), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n548), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT91), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT91), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n562), .B(new_n548), .C1(new_n558), .C2(new_n559), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n542), .B1(new_n564), .B2(KEYINPUT21), .ZN(new_n565));
  XNOR2_X1  g364(.A(G127gat), .B(G155gat), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n566), .B(KEYINPUT92), .Z(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT21), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n561), .A2(new_n569), .A3(new_n563), .A4(new_n541), .ZN(new_n570));
  AND3_X1   g369(.A1(new_n565), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n568), .B1(new_n565), .B2(new_n570), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n540), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n565), .A2(new_n570), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(new_n567), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n565), .A2(new_n568), .A3(new_n570), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n575), .A2(new_n539), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n564), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n231), .B1(new_n578), .B2(new_n569), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n573), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n579), .B1(new_n573), .B2(new_n577), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n538), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n579), .ZN(new_n583));
  NOR3_X1   g382(.A1(new_n571), .A2(new_n572), .A3(new_n540), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n539), .B1(new_n575), .B2(new_n576), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n573), .A2(new_n577), .A3(new_n579), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(new_n537), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G183gat), .B(G211gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n582), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n590), .B1(new_n582), .B2(new_n588), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n536), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT100), .ZN(new_n594));
  NAND2_X1  g393(.A1(G99gat), .A2(G106gat), .ZN(new_n595));
  INV_X1    g394(.A(G85gat), .ZN(new_n596));
  INV_X1    g395(.A(G92gat), .ZN(new_n597));
  AOI22_X1  g396(.A1(KEYINPUT8), .A2(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT98), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT97), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n600), .A2(G85gat), .A3(G92gat), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n601), .B(KEYINPUT7), .Z(new_n602));
  OAI21_X1  g401(.A(KEYINPUT99), .B1(new_n599), .B2(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(G99gat), .B(G106gat), .Z(new_n604));
  INV_X1    g403(.A(KEYINPUT98), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n598), .B(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT99), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n601), .B(KEYINPUT7), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n603), .A2(new_n604), .A3(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n604), .B1(new_n603), .B2(new_n609), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n594), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n604), .ZN(new_n614));
  NOR3_X1   g413(.A1(new_n599), .A2(new_n602), .A3(KEYINPUT99), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n607), .B1(new_n606), .B2(new_n608), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n617), .A2(KEYINPUT100), .A3(new_n610), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n221), .A2(new_n222), .ZN(new_n619));
  AOI22_X1  g418(.A1(new_n613), .A2(new_n618), .B1(new_n619), .B2(new_n219), .ZN(new_n620));
  NAND2_X1  g419(.A1(G232gat), .A2(G233gat), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT41), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(KEYINPUT101), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  NOR3_X1   g423(.A1(new_n611), .A2(new_n594), .A3(new_n612), .ZN(new_n625));
  AOI21_X1  g424(.A(KEYINPUT100), .B1(new_n617), .B2(new_n610), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n223), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT101), .ZN(new_n628));
  INV_X1    g427(.A(new_n623), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n625), .A2(new_n626), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n224), .ZN(new_n633));
  XNOR2_X1  g432(.A(G190gat), .B(G218gat), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n631), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G134gat), .B(G162gat), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  AOI22_X1  g440(.A1(new_n624), .A2(new_n630), .B1(new_n224), .B2(new_n632), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(new_n635), .ZN(new_n643));
  OAI21_X1  g442(.A(KEYINPUT103), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n631), .A2(new_n633), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n634), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT103), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n646), .A2(new_n647), .A3(new_n636), .A4(new_n640), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT102), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n642), .A2(new_n650), .A3(new_n635), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(new_n639), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n643), .A2(new_n650), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n652), .B1(new_n653), .B2(new_n636), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(G230gat), .A2(G233gat), .ZN(new_n656));
  INV_X1    g455(.A(new_n560), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n657), .B1(new_n611), .B2(new_n612), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n617), .A2(new_n561), .A3(new_n563), .A4(new_n610), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT104), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n578), .A2(KEYINPUT104), .A3(new_n610), .A4(new_n617), .ZN(new_n662));
  AOI21_X1  g461(.A(KEYINPUT10), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n564), .A2(KEYINPUT10), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n632), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n656), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(G120gat), .B(G148gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(G176gat), .B(G204gat), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n667), .B(new_n668), .Z(new_n669));
  NAND2_X1  g468(.A1(new_n661), .A2(new_n662), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n670), .A2(new_n656), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n666), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT106), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n656), .B(KEYINPUT105), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n676), .B1(new_n663), .B2(new_n665), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n671), .ZN(new_n678));
  INV_X1    g477(.A(new_n669), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n674), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n678), .A2(new_n674), .A3(new_n679), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n673), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n580), .A2(new_n581), .A3(new_n538), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n537), .B1(new_n586), .B2(new_n587), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n589), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n582), .A2(new_n588), .A3(new_n590), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n686), .A2(new_n535), .A3(new_n687), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n593), .A2(new_n655), .A3(new_n683), .A4(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n534), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n362), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(G1gat), .ZN(G1324gat));
  INV_X1    g493(.A(new_n515), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT16), .B(G8gat), .Z(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT42), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n692), .A2(new_n515), .ZN(new_n700));
  AOI22_X1  g499(.A1(new_n698), .A2(new_n699), .B1(new_n700), .B2(G8gat), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(new_n699), .B2(new_n698), .ZN(G1325gat));
  XNOR2_X1  g501(.A(new_n502), .B(KEYINPUT107), .ZN(new_n703));
  OAI21_X1  g502(.A(G15gat), .B1(new_n691), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n527), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n705), .A2(G15gat), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n704), .B1(new_n691), .B2(new_n706), .ZN(G1326gat));
  OR3_X1    g506(.A1(new_n691), .A2(KEYINPUT108), .A3(new_n318), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT108), .B1(new_n691), .B2(new_n318), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT43), .B(G22gat), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n710), .B(new_n712), .ZN(G1327gat));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n500), .A2(KEYINPUT110), .A3(new_n317), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT110), .B1(new_n500), .B2(new_n317), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n715), .A2(new_n716), .A3(new_n496), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n532), .B1(new_n717), .B2(new_n524), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n714), .B1(new_n718), .B2(new_n655), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n525), .A2(new_n533), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n655), .A2(new_n714), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n593), .A2(KEYINPUT109), .A3(new_n688), .ZN(new_n724));
  AOI21_X1  g523(.A(KEYINPUT109), .B1(new_n593), .B2(new_n688), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n682), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n672), .B1(new_n727), .B2(new_n680), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n726), .A2(new_n254), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n723), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(G29gat), .B1(new_n730), .B2(new_n499), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n593), .A2(new_n688), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n733), .A2(new_n655), .A3(new_n728), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n499), .A2(G29gat), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n534), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT45), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n731), .A2(new_n737), .ZN(G1328gat));
  OAI21_X1  g537(.A(G36gat), .B1(new_n730), .B2(new_n695), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n695), .A2(G36gat), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n534), .A2(new_n734), .A3(new_n740), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(KEYINPUT46), .Z(new_n742));
  NAND2_X1  g541(.A1(new_n739), .A2(new_n742), .ZN(G1329gat));
  NAND3_X1  g542(.A1(new_n723), .A2(new_n496), .A3(new_n729), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(G43gat), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT47), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n705), .A2(G43gat), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n534), .A2(new_n734), .A3(new_n747), .ZN(new_n748));
  OR2_X1    g547(.A1(new_n748), .A2(KEYINPUT111), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(KEYINPUT111), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n746), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n745), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n703), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n723), .A2(new_n753), .A3(new_n729), .ZN(new_n754));
  AOI22_X1  g553(.A1(new_n754), .A2(G43gat), .B1(new_n750), .B2(new_n749), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n752), .B1(new_n755), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g555(.A(KEYINPUT113), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n719), .A2(new_n317), .A3(new_n722), .A4(new_n729), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n757), .B1(new_n758), .B2(G50gat), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n317), .A2(new_n202), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(KEYINPUT112), .Z(new_n761));
  AND3_X1   g560(.A1(new_n534), .A2(new_n734), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n762), .B1(new_n758), .B2(G50gat), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT48), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n759), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  AOI221_X4 g564(.A(new_n762), .B1(new_n757), .B2(KEYINPUT48), .C1(new_n758), .C2(G50gat), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(G1331gat));
  NOR2_X1   g566(.A1(new_n716), .A2(new_n496), .ZN(new_n768));
  INV_X1    g567(.A(new_n715), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n768), .A2(new_n769), .A3(new_n524), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n533), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n646), .A2(KEYINPUT102), .A3(new_n636), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n644), .B(new_n648), .C1(new_n772), .C2(new_n652), .ZN(new_n773));
  NOR4_X1   g572(.A1(new_n732), .A2(new_n253), .A3(new_n773), .A4(new_n683), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n362), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g577(.A1(new_n775), .A2(new_n695), .ZN(new_n779));
  NOR2_X1   g578(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n780));
  AND2_X1   g579(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n782), .B1(new_n779), .B2(new_n780), .ZN(G1333gat));
  NAND3_X1  g582(.A1(new_n776), .A2(G71gat), .A3(new_n753), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n775), .A2(new_n705), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n785), .A2(KEYINPUT114), .ZN(new_n786));
  INV_X1    g585(.A(G71gat), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(new_n785), .B2(KEYINPUT114), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n784), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT50), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n791), .B(new_n784), .C1(new_n786), .C2(new_n788), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(G1334gat));
  NOR2_X1   g592(.A1(new_n775), .A2(new_n318), .ZN(new_n794));
  XNOR2_X1  g593(.A(KEYINPUT115), .B(G78gat), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n794), .B(new_n795), .ZN(G1335gat));
  NAND3_X1  g595(.A1(new_n732), .A2(new_n254), .A3(new_n728), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n719), .A2(new_n722), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(G85gat), .B1(new_n800), .B2(new_n499), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n655), .B1(new_n770), .B2(new_n533), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n733), .A2(new_n253), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT51), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n802), .A2(KEYINPUT51), .A3(new_n803), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n807), .A2(new_n596), .A3(new_n362), .A4(new_n728), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n801), .A2(new_n808), .ZN(G1336gat));
  NAND2_X1  g608(.A1(new_n799), .A2(new_n515), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G92gat), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n515), .A2(new_n597), .A3(new_n728), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(KEYINPUT116), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(new_n805), .B2(new_n806), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n811), .A2(new_n812), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n597), .B1(new_n799), .B2(new_n515), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT52), .B1(new_n819), .B2(new_n816), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(G1337gat));
  OAI21_X1  g620(.A(G99gat), .B1(new_n800), .B2(new_n703), .ZN(new_n822));
  INV_X1    g621(.A(G99gat), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n705), .A2(new_n683), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n807), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n822), .A2(new_n825), .ZN(G1338gat));
  NOR2_X1   g625(.A1(new_n318), .A2(G106gat), .ZN(new_n827));
  INV_X1    g626(.A(new_n806), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n728), .B(new_n827), .C1(new_n828), .C2(new_n804), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT117), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n719), .A2(new_n317), .A3(new_n722), .A4(new_n798), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(G106gat), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n830), .A2(new_n833), .A3(KEYINPUT53), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n829), .B(new_n832), .C1(KEYINPUT117), .C2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(new_n836), .ZN(G1339gat));
  INV_X1    g636(.A(KEYINPUT55), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT10), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n670), .A2(new_n839), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n632), .A2(new_n664), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(new_n841), .A3(new_n675), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n842), .A2(KEYINPUT54), .A3(new_n666), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n844), .B(new_n676), .C1(new_n663), .C2(new_n665), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n679), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n838), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n847), .A2(new_n672), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n233), .B1(new_n232), .B2(new_n235), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n850));
  OAI22_X1  g649(.A1(new_n849), .A2(new_n850), .B1(new_n240), .B2(new_n241), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n849), .A2(new_n850), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n248), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n252), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n842), .A2(new_n666), .A3(KEYINPUT54), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n856), .A2(KEYINPUT55), .A3(new_n679), .A4(new_n845), .ZN(new_n857));
  AND4_X1   g656(.A1(new_n773), .A2(new_n848), .A3(new_n855), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n728), .A2(new_n855), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n847), .A2(new_n253), .A3(new_n672), .A4(new_n857), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n773), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI22_X1  g660(.A1(new_n724), .A2(new_n725), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n690), .A2(new_n254), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n317), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n362), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n865), .A2(new_n515), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n253), .A3(new_n527), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g667(.A1(new_n866), .A2(new_n824), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g669(.A1(new_n866), .A2(new_n527), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n324), .B1(new_n871), .B2(new_n732), .ZN(new_n872));
  INV_X1    g671(.A(new_n726), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(new_n324), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(KEYINPUT119), .B1(new_n871), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n871), .A2(KEYINPUT119), .A3(new_n875), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n877), .A2(new_n878), .ZN(G1342gat));
  NOR2_X1   g678(.A1(new_n655), .A2(new_n515), .ZN(new_n880));
  XOR2_X1   g679(.A(KEYINPUT69), .B(G134gat), .Z(new_n881));
  NAND3_X1  g680(.A1(new_n880), .A2(new_n527), .A3(new_n881), .ZN(new_n882));
  OR3_X1    g681(.A1(new_n865), .A2(KEYINPUT120), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT120), .B1(new_n865), .B2(new_n882), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT56), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(G134gat), .B1(new_n871), .B2(new_n655), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n883), .A2(KEYINPUT56), .A3(new_n884), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(G1343gat));
  NOR2_X1   g689(.A1(new_n515), .A2(new_n499), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n502), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n318), .B1(new_n862), .B2(new_n863), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n689), .A2(new_n253), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n773), .A2(new_n848), .A3(new_n855), .A4(new_n857), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n683), .A2(new_n854), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n847), .A2(new_n857), .A3(new_n672), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n254), .B1(new_n899), .B2(KEYINPUT121), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n847), .A2(new_n857), .A3(new_n901), .A4(new_n672), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n898), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n897), .B1(new_n903), .B2(new_n773), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n896), .B1(new_n904), .B2(new_n732), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT57), .B1(new_n905), .B2(new_n318), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n895), .A2(new_n906), .A3(new_n253), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(G141gat), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n893), .A2(new_n703), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n254), .A2(G141gat), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(new_n891), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n908), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n910), .A2(new_n914), .A3(KEYINPUT58), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT58), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n908), .B(new_n913), .C1(new_n909), .C2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(G1344gat));
  NOR2_X1   g717(.A1(new_n683), .A2(G148gat), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n911), .A2(new_n891), .A3(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n921));
  INV_X1    g720(.A(new_n892), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n904), .A2(new_n732), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(new_n863), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT57), .B1(new_n924), .B2(new_n317), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n893), .A2(KEYINPUT57), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n728), .B(new_n922), .C1(new_n925), .C2(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n921), .B1(new_n927), .B2(G148gat), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n895), .A2(new_n906), .A3(new_n728), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n929), .A2(new_n921), .A3(G148gat), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n920), .B1(new_n928), .B2(new_n930), .ZN(G1345gat));
  NAND2_X1  g730(.A1(new_n895), .A2(new_n906), .ZN(new_n932));
  OAI21_X1  g731(.A(G155gat), .B1(new_n932), .B2(new_n873), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n911), .A2(new_n256), .A3(new_n733), .A4(new_n891), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1346gat));
  OAI21_X1  g734(.A(G162gat), .B1(new_n932), .B2(new_n655), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n911), .A2(new_n257), .A3(new_n362), .A4(new_n880), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1347gat));
  NOR2_X1   g737(.A1(new_n695), .A2(new_n362), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n864), .A2(new_n527), .A3(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT123), .ZN(new_n941));
  OAI22_X1  g740(.A1(new_n940), .A2(new_n254), .B1(new_n941), .B2(G169gat), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(G169gat), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n942), .B(new_n943), .ZN(G1348gat));
  NOR2_X1   g743(.A1(new_n940), .A2(new_n683), .ZN(new_n945));
  XOR2_X1   g744(.A(new_n945), .B(G176gat), .Z(G1349gat));
  OAI21_X1  g745(.A(G183gat), .B1(new_n940), .B2(new_n873), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT124), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n733), .A2(new_n385), .A3(new_n387), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n947), .B(new_n948), .C1(new_n940), .C2(new_n949), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT60), .ZN(G1350gat));
  NOR3_X1   g750(.A1(new_n940), .A2(G190gat), .A3(new_n655), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT125), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n940), .A2(new_n655), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n954), .A2(new_n375), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n955), .A2(KEYINPUT61), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(KEYINPUT61), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n953), .A2(new_n956), .A3(new_n957), .ZN(G1351gat));
  NOR2_X1   g757(.A1(new_n925), .A2(new_n926), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n703), .A2(new_n939), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT126), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n962), .A2(new_n271), .A3(new_n254), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n911), .A2(new_n253), .A3(new_n939), .ZN(new_n964));
  AOI22_X1  g763(.A1(new_n960), .A2(new_n963), .B1(new_n964), .B2(new_n271), .ZN(G1352gat));
  NAND4_X1  g764(.A1(new_n911), .A2(new_n272), .A3(new_n728), .A4(new_n939), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n966), .A2(KEYINPUT62), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(KEYINPUT62), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n959), .A2(new_n683), .A3(new_n962), .ZN(new_n969));
  OAI211_X1 g768(.A(new_n967), .B(new_n968), .C1(new_n969), .C2(new_n272), .ZN(G1353gat));
  INV_X1    g769(.A(G211gat), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT63), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n971), .B1(KEYINPUT127), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n703), .A2(new_n733), .A3(new_n939), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n973), .B1(new_n959), .B2(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n975), .A2(new_n976), .A3(KEYINPUT63), .ZN(new_n977));
  OAI221_X1 g776(.A(new_n973), .B1(KEYINPUT127), .B2(new_n972), .C1(new_n959), .C2(new_n974), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n911), .A2(new_n971), .A3(new_n733), .A4(new_n939), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(G1354gat));
  INV_X1    g779(.A(G218gat), .ZN(new_n981));
  NOR3_X1   g780(.A1(new_n962), .A2(new_n981), .A3(new_n655), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n911), .A2(new_n773), .A3(new_n939), .ZN(new_n983));
  AOI22_X1  g782(.A1(new_n960), .A2(new_n982), .B1(new_n983), .B2(new_n981), .ZN(G1355gat));
endmodule


