//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 0 0 0 1 1 0 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 1 1 0 0 1 0 0 0 0 0 1 1 1 1 0 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991;
  XNOR2_X1  g000(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G50gat), .ZN(new_n203));
  XOR2_X1   g002(.A(G78gat), .B(G106gat), .Z(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  AND2_X1   g004(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n207));
  OAI21_X1  g006(.A(G148gat), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G141gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(G148gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT2), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G155gat), .ZN(new_n216));
  INV_X1    g015(.A(G162gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G148gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(G141gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n214), .B1(new_n210), .B2(new_n220), .ZN(new_n221));
  AND2_X1   g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n222), .A2(new_n213), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n212), .A2(new_n218), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT29), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G197gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT73), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n230), .A2(G204gat), .ZN(new_n231));
  INV_X1    g030(.A(G204gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n232), .A2(KEYINPUT73), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n229), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT22), .ZN(new_n235));
  INV_X1    g034(.A(G211gat), .ZN(new_n236));
  INV_X1    g035(.A(G218gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n232), .A2(KEYINPUT73), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n230), .A2(G204gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(new_n240), .A3(G197gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n234), .A2(new_n238), .A3(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G211gat), .B(G218gat), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT74), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n242), .B(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n228), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(G228gat), .A2(G233gat), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n242), .A2(new_n245), .A3(new_n244), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n246), .A2(new_n238), .A3(new_n241), .A4(new_n234), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT3), .B1(new_n253), .B2(new_n227), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n248), .B(new_n250), .C1(new_n254), .C2(new_n224), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n249), .B(KEYINPUT86), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n242), .A2(new_n243), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n234), .A2(new_n244), .A3(new_n238), .A4(new_n241), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(new_n227), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n224), .B1(new_n259), .B2(new_n225), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT29), .B1(new_n224), .B2(new_n225), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n261), .A2(new_n253), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n256), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n255), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(G22gat), .ZN(new_n265));
  INV_X1    g064(.A(G22gat), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n255), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT88), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n265), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n264), .A2(KEYINPUT88), .A3(G22gat), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n205), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n205), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT87), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n255), .A2(new_n263), .A3(new_n266), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n265), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n255), .A2(new_n263), .A3(KEYINPUT87), .A4(new_n266), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n272), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(KEYINPUT89), .B1(new_n271), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n266), .B1(new_n255), .B2(new_n263), .ZN(new_n279));
  NOR3_X1   g078(.A1(new_n267), .A2(new_n279), .A3(KEYINPUT87), .ZN(new_n280));
  INV_X1    g079(.A(new_n276), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n205), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT89), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n279), .B1(KEYINPUT88), .B2(new_n274), .ZN(new_n284));
  INV_X1    g083(.A(new_n270), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n272), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n282), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n278), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT68), .ZN(new_n289));
  NOR2_X1   g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT26), .ZN(new_n292));
  NAND2_X1  g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G183gat), .A2(G190gat), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(new_n291), .B2(new_n292), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT67), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT27), .ZN(new_n299));
  INV_X1    g098(.A(G183gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n302));
  AOI21_X1  g101(.A(G190gat), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT66), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n298), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n294), .B(new_n297), .C1(new_n305), .C2(KEYINPUT28), .ZN(new_n306));
  INV_X1    g105(.A(G190gat), .ZN(new_n307));
  AND2_X1   g106(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT67), .B1(new_n310), .B2(KEYINPUT66), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n301), .A2(new_n302), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n298), .B1(new_n312), .B2(new_n307), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT28), .ZN(new_n314));
  NOR3_X1   g113(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n289), .B1(new_n306), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n296), .B1(new_n311), .B2(new_n314), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n310), .A2(KEYINPUT67), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n305), .A2(KEYINPUT28), .A3(new_n318), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n317), .A2(new_n319), .A3(KEYINPUT68), .A4(new_n294), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(KEYINPUT64), .B(G176gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT23), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n323), .A2(G169gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT65), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT65), .ZN(new_n327));
  INV_X1    g126(.A(G176gat), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n328), .A2(KEYINPUT64), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(KEYINPUT64), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n327), .B(new_n324), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n323), .B1(G169gat), .B2(G176gat), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT24), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n333), .A2(G183gat), .A3(G190gat), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n332), .A2(new_n334), .A3(new_n293), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n300), .A2(new_n307), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n336), .A2(KEYINPUT24), .A3(new_n295), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n326), .A2(new_n331), .A3(new_n335), .A4(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT25), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n335), .A2(new_n337), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n339), .B1(new_n290), .B2(KEYINPUT23), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n321), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(G134gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(G127gat), .ZN(new_n347));
  INV_X1    g146(.A(G127gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G134gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G113gat), .B(G120gat), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n350), .B1(new_n351), .B2(KEYINPUT1), .ZN(new_n352));
  INV_X1    g151(.A(G120gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(G113gat), .ZN(new_n354));
  INV_X1    g153(.A(G113gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G120gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G127gat), .B(G134gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT1), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n352), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G227gat), .ZN(new_n363));
  INV_X1    g162(.A(G233gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n338), .A2(new_n339), .B1(new_n341), .B2(new_n342), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n367), .B1(new_n316), .B2(new_n320), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n352), .A2(new_n360), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n362), .A2(new_n366), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT71), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT72), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT34), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT34), .B1(new_n371), .B2(KEYINPUT72), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n375), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n369), .B1(new_n321), .B2(new_n344), .ZN(new_n378));
  AOI211_X1 g177(.A(new_n361), .B(new_n367), .C1(new_n316), .C2(new_n320), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n365), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT33), .ZN(new_n381));
  XNOR2_X1  g180(.A(G15gat), .B(G43gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(G71gat), .ZN(new_n383));
  INV_X1    g182(.A(G99gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT69), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n381), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(new_n386), .B2(new_n385), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n380), .A2(KEYINPUT32), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT70), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n380), .A2(KEYINPUT70), .A3(KEYINPUT32), .A4(new_n388), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n380), .B1(KEYINPUT32), .B2(new_n381), .ZN(new_n393));
  AOI22_X1  g192(.A1(new_n391), .A2(new_n392), .B1(new_n385), .B2(new_n393), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n377), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n377), .A2(new_n394), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n288), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G226gat), .A2(G233gat), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n345), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n317), .A2(new_n319), .A3(new_n294), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT29), .B1(new_n344), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT75), .B1(new_n402), .B2(new_n399), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n306), .A2(new_n315), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n227), .B1(new_n404), .B2(new_n367), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT75), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(new_n406), .A3(new_n398), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n400), .A2(new_n403), .A3(new_n407), .A4(new_n253), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n344), .A2(new_n399), .A3(new_n401), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n398), .A2(new_n227), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n247), .B(new_n409), .C1(new_n368), .C2(new_n410), .ZN(new_n411));
  XOR2_X1   g210(.A(G8gat), .B(G36gat), .Z(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(G64gat), .ZN(new_n413));
  INV_X1    g212(.A(G92gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n408), .A2(new_n411), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT30), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT77), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n408), .A2(new_n411), .A3(KEYINPUT76), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT76), .B1(new_n408), .B2(new_n411), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n421), .B1(new_n424), .B2(new_n415), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n411), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT76), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n408), .A2(new_n411), .A3(KEYINPUT76), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n428), .A2(new_n421), .A3(new_n429), .A4(new_n415), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n420), .B1(new_n425), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT90), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n428), .A2(new_n429), .A3(new_n415), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT77), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n419), .B1(new_n436), .B2(new_n430), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT90), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n397), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(G141gat), .B(G148gat), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n223), .B1(new_n440), .B2(KEYINPUT2), .ZN(new_n441));
  XNOR2_X1  g240(.A(KEYINPUT78), .B(G141gat), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n210), .B1(new_n442), .B2(G148gat), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n222), .B1(new_n214), .B2(new_n213), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n441), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT3), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n226), .A2(new_n446), .A3(new_n361), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT4), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n369), .A2(new_n224), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT79), .B1(new_n445), .B2(new_n361), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT79), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n369), .A2(new_n224), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(G225gat), .A2(G233gat), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n455), .A2(new_n448), .ZN(new_n456));
  OAI221_X1 g255(.A(new_n447), .B1(new_n448), .B2(new_n449), .C1(new_n453), .C2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT5), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n450), .B(new_n452), .C1(new_n369), .C2(new_n224), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n458), .B1(new_n459), .B2(new_n455), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n445), .A2(new_n361), .A3(KEYINPUT79), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n451), .B1(new_n369), .B2(new_n224), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT4), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT4), .B1(new_n369), .B2(new_n224), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n464), .A2(KEYINPUT81), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT81), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n448), .B1(new_n450), .B2(new_n452), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n468), .B1(new_n469), .B2(new_n465), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n455), .A2(KEYINPUT5), .ZN(new_n472));
  AND4_X1   g271(.A1(KEYINPUT82), .A2(new_n471), .A3(new_n447), .A4(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n447), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n474), .B1(new_n467), .B2(new_n470), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT82), .B1(new_n475), .B2(new_n472), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n461), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  XOR2_X1   g276(.A(G1gat), .B(G29gat), .Z(new_n478));
  XNOR2_X1  g277(.A(G57gat), .B(G85gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n478), .B(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n481));
  XOR2_X1   g280(.A(new_n480), .B(new_n481), .Z(new_n482));
  NAND2_X1  g281(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n461), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT81), .B1(new_n464), .B2(new_n466), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n469), .A2(new_n468), .A3(new_n465), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n447), .B(new_n472), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT82), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n475), .A2(KEYINPUT82), .A3(new_n472), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n484), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n482), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT6), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n483), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT93), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n495), .A2(KEYINPUT93), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT83), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n489), .A2(new_n490), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n492), .B1(new_n499), .B2(new_n461), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n498), .B1(new_n500), .B2(KEYINPUT6), .ZN(new_n501));
  NOR4_X1   g300(.A1(new_n491), .A2(KEYINPUT83), .A3(new_n494), .A4(new_n492), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT94), .ZN(new_n503));
  NOR3_X1   g302(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n477), .A2(KEYINPUT6), .A3(new_n482), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT83), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n500), .A2(new_n498), .A3(KEYINPUT6), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT94), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n496), .B(new_n497), .C1(new_n504), .C2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT35), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n439), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT95), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n506), .A2(new_n495), .A3(new_n507), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n437), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT84), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT84), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n513), .A2(new_n516), .A3(new_n437), .ZN(new_n517));
  INV_X1    g316(.A(new_n397), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n515), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT35), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT95), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n439), .A2(new_n509), .A3(new_n521), .A4(new_n510), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n512), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT39), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n471), .A2(new_n447), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT91), .B1(new_n525), .B2(new_n455), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT91), .ZN(new_n527));
  NOR3_X1   g326(.A1(new_n475), .A2(new_n527), .A3(new_n454), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n524), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT92), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n529), .A2(new_n530), .A3(new_n492), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n525), .A2(KEYINPUT91), .A3(new_n455), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n527), .B1(new_n475), .B2(new_n454), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT39), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT92), .B1(new_n534), .B2(new_n482), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n526), .A2(new_n528), .ZN(new_n536));
  INV_X1    g335(.A(new_n459), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n524), .B1(new_n537), .B2(new_n454), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n531), .A2(new_n535), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n500), .B1(new_n539), .B2(KEYINPUT40), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT40), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n531), .A2(new_n535), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n536), .A2(new_n538), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n540), .A2(new_n544), .A3(new_n434), .A4(new_n438), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n426), .A2(KEYINPUT37), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n546), .A2(new_n415), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT38), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n253), .B(new_n409), .C1(new_n368), .C2(new_n410), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n400), .A2(new_n403), .A3(new_n407), .ZN(new_n550));
  OAI211_X1 g349(.A(KEYINPUT37), .B(new_n549), .C1(new_n550), .C2(new_n253), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n547), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n424), .A2(KEYINPUT37), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n547), .A2(new_n553), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n417), .B(new_n552), .C1(new_n554), .C2(new_n548), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n545), .B(new_n288), .C1(new_n509), .C2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n395), .ZN(new_n557));
  INV_X1    g356(.A(new_n396), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT36), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n515), .A2(new_n517), .ZN(new_n561));
  INV_X1    g360(.A(new_n288), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n556), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n523), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G15gat), .B(G22gat), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT16), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n566), .B1(new_n567), .B2(G1gat), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n568), .B1(G1gat), .B2(new_n566), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n569), .B(G8gat), .Z(new_n570));
  INV_X1    g369(.A(KEYINPUT21), .ZN(new_n571));
  XNOR2_X1  g370(.A(G57gat), .B(G64gat), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n573));
  OR3_X1    g372(.A1(new_n572), .A2(KEYINPUT101), .A3(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(G71gat), .B(G78gat), .Z(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n570), .B1(new_n571), .B2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT102), .ZN(new_n578));
  AND2_X1   g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n571), .ZN(new_n581));
  XOR2_X1   g380(.A(G127gat), .B(G155gat), .Z(new_n582));
  XOR2_X1   g381(.A(new_n581), .B(new_n582), .Z(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n586));
  XNOR2_X1  g385(.A(G183gat), .B(G211gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n580), .A2(new_n584), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n585), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n588), .B1(new_n585), .B2(new_n589), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G43gat), .B(G50gat), .Z(new_n593));
  INV_X1    g392(.A(KEYINPUT96), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G43gat), .B(G50gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT96), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n595), .A2(KEYINPUT15), .A3(new_n597), .ZN(new_n598));
  NOR3_X1   g397(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n599), .A2(KEYINPUT97), .B1(G29gat), .B2(G36gat), .ZN(new_n600));
  INV_X1    g399(.A(G29gat), .ZN(new_n601));
  INV_X1    g400(.A(G36gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT14), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n600), .B1(new_n604), .B2(KEYINPUT97), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n598), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n595), .A2(KEYINPUT15), .A3(new_n597), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT15), .ZN(new_n608));
  INV_X1    g407(.A(G43gat), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n609), .A2(KEYINPUT98), .A3(G50gat), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n608), .B(new_n610), .C1(new_n593), .C2(KEYINPUT98), .ZN(new_n611));
  NAND2_X1  g410(.A1(G29gat), .A2(G36gat), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n612), .B(KEYINPUT99), .Z(new_n613));
  NAND4_X1  g412(.A1(new_n607), .A2(new_n604), .A3(new_n611), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n606), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT17), .ZN(new_n616));
  NAND2_X1  g415(.A1(G85gat), .A2(G92gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT7), .ZN(new_n618));
  NAND2_X1  g417(.A1(G99gat), .A2(G106gat), .ZN(new_n619));
  INV_X1    g418(.A(G85gat), .ZN(new_n620));
  AOI22_X1  g419(.A1(KEYINPUT8), .A2(new_n619), .B1(new_n620), .B2(new_n414), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G99gat), .B(G106gat), .Z(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT103), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n622), .A2(new_n623), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n625), .B(new_n626), .Z(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n616), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT104), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(G232gat), .A2(G233gat), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n627), .A2(new_n615), .B1(KEYINPUT41), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G134gat), .B(G162gat), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n632), .A2(KEYINPUT41), .ZN(new_n637));
  XNOR2_X1  g436(.A(G190gat), .B(G218gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n635), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n631), .A2(new_n640), .A3(new_n633), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n636), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n639), .B1(new_n636), .B2(new_n641), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n592), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n615), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n646), .A2(new_n570), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n616), .B2(new_n570), .ZN(new_n648));
  NAND2_X1  g447(.A1(G229gat), .A2(G233gat), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT100), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n651), .A2(KEYINPUT18), .ZN(new_n652));
  OR2_X1    g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n646), .B(new_n570), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n649), .B(KEYINPUT13), .Z(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n650), .A2(new_n652), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n653), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT11), .B(G169gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G197gat), .ZN(new_n660));
  XOR2_X1   g459(.A(G113gat), .B(G141gat), .Z(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT12), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n653), .A2(new_n663), .A3(new_n656), .A4(new_n657), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n626), .A2(KEYINPUT105), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(new_n624), .ZN(new_n670));
  INV_X1    g469(.A(new_n576), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n627), .A2(new_n576), .ZN(new_n673));
  AOI21_X1  g472(.A(KEYINPUT10), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n627), .A2(KEYINPUT10), .A3(new_n671), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(G230gat), .ZN(new_n677));
  OAI22_X1  g476(.A1(new_n674), .A2(new_n676), .B1(new_n677), .B2(new_n364), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n364), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n672), .A2(new_n673), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(KEYINPUT106), .ZN(new_n682));
  XNOR2_X1  g481(.A(G120gat), .B(G148gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(new_n328), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(new_n232), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n682), .B(new_n686), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n645), .A2(new_n668), .A3(new_n687), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n565), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n513), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g491(.A1(new_n434), .A2(new_n438), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT16), .B(G8gat), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n695), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n697), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n699), .B1(KEYINPUT107), .B2(KEYINPUT42), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT42), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n701), .B1(new_n695), .B2(G8gat), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n689), .A2(new_n694), .A3(new_n699), .ZN(new_n703));
  AOI22_X1  g502(.A1(new_n698), .A2(new_n700), .B1(new_n702), .B2(new_n703), .ZN(G1325gat));
  AOI21_X1  g503(.A(G15gat), .B1(new_n689), .B2(new_n559), .ZN(new_n705));
  INV_X1    g504(.A(new_n560), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n689), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n705), .B1(G15gat), .B2(new_n707), .ZN(G1326gat));
  NAND2_X1  g507(.A1(new_n689), .A2(new_n562), .ZN(new_n709));
  XNOR2_X1  g508(.A(KEYINPUT43), .B(G22gat), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1327gat));
  AOI21_X1  g510(.A(new_n644), .B1(new_n523), .B2(new_n564), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n592), .A2(new_n668), .A3(new_n687), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n716), .A2(new_n601), .A3(new_n690), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT45), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n642), .B2(new_n643), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n636), .A2(new_n641), .ZN(new_n721));
  INV_X1    g520(.A(new_n639), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n636), .A2(new_n639), .A3(new_n641), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n723), .A2(KEYINPUT108), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n720), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n565), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n727), .B2(new_n712), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n731), .A2(new_n714), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n690), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n718), .B1(new_n734), .B2(new_n601), .ZN(G1328gat));
  NAND3_X1  g534(.A1(new_n716), .A2(new_n602), .A3(new_n694), .ZN(new_n736));
  XOR2_X1   g535(.A(KEYINPUT109), .B(KEYINPUT46), .Z(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n732), .A2(new_n694), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n740), .B2(new_n602), .ZN(G1329gat));
  AND4_X1   g540(.A1(new_n609), .A2(new_n712), .A3(new_n559), .A4(new_n714), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n731), .A2(new_n706), .A3(new_n714), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n742), .B1(new_n743), .B2(G43gat), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g544(.A1(new_n731), .A2(G50gat), .A3(new_n562), .A4(new_n714), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n712), .A2(KEYINPUT110), .A3(new_n714), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT110), .B1(new_n712), .B2(new_n714), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n747), .A2(new_n748), .A3(new_n288), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n746), .B1(new_n749), .B2(G50gat), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT48), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT48), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n746), .B(new_n752), .C1(new_n749), .C2(G50gat), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(G1331gat));
  NOR2_X1   g553(.A1(new_n645), .A2(new_n667), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n565), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n687), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n690), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g559(.A(KEYINPUT49), .B(G64gat), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n758), .A2(new_n694), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n763));
  OAI22_X1  g562(.A1(new_n757), .A2(new_n693), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n763), .B1(new_n762), .B2(new_n764), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(G1333gat));
  INV_X1    g566(.A(G71gat), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n758), .A2(new_n768), .A3(new_n559), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT50), .ZN(new_n770));
  OAI21_X1  g569(.A(G71gat), .B1(new_n757), .B2(new_n560), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n770), .B1(new_n769), .B2(new_n771), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(G1334gat));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n562), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G78gat), .ZN(G1335gat));
  INV_X1    g575(.A(new_n687), .ZN(new_n777));
  INV_X1    g576(.A(new_n644), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n592), .A2(new_n667), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n565), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT51), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g582(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n712), .A2(new_n779), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n777), .B1(new_n783), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(G85gat), .B1(new_n787), .B2(new_n690), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n779), .A2(new_n687), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(KEYINPUT112), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n731), .A2(G85gat), .A3(new_n690), .A4(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(KEYINPUT114), .B1(new_n788), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n786), .ZN(new_n794));
  AOI22_X1  g593(.A1(new_n712), .A2(new_n779), .B1(new_n781), .B2(KEYINPUT51), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n690), .B(new_n687), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n620), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n797), .A2(new_n798), .A3(new_n791), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n793), .A2(new_n799), .ZN(G1336gat));
  XNOR2_X1  g599(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(G92gat), .B1(new_n787), .B2(new_n694), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n731), .A2(G92gat), .A3(new_n694), .A4(new_n790), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n802), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n694), .B(new_n687), .C1(new_n794), .C2(new_n795), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n414), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n808), .A2(new_n801), .A3(new_n804), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n806), .A2(new_n809), .ZN(G1337gat));
  NAND3_X1  g609(.A1(new_n787), .A2(new_n384), .A3(new_n559), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n731), .A2(new_n706), .A3(new_n790), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n811), .B1(new_n813), .B2(new_n384), .ZN(G1338gat));
  AOI21_X1  g613(.A(new_n727), .B1(new_n565), .B2(new_n778), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n728), .B1(new_n523), .B2(new_n564), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n562), .B(new_n790), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n731), .A2(KEYINPUT117), .A3(new_n562), .A4(new_n790), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n819), .A2(G106gat), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n783), .A2(new_n786), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n777), .A2(G106gat), .A3(new_n288), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(KEYINPUT116), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI22_X1  g626(.A1(new_n822), .A2(new_n824), .B1(new_n817), .B2(G106gat), .ZN(new_n828));
  OAI22_X1  g627(.A1(new_n821), .A2(new_n827), .B1(new_n826), .B2(new_n828), .ZN(G1339gat));
  NOR2_X1   g628(.A1(new_n681), .A2(new_n685), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n672), .A2(new_n673), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT10), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n833), .A2(new_n679), .A3(new_n675), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n834), .A2(new_n678), .A3(KEYINPUT54), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n685), .B1(new_n678), .B2(KEYINPUT54), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n830), .B1(new_n837), .B2(KEYINPUT55), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n839), .B1(new_n835), .B2(new_n836), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n834), .A2(new_n678), .A3(KEYINPUT54), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n843), .B(new_n685), .C1(KEYINPUT54), .C2(new_n678), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n844), .A2(KEYINPUT118), .A3(new_n839), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n838), .A2(new_n842), .A3(new_n845), .A4(new_n667), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n648), .A2(new_n649), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n654), .A2(new_n655), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n662), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n666), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n687), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n846), .A2(new_n851), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n720), .A2(new_n725), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n838), .A2(new_n842), .A3(new_n845), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n726), .A2(new_n855), .A3(new_n850), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n592), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n645), .A2(new_n667), .A3(new_n687), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n859), .A2(new_n513), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n439), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(new_n668), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(new_n355), .ZN(G1340gat));
  OAI21_X1  g662(.A(G120gat), .B1(new_n861), .B2(new_n777), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n687), .A2(new_n353), .ZN(new_n865));
  XOR2_X1   g664(.A(new_n865), .B(KEYINPUT119), .Z(new_n866));
  OAI21_X1  g665(.A(new_n864), .B1(new_n861), .B2(new_n866), .ZN(G1341gat));
  INV_X1    g666(.A(new_n592), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n861), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(new_n348), .ZN(G1342gat));
  NAND3_X1  g669(.A1(new_n860), .A2(new_n439), .A3(new_n778), .ZN(new_n871));
  OR3_X1    g670(.A1(new_n871), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(G134gat), .ZN(new_n873));
  OAI21_X1  g672(.A(KEYINPUT56), .B1(new_n871), .B2(G134gat), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(G1343gat));
  INV_X1    g674(.A(KEYINPUT120), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n876), .B(new_n690), .C1(new_n857), .C2(new_n858), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n560), .A2(new_n562), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT120), .B1(new_n859), .B2(new_n513), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n667), .A2(new_n209), .ZN(new_n882));
  XOR2_X1   g681(.A(new_n882), .B(KEYINPUT121), .Z(new_n883));
  NAND4_X1  g682(.A1(new_n880), .A2(new_n693), .A3(new_n881), .A4(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n838), .A2(new_n842), .A3(new_n845), .A4(new_n850), .ZN(new_n886));
  AOI22_X1  g685(.A1(new_n665), .A2(new_n666), .B1(new_n844), .B2(new_n839), .ZN(new_n887));
  AOI22_X1  g686(.A1(new_n887), .A2(new_n838), .B1(new_n687), .B2(new_n850), .ZN(new_n888));
  OAI22_X1  g687(.A1(new_n853), .A2(new_n886), .B1(new_n888), .B2(new_n778), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n858), .B1(new_n889), .B2(new_n868), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT57), .B1(new_n890), .B2(new_n288), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n892), .B(new_n562), .C1(new_n857), .C2(new_n858), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n706), .A2(new_n513), .A3(new_n694), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n891), .A2(new_n893), .A3(new_n667), .A4(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n442), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n884), .A2(new_n885), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n885), .B1(new_n884), .B2(new_n897), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT58), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n895), .A2(new_n896), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n877), .A2(new_n693), .A3(new_n879), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n726), .B1(new_n846), .B2(new_n851), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n853), .A2(new_n886), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n868), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n858), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n876), .B1(new_n908), .B2(new_n690), .ZN(new_n909));
  INV_X1    g708(.A(new_n883), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n903), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT122), .B1(new_n902), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n884), .A2(new_n885), .A3(new_n897), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT58), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n901), .A2(new_n914), .ZN(G1344gat));
  INV_X1    g714(.A(KEYINPUT59), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT57), .B1(new_n859), .B2(new_n288), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n888), .A2(new_n778), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n855), .A2(new_n778), .A3(new_n850), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n592), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n892), .B(new_n562), .C1(new_n920), .C2(new_n858), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n687), .A3(new_n894), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n916), .B1(new_n923), .B2(G148gat), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n916), .B1(new_n925), .B2(new_n777), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n926), .A2(new_n219), .ZN(new_n927));
  INV_X1    g726(.A(new_n903), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n881), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n687), .A2(new_n219), .ZN(new_n930));
  OAI22_X1  g729(.A1(new_n924), .A2(new_n927), .B1(new_n929), .B2(new_n930), .ZN(G1345gat));
  NOR3_X1   g730(.A1(new_n925), .A2(new_n216), .A3(new_n868), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n928), .A2(new_n592), .A3(new_n881), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(new_n933), .B2(new_n216), .ZN(G1346gat));
  NAND4_X1  g733(.A1(new_n928), .A2(new_n217), .A3(new_n778), .A4(new_n881), .ZN(new_n935));
  OAI21_X1  g734(.A(G162gat), .B1(new_n925), .B2(new_n853), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT123), .ZN(G1347gat));
  NOR4_X1   g737(.A1(new_n859), .A2(new_n690), .A3(new_n693), .A4(new_n397), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(G169gat), .B1(new_n940), .B2(new_n668), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n859), .A2(new_n690), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(KEYINPUT124), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n944), .B1(new_n859), .B2(new_n690), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n943), .A2(new_n945), .A3(new_n694), .A4(new_n518), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n946), .A2(G169gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n941), .B1(new_n947), .B2(new_n668), .ZN(G1348gat));
  AND3_X1   g747(.A1(new_n939), .A2(new_n322), .A3(new_n687), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n946), .A2(new_n777), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n949), .B1(new_n950), .B2(new_n328), .ZN(G1349gat));
  NAND4_X1  g750(.A1(new_n942), .A2(new_n694), .A3(new_n518), .A4(new_n592), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(KEYINPUT125), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT125), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n939), .A2(new_n954), .A3(new_n592), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n953), .A2(G183gat), .A3(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n592), .A2(new_n312), .ZN(new_n958));
  OAI21_X1  g757(.A(KEYINPUT126), .B1(new_n946), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(KEYINPUT60), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n946), .A2(new_n958), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT60), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n961), .A2(KEYINPUT126), .A3(new_n956), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n960), .A2(new_n963), .ZN(G1350gat));
  OAI21_X1  g763(.A(G190gat), .B1(new_n940), .B2(new_n644), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n965), .A2(KEYINPUT61), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n965), .A2(KEYINPUT61), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n726), .A2(new_n307), .ZN(new_n968));
  OAI22_X1  g767(.A1(new_n966), .A2(new_n967), .B1(new_n946), .B2(new_n968), .ZN(G1351gat));
  NOR3_X1   g768(.A1(new_n706), .A2(new_n690), .A3(new_n693), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n922), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g770(.A(G197gat), .B1(new_n971), .B2(new_n668), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n943), .A2(new_n945), .A3(new_n694), .A4(new_n879), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n973), .A2(G197gat), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n972), .B1(new_n974), .B2(new_n668), .ZN(G1352gat));
  NAND2_X1  g774(.A1(new_n687), .A2(new_n232), .ZN(new_n976));
  OR3_X1    g775(.A1(new_n973), .A2(KEYINPUT62), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g776(.A(KEYINPUT62), .B1(new_n973), .B2(new_n976), .ZN(new_n978));
  AND3_X1   g777(.A1(new_n922), .A2(new_n687), .A3(new_n970), .ZN(new_n979));
  OAI211_X1 g778(.A(new_n977), .B(new_n978), .C1(new_n232), .C2(new_n979), .ZN(G1353gat));
  NAND4_X1  g779(.A1(new_n917), .A2(new_n592), .A3(new_n921), .A4(new_n970), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(G211gat), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT63), .ZN(new_n983));
  XNOR2_X1  g782(.A(new_n982), .B(new_n983), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n973), .A2(new_n868), .ZN(new_n985));
  AOI21_X1  g784(.A(KEYINPUT127), .B1(new_n985), .B2(new_n236), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT127), .ZN(new_n987));
  NOR4_X1   g786(.A1(new_n973), .A2(new_n987), .A3(G211gat), .A4(new_n868), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n984), .B1(new_n986), .B2(new_n988), .ZN(G1354gat));
  NOR3_X1   g788(.A1(new_n971), .A2(new_n237), .A3(new_n644), .ZN(new_n990));
  OR2_X1    g789(.A1(new_n973), .A2(new_n853), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n990), .B1(new_n237), .B2(new_n991), .ZN(G1355gat));
endmodule


