//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 0 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1279,
    new_n1280, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1346, new_n1347,
    new_n1348;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G58), .ZN(new_n206));
  INV_X1    g0006(.A(G68), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G50), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  OR3_X1    g0011(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G1), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n210), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT0), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT65), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n220), .A2(KEYINPUT66), .A3(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT64), .B(G68), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n226), .B1(G238), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n222), .A2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(KEYINPUT66), .B1(new_n220), .B2(new_n221), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n215), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n212), .B(new_n218), .C1(new_n231), .C2(KEYINPUT1), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT67), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT68), .B(KEYINPUT69), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT70), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n247), .B(new_n251), .ZN(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n211), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G33), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n256), .A2(new_n258), .A3(new_n210), .A4(G87), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT22), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT3), .B(G33), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT22), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n261), .A2(new_n262), .A3(new_n210), .A4(G87), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT23), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(new_n203), .A3(G20), .ZN(new_n266));
  INV_X1    g0066(.A(G116), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n210), .A2(G33), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n203), .A2(KEYINPUT73), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT73), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G107), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n270), .A2(new_n272), .A3(G20), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n269), .B1(KEYINPUT23), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT24), .ZN(new_n275));
  AND3_X1   g0075(.A1(new_n264), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n275), .B1(new_n264), .B2(new_n274), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n254), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G13), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(G1), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(G20), .A3(new_n203), .ZN(new_n281));
  XNOR2_X1  g0081(.A(new_n281), .B(KEYINPUT25), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n213), .A2(G13), .A3(G20), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n213), .A2(G33), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n283), .A2(new_n284), .A3(new_n211), .A4(new_n253), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(new_n203), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n278), .A2(new_n287), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n256), .A2(new_n258), .A3(G257), .A4(G1698), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n256), .A2(new_n258), .A3(G250), .A4(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G294), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n289), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G45), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(G1), .ZN(new_n297));
  NAND2_X1  g0097(.A1(KEYINPUT5), .A2(G41), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(KEYINPUT5), .A2(G41), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n297), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G41), .ZN(new_n302));
  OAI211_X1 g0102(.A(G1), .B(G13), .C1(new_n255), .C2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n301), .A2(G264), .A3(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n297), .B(G274), .C1(new_n300), .C2(new_n299), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n295), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT85), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n295), .A2(new_n304), .A3(KEYINPUT85), .A4(new_n305), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G190), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AND3_X1   g0112(.A1(new_n295), .A2(new_n304), .A3(new_n305), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n313), .A2(G200), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n288), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n287), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n264), .A2(new_n274), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT24), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n264), .A2(new_n274), .A3(new_n275), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n317), .B1(new_n321), .B2(new_n254), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n308), .A2(G169), .A3(new_n309), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n313), .A2(G179), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n322), .B1(new_n325), .B2(KEYINPUT86), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT86), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n323), .A2(new_n327), .A3(new_n324), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n316), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n283), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(new_n254), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n213), .A2(G20), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G50), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G50), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n331), .A2(new_n334), .B1(new_n335), .B2(new_n330), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT8), .B(G58), .ZN(new_n337));
  INV_X1    g0137(.A(G150), .ZN(new_n338));
  NOR2_X1   g0138(.A1(G20), .A2(G33), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  OAI22_X1  g0140(.A1(new_n337), .A2(new_n268), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(G50), .A2(G58), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n210), .B1(new_n342), .B2(new_n207), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g0144(.A1(new_n253), .A2(new_n211), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n336), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n346), .A2(KEYINPUT9), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(KEYINPUT9), .ZN(new_n348));
  AOI21_X1  g0148(.A(G1), .B1(new_n302), .B2(new_n296), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n294), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G226), .ZN(new_n351));
  OR2_X1    g0151(.A1(KEYINPUT71), .A2(G45), .ZN(new_n352));
  NAND2_X1  g0152(.A1(KEYINPUT71), .A2(G45), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(new_n302), .A3(new_n353), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n213), .A2(G274), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n261), .A2(G222), .A3(new_n290), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n261), .A2(G1698), .ZN(new_n359));
  INV_X1    g0159(.A(G223), .ZN(new_n360));
  OAI221_X1 g0160(.A(new_n358), .B1(new_n224), .B2(new_n261), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n357), .B1(new_n361), .B2(new_n294), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n347), .A2(new_n348), .B1(G190), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT75), .ZN(new_n364));
  INV_X1    g0164(.A(G200), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n364), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n361), .A2(new_n294), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n367), .A2(new_n356), .A3(new_n351), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n368), .A2(KEYINPUT75), .A3(G200), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n363), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT10), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT10), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n363), .A2(new_n366), .A3(new_n372), .A4(new_n369), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n368), .A2(G179), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n346), .B1(new_n362), .B2(G169), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g0177(.A(new_n377), .B(KEYINPUT72), .ZN(new_n378));
  OAI22_X1  g0178(.A1(new_n337), .A2(new_n340), .B1(new_n210), .B2(new_n224), .ZN(new_n379));
  XNOR2_X1  g0179(.A(KEYINPUT15), .B(G87), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n380), .A2(new_n268), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n254), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT74), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n382), .B(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n332), .A2(G77), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n331), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n330), .A2(new_n224), .ZN(new_n388));
  AND2_X1   g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n261), .A2(G232), .A3(new_n290), .ZN(new_n391));
  XNOR2_X1  g0191(.A(KEYINPUT73), .B(G107), .ZN(new_n392));
  INV_X1    g0192(.A(G238), .ZN(new_n393));
  OAI221_X1 g0193(.A(new_n391), .B1(new_n261), .B2(new_n392), .C1(new_n359), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n294), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n350), .A2(G244), .B1(new_n355), .B2(new_n354), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G169), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n390), .B(new_n399), .C1(G179), .C2(new_n397), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n397), .A2(G200), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n395), .A2(G190), .A3(new_n396), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n401), .A2(new_n384), .A3(new_n389), .A4(new_n402), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n374), .A2(new_n378), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT16), .ZN(new_n406));
  AND2_X1   g0206(.A1(KEYINPUT64), .A2(G68), .ZN(new_n407));
  NOR2_X1   g0207(.A1(KEYINPUT64), .A2(G68), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n208), .B1(new_n409), .B2(new_n206), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G20), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n339), .A2(G159), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT7), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(new_n261), .B2(G20), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n256), .A2(new_n258), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n416), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n409), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n406), .B1(new_n413), .B2(new_n418), .ZN(new_n419));
  NOR3_X1   g0219(.A1(new_n261), .A2(new_n414), .A3(G20), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT7), .B1(new_n416), .B2(new_n210), .ZN(new_n421));
  OAI21_X1  g0221(.A(G68), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n422), .A2(KEYINPUT16), .A3(new_n411), .A4(new_n412), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n419), .A2(new_n423), .A3(new_n254), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n337), .B1(new_n213), .B2(G20), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n425), .A2(new_n331), .B1(new_n330), .B2(new_n337), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n256), .A2(new_n258), .A3(G226), .A4(G1698), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n256), .A2(new_n258), .A3(G223), .A4(new_n290), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G33), .A2(G87), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n294), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n350), .A2(G232), .B1(new_n355), .B2(new_n354), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(G169), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n432), .A2(new_n433), .A3(G179), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n427), .A2(KEYINPUT18), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT79), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n427), .A2(KEYINPUT79), .A3(KEYINPUT18), .A4(new_n437), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n427), .A2(new_n437), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT18), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n440), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT80), .B1(new_n434), .B2(G190), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n434), .A2(new_n365), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT80), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n432), .A2(new_n433), .A3(new_n448), .A4(new_n311), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n446), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(new_n424), .A3(new_n426), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT17), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n450), .A2(KEYINPUT17), .A3(new_n424), .A4(new_n426), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n445), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g0256(.A(KEYINPUT78), .B(KEYINPUT14), .Z(new_n457));
  NAND4_X1  g0257(.A1(new_n256), .A2(new_n258), .A3(G232), .A4(G1698), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n256), .A2(new_n258), .A3(G226), .A4(new_n290), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n458), .B(new_n459), .C1(new_n255), .C2(new_n202), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n294), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n350), .A2(G238), .B1(new_n355), .B2(new_n354), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT13), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n463), .B1(new_n461), .B2(new_n462), .ZN(new_n465));
  OAI211_X1 g0265(.A(G169), .B(new_n457), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n461), .A2(new_n462), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT13), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n468), .A2(G179), .A3(new_n469), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n398), .B1(new_n468), .B2(new_n469), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT14), .B1(new_n472), .B2(KEYINPUT77), .ZN(new_n473));
  OAI211_X1 g0273(.A(KEYINPUT77), .B(G169), .C1(new_n464), .C2(new_n465), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n471), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n227), .A2(new_n210), .ZN(new_n477));
  OAI22_X1  g0277(.A1(new_n340), .A2(new_n335), .B1(new_n268), .B2(new_n224), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n254), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT11), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(KEYINPUT11), .B(new_n254), .C1(new_n477), .C2(new_n478), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT76), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT76), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n481), .A2(new_n485), .A3(new_n482), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n477), .A2(KEYINPUT12), .A3(new_n280), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n331), .A2(G68), .A3(new_n332), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT12), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n489), .B1(new_n283), .B2(G68), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n487), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n484), .A2(new_n486), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n476), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n492), .ZN(new_n494));
  OAI21_X1  g0294(.A(G200), .B1(new_n464), .B2(new_n465), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n468), .A2(G190), .A3(new_n469), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n405), .A2(new_n456), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n301), .A2(G270), .A3(new_n303), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n500), .A2(new_n305), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n256), .A2(new_n258), .A3(G264), .A4(G1698), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n256), .A2(new_n258), .A3(G257), .A4(new_n290), .ZN(new_n503));
  INV_X1    g0303(.A(G303), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n502), .B(new_n503), .C1(new_n504), .C2(new_n261), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n294), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT84), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n501), .A2(new_n506), .A3(KEYINPUT84), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G283), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n511), .B(new_n210), .C1(G33), .C2(new_n202), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n267), .A2(G20), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n512), .A2(new_n254), .A3(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT20), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n512), .A2(KEYINPUT20), .A3(new_n254), .A4(new_n513), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n283), .A2(G116), .ZN(new_n519));
  INV_X1    g0319(.A(new_n285), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n519), .B1(new_n520), .B2(G116), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n398), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n509), .A2(new_n510), .A3(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT21), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n501), .A2(new_n506), .A3(G179), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n518), .A2(new_n521), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n509), .A2(KEYINPUT21), .A3(new_n510), .A4(new_n522), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n525), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n501), .A2(new_n506), .A3(KEYINPUT84), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT84), .B1(new_n501), .B2(new_n506), .ZN(new_n532));
  OAI21_X1  g0332(.A(G190), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n509), .A2(G200), .A3(new_n510), .ZN(new_n534));
  INV_X1    g0334(.A(new_n527), .ZN(new_n535));
  AND3_X1   g0335(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n530), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n301), .A2(G257), .A3(new_n303), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT82), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n538), .A2(new_n539), .A3(new_n305), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n539), .B1(new_n538), .B2(new_n305), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n256), .A2(new_n258), .A3(G244), .A4(new_n290), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT4), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n261), .A2(KEYINPUT4), .A3(G244), .A4(new_n290), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n261), .A2(G250), .A3(G1698), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n511), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n294), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n542), .A2(G190), .A3(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n283), .A2(G97), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(new_n520), .B2(G97), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n392), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n420), .B2(new_n421), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n339), .A2(G77), .ZN(new_n556));
  XNOR2_X1  g0356(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G97), .A2(G107), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n204), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT6), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n560), .A2(KEYINPUT81), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n560), .A2(KEYINPUT81), .ZN(new_n562));
  OAI22_X1  g0362(.A1(new_n561), .A2(new_n562), .B1(new_n202), .B2(G107), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n559), .A2(new_n563), .A3(G20), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n555), .A2(new_n556), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n553), .B1(new_n565), .B2(new_n254), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n538), .A2(new_n305), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT82), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n538), .A2(new_n539), .A3(new_n305), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n549), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n550), .B(new_n566), .C1(new_n570), .C2(new_n365), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n549), .A2(new_n568), .A3(new_n569), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n398), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n564), .A2(new_n556), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n392), .B1(new_n415), .B2(new_n417), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n254), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n552), .ZN(new_n577));
  INV_X1    g0377(.A(G179), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n542), .A2(new_n578), .A3(new_n549), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n573), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n256), .A2(new_n258), .A3(new_n210), .A4(G68), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT19), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n268), .B2(new_n202), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(G87), .A2(G97), .ZN(new_n585));
  NAND3_X1  g0385(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n392), .A2(new_n585), .B1(new_n210), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n254), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n380), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n589), .A2(new_n283), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n285), .A2(new_n380), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n588), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n393), .A2(new_n290), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n225), .A2(G1698), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n256), .A2(new_n595), .A3(new_n258), .A4(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n255), .A2(new_n267), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n303), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(G250), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n601), .B1(new_n213), .B2(G45), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n303), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n355), .A2(G45), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n398), .B1(new_n600), .B2(new_n605), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n303), .A2(new_n602), .B1(new_n355), .B2(G45), .ZN(new_n607));
  NOR2_X1   g0407(.A1(G238), .A2(G1698), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(new_n225), .B2(G1698), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n598), .B1(new_n609), .B2(new_n261), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n578), .B(new_n607), .C1(new_n610), .C2(new_n303), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n594), .A2(new_n606), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n270), .A2(new_n272), .A3(new_n585), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n586), .A2(new_n210), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n615), .A2(new_n581), .A3(new_n583), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n590), .B1(new_n616), .B2(new_n254), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n520), .A2(G87), .ZN(new_n618));
  OAI21_X1  g0418(.A(G200), .B1(new_n600), .B2(new_n605), .ZN(new_n619));
  OAI211_X1 g0419(.A(G190), .B(new_n607), .C1(new_n610), .C2(new_n303), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n617), .A2(new_n618), .A3(new_n619), .A4(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT83), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n612), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n622), .B1(new_n612), .B2(new_n621), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n571), .B(new_n580), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  AND4_X1   g0426(.A1(new_n329), .A2(new_n499), .A3(new_n537), .A4(new_n626), .ZN(G372));
  INV_X1    g0427(.A(new_n378), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n493), .B1(new_n629), .B2(new_n400), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n455), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n444), .A2(new_n438), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n628), .B1(new_n633), .B2(new_n374), .ZN(new_n634));
  AOI211_X1 g0434(.A(new_n592), .B(new_n590), .C1(new_n616), .C2(new_n254), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n606), .A2(new_n611), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n619), .A2(new_n620), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n588), .A2(new_n591), .A3(new_n618), .ZN(new_n638));
  OAI22_X1  g0438(.A1(new_n635), .A2(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT83), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n612), .A2(new_n621), .A3(new_n622), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n580), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT26), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n643), .B1(new_n580), .B2(new_n639), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT88), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n642), .A2(KEYINPUT26), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n640), .A2(new_n641), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n573), .A2(new_n577), .A3(new_n579), .ZN(new_n648));
  AND4_X1   g0448(.A1(new_n645), .A2(new_n647), .A3(KEYINPUT26), .A4(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n612), .A2(KEYINPUT87), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT87), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n594), .A2(new_n652), .A3(new_n606), .A4(new_n611), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n530), .B1(new_n288), .B2(new_n325), .ZN(new_n656));
  AOI21_X1  g0456(.A(G190), .B1(new_n308), .B2(new_n309), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n322), .B1(new_n657), .B2(new_n314), .ZN(new_n658));
  INV_X1    g0458(.A(new_n639), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n658), .A2(new_n659), .A3(new_n580), .A4(new_n571), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n655), .B1(new_n656), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n499), .B1(new_n650), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n634), .A2(new_n662), .ZN(G369));
  INV_X1    g0463(.A(new_n280), .ZN(new_n664));
  OR3_X1    g0464(.A1(new_n664), .A2(KEYINPUT27), .A3(G20), .ZN(new_n665));
  OAI21_X1  g0465(.A(KEYINPUT27), .B1(new_n664), .B2(G20), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(G213), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G343), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(new_n535), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n530), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n537), .ZN(new_n673));
  OAI211_X1 g0473(.A(KEYINPUT89), .B(new_n672), .C1(new_n673), .C2(new_n671), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n672), .A2(KEYINPUT89), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G330), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n329), .B1(new_n322), .B2(new_n670), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n326), .A2(new_n328), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n678), .B1(new_n679), .B2(new_n670), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n530), .A2(new_n670), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n329), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n325), .A2(new_n288), .A3(new_n670), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n681), .A2(new_n686), .ZN(G399));
  INV_X1    g0487(.A(new_n216), .ZN(new_n688));
  OAI21_X1  g0488(.A(KEYINPUT90), .B1(new_n688), .B2(G41), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n688), .A2(KEYINPUT90), .A3(G41), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n613), .A2(G116), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(G1), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n209), .B2(new_n693), .ZN(new_n696));
  XOR2_X1   g0496(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT92), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n696), .B(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n642), .A2(new_n645), .A3(KEYINPUT26), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n647), .A2(KEYINPUT26), .A3(new_n648), .ZN(new_n701));
  AOI22_X1  g0501(.A1(new_n572), .A2(new_n398), .B1(new_n576), .B2(new_n552), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n659), .A2(new_n702), .A3(new_n579), .ZN(new_n703));
  AOI21_X1  g0503(.A(KEYINPUT88), .B1(new_n703), .B2(new_n643), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n700), .B1(new_n701), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n571), .A2(new_n580), .A3(new_n659), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(new_n316), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n325), .A2(new_n288), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n708), .A2(new_n525), .A3(new_n528), .A4(new_n529), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n654), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n669), .B1(new_n705), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT29), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n329), .A2(new_n537), .A3(new_n626), .A4(new_n670), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n600), .A2(new_n605), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n715), .A2(new_n304), .A3(new_n295), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n716), .A2(new_n526), .A3(new_n549), .A4(new_n542), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT30), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(KEYINPUT93), .B1(new_n600), .B2(new_n605), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT93), .ZN(new_n721));
  OAI211_X1 g0521(.A(new_n721), .B(new_n607), .C1(new_n610), .C2(new_n303), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n720), .A2(new_n722), .A3(new_n578), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(new_n313), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n724), .A2(new_n509), .A3(new_n510), .A4(new_n572), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n570), .A2(KEYINPUT30), .A3(new_n526), .A4(new_n716), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n719), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n669), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT31), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n727), .A2(KEYINPUT31), .A3(new_n669), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n714), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G330), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n654), .A2(KEYINPUT94), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT94), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n651), .A2(new_n735), .A3(new_n653), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n643), .B1(new_n648), .B2(new_n659), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n642), .A2(new_n643), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n530), .B1(new_n326), .B2(new_n328), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n739), .B(new_n740), .C1(new_n660), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n670), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n713), .B(new_n733), .C1(new_n744), .C2(new_n712), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT95), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n745), .B(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n699), .B1(new_n747), .B2(G1), .ZN(G364));
  AND2_X1   g0548(.A1(new_n674), .A2(new_n675), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n749), .A2(G330), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n279), .A2(G20), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n213), .B1(new_n751), .B2(G45), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n692), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT96), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n676), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n674), .A2(KEYINPUT96), .A3(G330), .A4(new_n675), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n750), .A2(new_n755), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G13), .A2(G33), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n211), .B1(G20), .B2(new_n398), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n688), .A2(new_n261), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n352), .A2(new_n353), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n766), .B1(new_n209), .B2(new_n767), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT97), .Z(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(new_n247), .B2(new_n296), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n688), .A2(new_n416), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n771), .A2(G355), .B1(new_n267), .B2(new_n688), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n765), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n311), .A2(G179), .A3(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n210), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n210), .A2(G179), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n777), .A2(G190), .A3(G200), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n776), .A2(G97), .B1(new_n779), .B2(G87), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n210), .A2(new_n578), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G200), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G190), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n777), .A2(new_n311), .A3(G200), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n780), .B1(new_n207), .B2(new_n784), .C1(new_n203), .C2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G190), .A2(G200), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n777), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G159), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n788), .A2(KEYINPUT32), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(KEYINPUT32), .B1(new_n788), .B2(new_n789), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n782), .A2(new_n311), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n791), .B1(new_n793), .B2(new_n335), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n781), .A2(new_n787), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n781), .A2(G190), .A3(new_n365), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n261), .B1(new_n795), .B2(new_n224), .C1(new_n206), .C2(new_n796), .ZN(new_n797));
  NOR4_X1   g0597(.A1(new_n786), .A2(new_n790), .A3(new_n794), .A4(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G317), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(KEYINPUT33), .ZN(new_n800));
  OR2_X1    g0600(.A1(new_n799), .A2(KEYINPUT33), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n783), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G294), .ZN(new_n803));
  INV_X1    g0603(.A(G326), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n802), .B1(new_n803), .B2(new_n775), .C1(new_n804), .C2(new_n793), .ZN(new_n805));
  INV_X1    g0605(.A(new_n796), .ZN(new_n806));
  INV_X1    g0606(.A(new_n788), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n806), .A2(G322), .B1(new_n807), .B2(G329), .ZN(new_n808));
  INV_X1    g0608(.A(G311), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n808), .B(new_n416), .C1(new_n809), .C2(new_n795), .ZN(new_n810));
  INV_X1    g0610(.A(G283), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n811), .A2(new_n785), .B1(new_n778), .B2(new_n504), .ZN(new_n812));
  NOR3_X1   g0612(.A1(new_n805), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n798), .A2(new_n813), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n755), .B(new_n773), .C1(new_n763), .C2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n762), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n749), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n759), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT98), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G396));
  INV_X1    g0620(.A(new_n763), .ZN(new_n821));
  INV_X1    g0621(.A(new_n795), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n806), .A2(G143), .B1(new_n822), .B2(G159), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n792), .A2(G137), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n823), .B(new_n824), .C1(new_n338), .C2(new_n784), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT34), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n785), .A2(new_n207), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n416), .B(new_n829), .C1(G132), .C2(new_n807), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n776), .A2(G58), .B1(new_n779), .B2(G50), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n827), .A2(new_n828), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n811), .A2(new_n784), .B1(new_n793), .B2(new_n504), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(G107), .B2(new_n779), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n776), .A2(G97), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n796), .A2(new_n803), .B1(new_n788), .B2(new_n809), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n261), .B(new_n836), .C1(G116), .C2(new_n822), .ZN(new_n837));
  INV_X1    g0637(.A(new_n785), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(G87), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n834), .A2(new_n835), .A3(new_n837), .A4(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n821), .B1(new_n832), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n763), .A2(new_n760), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n755), .B(new_n841), .C1(new_n224), .C2(new_n842), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT99), .Z(new_n844));
  OR2_X1    g0644(.A1(new_n400), .A2(new_n669), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n390), .A2(new_n669), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n403), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n400), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n844), .B1(new_n761), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n404), .A2(new_n670), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(new_n705), .B2(new_n710), .ZN(new_n853));
  INV_X1    g0653(.A(new_n711), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n849), .B(KEYINPUT100), .Z(new_n855));
  AOI21_X1  g0655(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n754), .B1(new_n857), .B2(new_n733), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n857), .A2(new_n733), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n851), .B1(new_n859), .B2(new_n860), .ZN(G384));
  NOR2_X1   g0661(.A1(new_n751), .A2(new_n213), .ZN(new_n862));
  INV_X1    g0662(.A(G330), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n727), .A2(new_n669), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n729), .B1(new_n864), .B2(KEYINPUT106), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n727), .A2(KEYINPUT106), .A3(new_n669), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n731), .B(new_n714), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n492), .B(new_n669), .C1(new_n476), .C2(new_n629), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n492), .A2(new_n669), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n466), .A2(new_n470), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT14), .ZN(new_n871));
  OAI21_X1  g0671(.A(G169), .B1(new_n464), .B2(new_n465), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT77), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n870), .B1(new_n874), .B2(new_n474), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n497), .B(new_n869), .C1(new_n875), .C2(new_n494), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n849), .B1(new_n868), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n207), .B1(new_n415), .B2(new_n417), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n406), .B1(new_n413), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(new_n423), .A3(new_n254), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n426), .ZN(new_n881));
  INV_X1    g0681(.A(new_n667), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n456), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n881), .A2(new_n437), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n883), .A2(new_n886), .A3(KEYINPUT37), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n427), .A2(new_n882), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n442), .A2(new_n888), .A3(new_n451), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT37), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n887), .A2(new_n451), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT38), .B1(new_n885), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n883), .B1(new_n445), .B2(new_n455), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n889), .A2(new_n890), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n883), .A2(new_n886), .A3(new_n451), .A4(KEYINPUT37), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR3_X1   g0697(.A1(new_n893), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n867), .B(new_n877), .C1(new_n892), .C2(new_n898), .ZN(new_n899));
  XOR2_X1   g0699(.A(KEYINPUT105), .B(KEYINPUT40), .Z(new_n900));
  AND2_X1   g0700(.A1(new_n867), .A2(new_n877), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  XOR2_X1   g0702(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n903));
  AOI21_X1  g0703(.A(new_n667), .B1(new_n424), .B2(new_n426), .ZN(new_n904));
  OAI21_X1  g0704(.A(KEYINPUT37), .B1(new_n904), .B2(KEYINPUT104), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n889), .B(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n888), .B1(new_n455), .B2(new_n632), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n453), .A2(new_n454), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT18), .B1(new_n427), .B2(new_n437), .ZN(new_n910));
  AOI221_X4 g0710(.A(new_n443), .B1(new_n435), .B2(new_n436), .C1(new_n424), .C2(new_n426), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n910), .B1(new_n911), .B2(KEYINPUT79), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n909), .B1(new_n912), .B2(new_n440), .ZN(new_n913));
  OAI211_X1 g0713(.A(KEYINPUT38), .B(new_n891), .C1(new_n913), .C2(new_n883), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n902), .B1(new_n908), .B2(new_n914), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n899), .A2(new_n900), .B1(new_n901), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT107), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n867), .A2(new_n499), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n863), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n918), .B2(new_n917), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n868), .A2(new_n876), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n852), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n650), .B2(new_n661), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT101), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n845), .B(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n924), .A2(KEYINPUT102), .A3(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT102), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n853), .B2(new_n926), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n922), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n894), .B1(new_n893), .B2(new_n897), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n914), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n908), .A2(new_n914), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT39), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n476), .A2(new_n492), .A3(new_n670), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n932), .A2(new_n914), .A3(KEYINPUT39), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n444), .A2(new_n438), .A3(new_n667), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n934), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AOI211_X1 g0743(.A(KEYINPUT29), .B(new_n669), .C1(new_n705), .C2(new_n710), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n712), .B1(new_n742), .B2(new_n670), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n499), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n634), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n943), .B(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n862), .B1(new_n920), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n948), .B2(new_n920), .ZN(new_n950));
  NOR3_X1   g0750(.A1(new_n211), .A2(new_n210), .A3(new_n267), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n559), .A2(new_n563), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT35), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n953), .B2(new_n952), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT36), .Z(new_n956));
  AOI211_X1 g0756(.A(new_n224), .B(new_n209), .C1(new_n227), .C2(G58), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n207), .A2(G50), .ZN(new_n958));
  OAI211_X1 g0758(.A(G1), .B(new_n279), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n950), .A2(new_n956), .A3(new_n959), .ZN(G367));
  OAI22_X1  g0760(.A1(new_n784), .A2(new_n789), .B1(new_n778), .B2(new_n206), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(G68), .B2(new_n776), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n796), .A2(new_n338), .B1(new_n795), .B2(new_n335), .ZN(new_n963));
  XNOR2_X1  g0763(.A(KEYINPUT114), .B(G137), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n261), .B1(new_n788), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n792), .A2(G143), .B1(new_n838), .B2(G77), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n962), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n795), .A2(new_n811), .B1(new_n788), .B2(new_n799), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n261), .B(new_n969), .C1(G303), .C2(new_n806), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n554), .A2(new_n776), .B1(new_n783), .B2(G294), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n792), .A2(G311), .B1(new_n838), .B2(G97), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT46), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n778), .B2(new_n267), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n970), .A2(new_n971), .A3(new_n972), .A4(new_n974), .ZN(new_n975));
  NOR3_X1   g0775(.A1(new_n778), .A2(new_n973), .A3(new_n267), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT113), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n968), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT47), .Z(new_n979));
  NOR2_X1   g0779(.A1(new_n979), .A2(new_n821), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n669), .A2(new_n638), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n659), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n655), .B2(new_n981), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n983), .A2(new_n816), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n764), .B1(new_n216), .B2(new_n380), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(new_n766), .B2(new_n241), .ZN(new_n986));
  NOR4_X1   g0786(.A1(new_n980), .A2(new_n755), .A3(new_n984), .A4(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT115), .Z(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n983), .A2(KEYINPUT43), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n571), .B(new_n580), .C1(new_n566), .C2(new_n670), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n679), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n669), .B1(new_n993), .B2(new_n580), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT109), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n648), .A2(new_n669), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n995), .B1(new_n683), .B2(new_n998), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n682), .A2(new_n329), .A3(new_n997), .A4(KEYINPUT109), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n994), .B1(new_n1001), .B2(KEYINPUT42), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(KEYINPUT42), .B2(new_n1001), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT108), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n983), .A2(KEYINPUT43), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1004), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n991), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n681), .A2(new_n998), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(KEYINPUT108), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1012), .A2(new_n990), .A3(new_n1006), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1009), .A2(new_n1010), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT110), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1009), .A2(new_n1013), .A3(KEYINPUT110), .A4(new_n1010), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n1007), .A2(new_n1008), .A3(new_n991), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n990), .B1(new_n1012), .B2(new_n1006), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n1019), .A2(new_n1020), .B1(new_n681), .B2(new_n998), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n692), .B(KEYINPUT41), .Z(new_n1022));
  OAI21_X1  g0822(.A(new_n683), .B1(new_n680), .B2(new_n682), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n757), .A2(new_n758), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT112), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1023), .A2(new_n676), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n757), .A2(new_n1023), .A3(KEYINPUT112), .A4(new_n758), .ZN(new_n1028));
  AND3_X1   g0828(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n681), .ZN(new_n1030));
  OAI21_X1  g0830(.A(KEYINPUT111), .B1(new_n686), .B2(new_n997), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT111), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n685), .A2(new_n1032), .A3(new_n998), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1031), .A2(KEYINPUT44), .A3(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n686), .A2(KEYINPUT45), .A3(new_n997), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT45), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n685), .B2(new_n998), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(KEYINPUT44), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1030), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1040), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1042), .A2(new_n681), .A3(new_n1038), .A4(new_n1034), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1029), .A2(new_n747), .A3(new_n1041), .A4(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1022), .B1(new_n1044), .B2(new_n747), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1021), .B1(new_n1045), .B2(new_n753), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n989), .B1(new_n1018), .B2(new_n1046), .ZN(G387));
  OR2_X1    g0847(.A1(new_n680), .A2(new_n816), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n694), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n771), .A2(new_n1049), .B1(new_n203), .B2(new_n688), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT116), .Z(new_n1051));
  NAND2_X1  g0851(.A1(new_n238), .A2(new_n767), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n766), .ZN(new_n1053));
  AOI211_X1 g0853(.A(G45), .B(new_n1049), .C1(G68), .C2(G77), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n337), .A2(G50), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(KEYINPUT117), .B(KEYINPUT50), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1055), .B(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1053), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1051), .B1(new_n1052), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n754), .B1(new_n1059), .B2(new_n765), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n806), .A2(G317), .B1(new_n822), .B2(G303), .ZN(new_n1061));
  INV_X1    g0861(.A(G322), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1061), .B1(new_n793), .B2(new_n1062), .C1(new_n809), .C2(new_n784), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT48), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n811), .B2(new_n775), .C1(new_n803), .C2(new_n778), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1068), .A2(KEYINPUT49), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n416), .B1(new_n788), .B2(new_n804), .C1(new_n267), .C2(new_n785), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(KEYINPUT49), .B2(new_n1068), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n795), .A2(new_n207), .B1(new_n788), .B2(new_n338), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n416), .B(new_n1073), .C1(G50), .C2(new_n806), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n779), .A2(G77), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n337), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n589), .A2(new_n776), .B1(new_n783), .B2(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n792), .A2(G159), .B1(new_n838), .B2(G97), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1074), .A2(new_n1075), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1072), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1060), .B1(new_n1080), .B2(new_n763), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1029), .A2(new_n753), .B1(new_n1048), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1029), .A2(new_n747), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n692), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1029), .A2(new_n747), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1082), .B1(new_n1084), .B2(new_n1085), .ZN(G393));
  NAND3_X1  g0886(.A1(new_n1041), .A2(new_n1043), .A3(KEYINPUT118), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT118), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1030), .B(new_n1088), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1087), .A2(new_n1083), .A3(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1090), .A2(new_n692), .A3(new_n1044), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n998), .A2(new_n762), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n251), .A2(new_n1053), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n764), .B1(new_n202), .B2(new_n216), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n754), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n775), .A2(new_n224), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n1076), .B2(new_n822), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n335), .B2(new_n784), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT119), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(G150), .A2(new_n792), .B1(new_n806), .B2(G159), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT51), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n416), .B1(new_n807), .B2(G143), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1103), .B(new_n839), .C1(new_n409), .C2(new_n778), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n1100), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G317), .A2(new_n792), .B1(new_n806), .B2(G311), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT52), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n416), .B1(new_n788), .B2(new_n1062), .C1(new_n803), .C2(new_n795), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n784), .A2(new_n504), .B1(new_n785), .B2(new_n203), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n775), .A2(new_n267), .B1(new_n778), .B2(new_n811), .ZN(new_n1110));
  NOR4_X1   g0910(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  OR2_X1    g0911(.A1(new_n1105), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1096), .B1(new_n1112), .B2(new_n763), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1092), .A2(new_n753), .B1(new_n1093), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1091), .A2(new_n1114), .ZN(G390));
  AOI21_X1  g0915(.A(new_n761), .B1(new_n937), .B2(new_n940), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n842), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(G97), .A2(new_n822), .B1(new_n807), .B2(G294), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1118), .B(new_n416), .C1(new_n267), .C2(new_n796), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n829), .B(new_n1119), .C1(G87), .C2(new_n779), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n784), .A2(new_n392), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1097), .B(new_n1121), .C1(G283), .C2(new_n792), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n778), .A2(new_n338), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT53), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n784), .A2(new_n964), .B1(new_n335), .B2(new_n785), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n792), .A2(G128), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n789), .B2(new_n775), .ZN(new_n1127));
  INV_X1    g0927(.A(G125), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n261), .B1(new_n788), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(G132), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(KEYINPUT54), .B(G143), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n796), .A2(new_n1130), .B1(new_n795), .B2(new_n1131), .ZN(new_n1132));
  NOR4_X1   g0932(.A1(new_n1125), .A2(new_n1127), .A3(new_n1129), .A4(new_n1132), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1120), .A2(new_n1122), .B1(new_n1124), .B2(new_n1133), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n754), .B1(new_n1076), .B2(new_n1117), .C1(new_n1134), .C2(new_n821), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1116), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n937), .A2(new_n940), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n931), .B2(new_n939), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n927), .B1(new_n743), .B2(new_n849), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n938), .B(new_n935), .C1(new_n1140), .C2(new_n922), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n732), .A2(G330), .A3(new_n850), .ZN(new_n1142));
  OR2_X1    g0942(.A1(new_n1142), .A2(new_n922), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n1138), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n714), .A2(new_n731), .ZN(new_n1145));
  AOI21_X1  g0945(.A(KEYINPUT106), .B1(new_n727), .B2(new_n669), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n866), .A2(new_n1146), .A3(KEYINPUT31), .ZN(new_n1147));
  OAI211_X1 g0947(.A(G330), .B(new_n877), .C1(new_n1145), .C2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(KEYINPUT120), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT120), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n867), .A2(new_n1150), .A3(G330), .A4(new_n877), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1144), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1136), .B1(new_n1154), .B2(new_n753), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1138), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n935), .A2(new_n938), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n921), .B2(new_n1139), .ZN(new_n1158));
  AOI21_X1  g0958(.A(KEYINPUT102), .B1(new_n924), .B2(new_n927), .ZN(new_n1159));
  NOR3_X1   g0959(.A1(new_n853), .A2(new_n929), .A3(new_n926), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n921), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n938), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1158), .B1(new_n1162), .B2(new_n1137), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1156), .B1(new_n1163), .B2(new_n1152), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1142), .A2(new_n922), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1149), .A2(new_n1151), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n928), .A2(new_n930), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n867), .A2(G330), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n922), .B1(new_n1169), .B2(new_n855), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1170), .A2(new_n1143), .A3(new_n1140), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n499), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n946), .B(new_n634), .C1(new_n1173), .C2(new_n1169), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n693), .B1(new_n1164), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1174), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1156), .B(new_n1178), .C1(new_n1163), .C2(new_n1152), .ZN(new_n1179));
  AOI21_X1  g0979(.A(KEYINPUT121), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1176), .B1(new_n1144), .B2(new_n1153), .ZN(new_n1181));
  AND4_X1   g0981(.A1(KEYINPUT121), .A2(new_n1181), .A3(new_n692), .A4(new_n1179), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1155), .B1(new_n1180), .B2(new_n1182), .ZN(G378));
  OAI21_X1  g0983(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n346), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1185), .A2(new_n667), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  OR3_X1    g0990(.A1(new_n1187), .A2(new_n1188), .A3(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1190), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n899), .A2(new_n900), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n901), .A2(new_n915), .ZN(new_n1195));
  AND4_X1   g0995(.A1(G330), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1193), .B1(new_n916), .B2(G330), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n943), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n934), .A2(new_n941), .A3(new_n942), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1194), .A2(new_n1195), .A3(G330), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1193), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n916), .A2(G330), .A3(new_n1193), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1199), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1198), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1201), .A2(new_n760), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n754), .B1(G50), .B2(new_n1117), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n784), .A2(new_n202), .B1(new_n785), .B2(new_n206), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G116), .B2(new_n792), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n416), .A2(new_n302), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G283), .B2(new_n807), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n806), .A2(G107), .B1(new_n822), .B2(new_n589), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n776), .A2(G68), .B1(new_n779), .B2(G77), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1209), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT58), .ZN(new_n1215));
  AOI21_X1  g1015(.A(G50), .B1(new_n255), .B2(new_n302), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1214), .A2(new_n1215), .B1(new_n1210), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT122), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1218), .A2(G124), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(G124), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n807), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1221), .A2(new_n255), .A3(new_n302), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n1128), .A2(new_n793), .B1(new_n784), .B2(new_n1130), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n806), .A2(G128), .B1(new_n822), .B2(G137), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n778), .B2(new_n1131), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1223), .B(new_n1225), .C1(G150), .C2(new_n776), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT59), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1222), .B1(new_n789), .B2(new_n785), .C1(new_n1226), .C2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1226), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1229), .A2(KEYINPUT59), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1217), .B1(new_n1215), .B2(new_n1214), .C1(new_n1228), .C2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1207), .B1(new_n1231), .B2(new_n763), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1205), .A2(new_n753), .B1(new_n1206), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT57), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(new_n1198), .B2(new_n1204), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1179), .A2(new_n1175), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n692), .ZN(new_n1238));
  AOI21_X1  g1038(.A(KEYINPUT57), .B1(new_n1236), .B2(new_n1205), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1233), .B1(new_n1238), .B2(new_n1239), .ZN(G375));
  INV_X1    g1040(.A(new_n1022), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1168), .A2(new_n1174), .A3(new_n1171), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1176), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n922), .A2(new_n760), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n267), .A2(new_n784), .B1(new_n793), .B2(new_n803), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(G97), .B2(new_n779), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n261), .B1(new_n807), .B2(G303), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n806), .A2(G283), .B1(new_n822), .B2(new_n554), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n776), .A2(new_n589), .B1(new_n838), .B2(G77), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n796), .A2(new_n964), .B1(new_n795), .B2(new_n338), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n416), .B(new_n1251), .C1(G128), .C2(new_n807), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n775), .A2(new_n335), .B1(new_n778), .B2(new_n789), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(G132), .B2(new_n792), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1131), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n783), .A2(new_n1255), .B1(new_n838), .B2(G58), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1252), .A2(new_n1254), .A3(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n821), .B1(new_n1250), .B2(new_n1257), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n755), .B(new_n1258), .C1(new_n207), .C2(new_n842), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n1172), .A2(new_n753), .B1(new_n1244), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1243), .A2(new_n1260), .ZN(G381));
  NAND3_X1  g1061(.A1(new_n1181), .A2(new_n692), .A3(new_n1179), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1262), .A2(new_n1155), .A3(KEYINPUT123), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT123), .B1(new_n1262), .B2(new_n1155), .ZN(new_n1264));
  OR2_X1    g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1205), .A2(new_n753), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1206), .A2(new_n1232), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1236), .A2(new_n1205), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1234), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n693), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1268), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1265), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(G387), .ZN(new_n1274));
  INV_X1    g1074(.A(G381), .ZN(new_n1275));
  NOR4_X1   g1075(.A1(G390), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1273), .A2(new_n1274), .A3(new_n1275), .A4(new_n1276), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1277), .B(KEYINPUT124), .ZN(G407));
  INV_X1    g1078(.A(G213), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1279), .B1(new_n1273), .B2(new_n668), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G407), .A2(new_n1280), .ZN(G409));
  INV_X1    g1081(.A(KEYINPUT127), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT126), .ZN(new_n1283));
  INV_X1    g1083(.A(G390), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1283), .B1(G387), .B2(new_n1284), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(G393), .B(new_n819), .ZN(new_n1286));
  OR2_X1    g1086(.A1(new_n1045), .A2(new_n753), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1287), .A2(new_n1021), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1288));
  AOI21_X1  g1088(.A(G390), .B1(new_n1288), .B2(new_n989), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n989), .B(G390), .C1(new_n1018), .C2(new_n1046), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  OAI22_X1  g1091(.A1(new_n1285), .A2(new_n1286), .B1(new_n1289), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(G387), .A2(new_n1284), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1286), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1293), .A2(new_n1294), .A3(new_n1283), .A4(new_n1290), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1292), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT62), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1233), .B1(new_n1269), .B2(new_n1022), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1298), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1155), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT121), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1262), .A2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1177), .A2(KEYINPUT121), .A3(new_n1179), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1300), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1299), .B1(G375), .B2(new_n1304), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1279), .A2(G343), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT60), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1242), .A2(new_n1308), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1168), .A2(new_n1171), .A3(new_n1174), .A4(KEYINPUT60), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1309), .A2(new_n1176), .A3(new_n692), .A4(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1260), .ZN(new_n1312));
  INV_X1    g1112(.A(G384), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1311), .A2(G384), .A3(new_n1260), .ZN(new_n1315));
  AND2_X1   g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  AND4_X1   g1116(.A1(new_n1297), .A2(new_n1305), .A3(new_n1307), .A4(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1272), .A2(G378), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1306), .B1(new_n1318), .B2(new_n1299), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1297), .B1(new_n1319), .B2(new_n1316), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1317), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1319), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT125), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1306), .A2(G2897), .ZN(new_n1324));
  AND3_X1   g1124(.A1(new_n1316), .A2(new_n1323), .A3(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1324), .B1(new_n1316), .B2(new_n1323), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1316), .A2(new_n1323), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1325), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(KEYINPUT61), .B1(new_n1322), .B2(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1296), .B1(new_n1321), .B2(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1319), .A2(KEYINPUT63), .A3(new_n1316), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1296), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT61), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1316), .A2(new_n1323), .A3(new_n1324), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1333), .B1(new_n1336), .B2(new_n1319), .ZN(new_n1337));
  AOI21_X1  g1137(.A(KEYINPUT63), .B1(new_n1319), .B2(new_n1316), .ZN(new_n1338));
  NOR3_X1   g1138(.A1(new_n1332), .A2(new_n1337), .A3(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1282), .B1(new_n1330), .B2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1338), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1329), .A2(new_n1341), .A3(new_n1296), .A4(new_n1331), .ZN(new_n1342));
  NOR3_X1   g1142(.A1(new_n1337), .A2(new_n1320), .A3(new_n1317), .ZN(new_n1343));
  OAI211_X1 g1143(.A(new_n1342), .B(KEYINPUT127), .C1(new_n1343), .C2(new_n1296), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1340), .A2(new_n1344), .ZN(G405));
  NOR2_X1   g1145(.A1(G375), .A2(new_n1304), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1346), .B1(G375), .B2(new_n1265), .ZN(new_n1347));
  XNOR2_X1  g1147(.A(new_n1296), .B(new_n1347), .ZN(new_n1348));
  XNOR2_X1  g1148(.A(new_n1348), .B(new_n1316), .ZN(G402));
endmodule


