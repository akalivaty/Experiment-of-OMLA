//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 1 1 1 1 0 0 0 1 0 0 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 0 0 0 0 1 0 1 0 0 1 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1246, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  INV_X1    g0002(.A(G58), .ZN(new_n203));
  INV_X1    g0003(.A(G68), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NOR3_X1   g0005(.A1(new_n202), .A2(G77), .A3(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT65), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  INV_X1    g0015(.A(G13), .ZN(new_n216));
  OAI21_X1  g0016(.A(KEYINPUT66), .B1(new_n208), .B2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT66), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n218), .A2(G1), .A3(G13), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n221), .A2(new_n209), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n205), .A2(G50), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n226));
  INV_X1    g0026(.A(G238), .ZN(new_n227));
  INV_X1    g0027(.A(G77), .ZN(new_n228));
  INV_X1    g0028(.A(G244), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n226), .B1(new_n204), .B2(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT67), .ZN(new_n231));
  AOI22_X1  g0031(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT68), .ZN(new_n233));
  AOI22_X1  g0033(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g0035(.A(new_n211), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  OAI211_X1 g0036(.A(new_n215), .B(new_n225), .C1(KEYINPUT1), .C2(new_n236), .ZN(new_n237));
  AOI21_X1  g0037(.A(new_n237), .B1(KEYINPUT1), .B2(new_n236), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XOR2_X1   g0040(.A(KEYINPUT2), .B(G226), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G264), .B(G270), .Z(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G358));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT69), .B(G50), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(KEYINPUT88), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT70), .B(G1698), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n256), .A2(G250), .B1(G257), .B2(G1698), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT76), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT76), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n259), .A2(new_n261), .A3(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G294), .ZN(new_n266));
  OAI22_X1  g0066(.A1(new_n257), .A2(new_n265), .B1(new_n263), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  AND2_X1   g0068(.A1(new_n220), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n268), .A2(G1), .A3(G13), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n208), .A2(G45), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT5), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n272), .B1(new_n273), .B2(G41), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(KEYINPUT80), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT80), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT5), .ZN(new_n277));
  AOI21_X1  g0077(.A(G41), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT81), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n274), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI211_X1 g0080(.A(KEYINPUT81), .B(G41), .C1(new_n275), .C2(new_n277), .ZN(new_n281));
  OAI211_X1 g0081(.A(G264), .B(new_n271), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  AND3_X1   g0082(.A1(new_n270), .A2(G179), .A3(new_n282), .ZN(new_n283));
  OR2_X1    g0083(.A1(new_n278), .A2(new_n279), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n278), .A2(new_n279), .ZN(new_n285));
  AND2_X1   g0085(.A1(new_n271), .A2(G274), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n284), .A2(new_n285), .A3(new_n274), .A4(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n270), .A2(new_n282), .A3(new_n287), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n283), .A2(new_n287), .B1(new_n288), .B2(G169), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n217), .A2(new_n219), .A3(new_n290), .A4(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n263), .A2(G1), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G107), .ZN(new_n295));
  INV_X1    g0095(.A(G107), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n208), .A2(new_n296), .A3(G13), .A4(G20), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n297), .A2(KEYINPUT86), .A3(KEYINPUT25), .ZN(new_n298));
  XNOR2_X1  g0098(.A(KEYINPUT86), .B(KEYINPUT25), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n299), .A2(new_n297), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n295), .A2(KEYINPUT87), .A3(new_n298), .A4(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT87), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n292), .A2(new_n296), .A3(new_n293), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(new_n298), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(KEYINPUT85), .B1(new_n209), .B2(G107), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT23), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT23), .ZN(new_n309));
  OAI211_X1 g0109(.A(KEYINPUT85), .B(new_n309), .C1(new_n209), .C2(G107), .ZN(new_n310));
  INV_X1    g0110(.A(G116), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n263), .A2(new_n311), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n308), .A2(new_n310), .B1(new_n209), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT22), .ZN(new_n314));
  INV_X1    g0114(.A(G87), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n262), .A2(new_n209), .A3(new_n264), .A4(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n258), .A2(G33), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n264), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n209), .A2(G87), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n314), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n313), .A2(new_n317), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT24), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n217), .A2(new_n219), .A3(new_n290), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n313), .A2(new_n317), .A3(KEYINPUT24), .A4(new_n321), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n306), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n255), .B1(new_n289), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n288), .A2(G200), .ZN(new_n330));
  INV_X1    g0130(.A(G190), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n328), .B(new_n330), .C1(new_n331), .C2(new_n288), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n288), .A2(G169), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n270), .A2(new_n282), .A3(G179), .A4(new_n287), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n306), .A2(new_n327), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(KEYINPUT88), .A3(new_n336), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n329), .A2(new_n332), .A3(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n291), .A2(G77), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n209), .A2(G1), .ZN(new_n340));
  NOR3_X1   g0140(.A1(new_n292), .A2(new_n228), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G20), .A2(G77), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n209), .A2(new_n263), .ZN(new_n343));
  XNOR2_X1  g0143(.A(KEYINPUT8), .B(G58), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n315), .A2(KEYINPUT15), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT15), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G87), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n263), .A2(G20), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  OAI221_X1 g0151(.A(new_n342), .B1(new_n343), .B2(new_n344), .C1(new_n349), .C2(new_n351), .ZN(new_n352));
  AOI211_X1 g0152(.A(new_n339), .B(new_n341), .C1(new_n352), .C2(new_n325), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT3), .B(G33), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n354), .A2(new_n256), .A3(G232), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(G238), .A3(G1698), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n319), .A2(G107), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT71), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT71), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n355), .A2(new_n356), .A3(new_n360), .A4(new_n357), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(new_n269), .A3(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n364), .A2(new_n271), .A3(G274), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n271), .A2(new_n363), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n366), .B1(G244), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n362), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G169), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n353), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT72), .ZN(new_n372));
  OR2_X1    g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n372), .ZN(new_n374));
  INV_X1    g0174(.A(G179), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n362), .A2(new_n375), .A3(new_n368), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n339), .B1(new_n352), .B2(new_n325), .ZN(new_n378));
  INV_X1    g0178(.A(new_n341), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n380), .B1(new_n369), .B2(G200), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(new_n331), .B2(new_n369), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n383), .B(KEYINPUT73), .ZN(new_n384));
  INV_X1    g0184(.A(new_n292), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n344), .A2(new_n340), .ZN(new_n386));
  INV_X1    g0186(.A(new_n291), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n385), .A2(new_n386), .B1(new_n387), .B2(new_n344), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n325), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT77), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G58), .A2(G68), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n209), .B1(new_n205), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G159), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n343), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n391), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n392), .ZN(new_n397));
  NOR2_X1   g0197(.A1(G58), .A2(G68), .ZN(new_n398));
  OAI21_X1  g0198(.A(G20), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(G20), .A2(G33), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(G159), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(KEYINPUT77), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n396), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(G20), .B1(new_n262), .B2(new_n264), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT7), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n204), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n264), .ZN(new_n407));
  XNOR2_X1  g0207(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n407), .B1(new_n408), .B2(G33), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT7), .B1(new_n409), .B2(G20), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n403), .B1(new_n406), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n390), .B1(new_n411), .B2(KEYINPUT16), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT16), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n405), .A2(G20), .ZN(new_n414));
  AOI21_X1  g0214(.A(G33), .B1(new_n259), .B2(new_n261), .ZN(new_n415));
  INV_X1    g0215(.A(new_n318), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n405), .B1(new_n354), .B2(G20), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n204), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n413), .B1(new_n419), .B2(new_n403), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n389), .B1(new_n412), .B2(new_n420), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n367), .A2(G232), .B1(new_n286), .B2(new_n364), .ZN(new_n422));
  NAND2_X1  g0222(.A1(G226), .A2(G1698), .ZN(new_n423));
  INV_X1    g0223(.A(G1698), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT70), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT70), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(G1698), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(G223), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n423), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n430), .A2(new_n409), .B1(G33), .B2(G87), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n220), .A2(new_n268), .ZN(new_n432));
  OAI211_X1 g0232(.A(G179), .B(new_n422), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n367), .A2(G232), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n365), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n256), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n436));
  OAI22_X1  g0236(.A1(new_n436), .A2(new_n265), .B1(new_n263), .B2(new_n315), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n435), .B1(new_n437), .B2(new_n269), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n433), .B1(new_n438), .B2(new_n370), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT18), .B1(new_n421), .B2(new_n440), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n396), .A2(new_n402), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n265), .A2(new_n405), .A3(new_n209), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G68), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n404), .A2(new_n405), .ZN(new_n445));
  OAI211_X1 g0245(.A(KEYINPUT16), .B(new_n442), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n446), .A2(new_n325), .A3(new_n420), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n388), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT18), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(new_n449), .A3(new_n439), .ZN(new_n450));
  XNOR2_X1  g0250(.A(KEYINPUT78), .B(G190), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n451), .B(new_n422), .C1(new_n431), .C2(new_n432), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n438), .B2(G200), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n447), .A2(new_n388), .A3(new_n453), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n454), .A2(KEYINPUT17), .ZN(new_n455));
  XOR2_X1   g0255(.A(KEYINPUT79), .B(KEYINPUT17), .Z(new_n456));
  AND4_X1   g0256(.A1(new_n447), .A2(new_n453), .A3(new_n388), .A4(new_n456), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n441), .B(new_n450), .C1(new_n455), .C2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n209), .B1(new_n201), .B2(new_n398), .ZN(new_n460));
  INV_X1    g0260(.A(G150), .ZN(new_n461));
  OAI22_X1  g0261(.A1(new_n344), .A2(new_n351), .B1(new_n461), .B2(new_n343), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n325), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n340), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n385), .A2(G50), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G50), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n387), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n463), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n354), .A2(G223), .A3(G1698), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n354), .A2(new_n256), .A3(G222), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n469), .B(new_n470), .C1(new_n228), .C2(new_n354), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n269), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n366), .B1(G226), .B2(new_n367), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n468), .B1(new_n475), .B2(G169), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n476), .B1(new_n375), .B2(new_n475), .ZN(new_n477));
  INV_X1    g0277(.A(new_n468), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n475), .A2(G190), .B1(new_n478), .B2(KEYINPUT9), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT9), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n474), .A2(G200), .B1(new_n468), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  OR2_X1    g0282(.A1(new_n482), .A2(KEYINPUT10), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(KEYINPUT10), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n477), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G200), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G97), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n425), .A2(new_n427), .A3(G226), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G232), .A2(G1698), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n319), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n269), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n367), .A2(G238), .B1(new_n286), .B2(new_n364), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT13), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT13), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n492), .A2(new_n496), .A3(new_n493), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n486), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n400), .A2(G50), .B1(G20), .B2(new_n204), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(new_n351), .B2(new_n228), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n325), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT75), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n500), .A2(KEYINPUT75), .A3(new_n325), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT11), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT11), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n503), .A2(new_n507), .A3(new_n504), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n292), .A2(new_n204), .A3(new_n340), .ZN(new_n509));
  OAI21_X1  g0309(.A(KEYINPUT12), .B1(new_n291), .B2(G68), .ZN(new_n510));
  OR3_X1    g0310(.A1(new_n291), .A2(KEYINPUT12), .A3(G68), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n506), .A2(new_n508), .A3(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n498), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT74), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n497), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n492), .A2(KEYINPUT74), .A3(new_n496), .A4(new_n493), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n516), .A2(new_n495), .A3(G190), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n492), .A2(new_n496), .A3(new_n493), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n496), .B1(new_n492), .B2(new_n493), .ZN(new_n521));
  OAI21_X1  g0321(.A(G169), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT14), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT14), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n524), .B(G169), .C1(new_n520), .C2(new_n521), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n516), .A2(new_n495), .A3(G179), .A4(new_n517), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n513), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n459), .A2(new_n485), .A3(new_n519), .A4(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n384), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n425), .A2(new_n427), .A3(G257), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G264), .A2(G1698), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n409), .A2(new_n533), .B1(G303), .B2(new_n319), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT83), .ZN(new_n535));
  NOR3_X1   g0335(.A1(new_n534), .A2(new_n535), .A3(new_n432), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n319), .A2(G303), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n256), .A2(G257), .B1(G264), .B2(G1698), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n537), .B1(new_n538), .B2(new_n265), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT83), .B1(new_n539), .B2(new_n269), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT20), .ZN(new_n542));
  AOI21_X1  g0342(.A(G20), .B1(G33), .B2(G283), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n263), .A2(G97), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT84), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n545), .B1(new_n543), .B2(new_n544), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n311), .A2(G20), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n325), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n542), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(G33), .A2(G283), .ZN(new_n553));
  INV_X1    g0353(.A(G97), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n553), .B(new_n209), .C1(G33), .C2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT84), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n546), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n557), .A2(KEYINPUT20), .A3(new_n325), .A4(new_n550), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n552), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n291), .A2(new_n311), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n294), .B2(new_n311), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(G270), .B(new_n271), .C1(new_n280), .C2(new_n281), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n563), .A2(new_n287), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n541), .A2(new_n562), .A3(G179), .A4(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n370), .B1(new_n559), .B2(new_n561), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT21), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n535), .B1(new_n534), .B2(new_n432), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n539), .A2(KEYINPUT83), .A3(new_n269), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n568), .A2(new_n569), .A3(new_n287), .A4(new_n563), .ZN(new_n570));
  AND3_X1   g0370(.A1(new_n566), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n567), .B1(new_n566), .B2(new_n570), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n565), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n486), .B1(new_n541), .B2(new_n564), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n570), .A2(new_n451), .ZN(new_n575));
  NOR3_X1   g0375(.A1(new_n574), .A2(new_n575), .A3(new_n562), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(G257), .B(new_n271), .C1(new_n280), .C2(new_n281), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n578), .A2(new_n287), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n428), .A2(new_n229), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT4), .B1(new_n409), .B2(new_n580), .ZN(new_n581));
  AND2_X1   g0381(.A1(KEYINPUT4), .A2(G244), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n354), .A2(new_n256), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n354), .A2(G250), .A3(G1698), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n583), .A2(new_n584), .A3(new_n553), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n269), .B1(new_n581), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n579), .A2(new_n375), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(new_n287), .A3(new_n578), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n370), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT6), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n554), .A2(new_n296), .ZN(new_n591));
  NOR2_X1   g0391(.A1(G97), .A2(G107), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n296), .A2(KEYINPUT6), .A3(G97), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI22_X1  g0395(.A1(new_n595), .A2(new_n209), .B1(new_n228), .B2(new_n343), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n296), .B1(new_n417), .B2(new_n418), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n325), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n291), .A2(G97), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n294), .B2(G97), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n587), .A2(new_n589), .A3(new_n601), .ZN(new_n602));
  OR2_X1    g0402(.A1(new_n272), .A2(G274), .ZN(new_n603));
  INV_X1    g0403(.A(G250), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n272), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n603), .A2(new_n271), .A3(new_n605), .ZN(new_n606));
  OAI22_X1  g0406(.A1(new_n428), .A2(new_n227), .B1(new_n229), .B2(new_n424), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n312), .B1(new_n607), .B2(new_n409), .ZN(new_n608));
  OAI211_X1 g0408(.A(G179), .B(new_n606), .C1(new_n608), .C2(new_n432), .ZN(new_n609));
  INV_X1    g0409(.A(new_n606), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n256), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n611));
  OAI22_X1  g0411(.A1(new_n611), .A2(new_n265), .B1(new_n263), .B2(new_n311), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n610), .B1(new_n612), .B2(new_n269), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n609), .B1(new_n613), .B2(new_n370), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT82), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n609), .B(KEYINPUT82), .C1(new_n613), .C2(new_n370), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n409), .A2(new_n209), .A3(G68), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT19), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n350), .A2(new_n619), .A3(G97), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n592), .A2(new_n315), .B1(new_n487), .B2(new_n209), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n620), .B1(new_n621), .B2(new_n619), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n390), .B1(new_n618), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n348), .A2(new_n291), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n294), .A2(new_n348), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n624), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n616), .A2(new_n617), .A3(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n598), .A2(new_n600), .ZN(new_n630));
  AOI21_X1  g0430(.A(G200), .B1(new_n579), .B2(new_n586), .ZN(new_n631));
  AND4_X1   g0431(.A1(new_n331), .A2(new_n586), .A3(new_n287), .A4(new_n578), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n613), .A2(new_n486), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n292), .A2(new_n315), .A3(new_n293), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n623), .A2(new_n625), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n613), .A2(G190), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  AND4_X1   g0438(.A1(new_n602), .A2(new_n629), .A3(new_n633), .A4(new_n638), .ZN(new_n639));
  AND4_X1   g0439(.A1(new_n338), .A2(new_n530), .A3(new_n577), .A4(new_n639), .ZN(G372));
  INV_X1    g0440(.A(new_n602), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n641), .A2(new_n629), .A3(KEYINPUT26), .A4(new_n638), .ZN(new_n642));
  INV_X1    g0442(.A(new_n628), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT89), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n614), .A2(new_n644), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n609), .B(KEYINPUT89), .C1(new_n613), .C2(new_n370), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n647), .A2(new_n648), .A3(new_n602), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n642), .B1(new_n649), .B2(KEYINPUT26), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n335), .A2(new_n336), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n651), .B(new_n565), .C1(new_n571), .C2(new_n572), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n633), .A2(new_n602), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n647), .A2(new_n648), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n652), .A2(new_n653), .A3(new_n654), .A4(new_n332), .ZN(new_n655));
  INV_X1    g0455(.A(new_n647), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n650), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n530), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n377), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n659), .A2(new_n519), .B1(new_n513), .B2(new_n527), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n457), .B1(KEYINPUT17), .B2(new_n454), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n441), .B(new_n450), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n483), .A2(new_n484), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n477), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n658), .A2(new_n664), .ZN(G369));
  NAND3_X1  g0465(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT27), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n668), .A2(new_n208), .A3(new_n209), .A4(G13), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n667), .A2(G213), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G343), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT90), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n562), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n577), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n573), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n674), .B1(new_n675), .B2(new_n673), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT91), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G330), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n336), .A2(new_n672), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n338), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT92), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n335), .A2(new_n336), .A3(new_n672), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n682), .B1(new_n681), .B2(new_n683), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n679), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n672), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n573), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n681), .A2(new_n683), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT92), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n691), .B1(new_n693), .B2(new_n684), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n651), .A2(new_n672), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n689), .A2(new_n696), .ZN(G399));
  INV_X1    g0497(.A(KEYINPUT93), .ZN(new_n698));
  INV_X1    g0498(.A(new_n212), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n698), .B1(new_n699), .B2(G41), .ZN(new_n700));
  INV_X1    g0500(.A(G41), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n212), .A2(KEYINPUT93), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n592), .A2(new_n315), .A3(new_n311), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n704), .A2(new_n208), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n706), .B1(new_n224), .B2(new_n704), .ZN(new_n707));
  XOR2_X1   g0507(.A(new_n707), .B(KEYINPUT28), .Z(new_n708));
  NAND3_X1  g0508(.A1(new_n653), .A2(new_n654), .A3(new_n332), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n329), .A2(new_n337), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n709), .B1(new_n710), .B2(new_n675), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT26), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n641), .A2(new_n629), .A3(new_n712), .A4(new_n638), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n656), .B(new_n713), .C1(new_n649), .C2(new_n712), .ZN(new_n714));
  OAI211_X1 g0514(.A(KEYINPUT29), .B(new_n690), .C1(new_n711), .C2(new_n714), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n657), .A2(new_n690), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n715), .B1(new_n716), .B2(KEYINPUT29), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n338), .A2(new_n577), .A3(new_n639), .A4(new_n690), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n541), .A2(new_n564), .A3(new_n586), .A4(new_n579), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n283), .A2(new_n613), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n612), .A2(new_n269), .ZN(new_n723));
  AOI21_X1  g0523(.A(G179), .B1(new_n723), .B2(new_n606), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n724), .A2(new_n288), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT94), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n725), .A2(new_n726), .A3(new_n570), .A4(new_n588), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n570), .A2(new_n588), .ZN(new_n728));
  AND4_X1   g0528(.A1(G179), .A2(new_n613), .A3(new_n282), .A4(new_n270), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n728), .A2(KEYINPUT30), .A3(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n570), .A2(new_n588), .A3(new_n288), .A4(new_n724), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(KEYINPUT94), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n722), .A2(new_n727), .A3(new_n730), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n672), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT31), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n722), .A2(new_n730), .A3(new_n731), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(KEYINPUT31), .A3(new_n672), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n718), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G330), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n717), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n708), .B1(new_n742), .B2(G1), .ZN(G364));
  XNOR2_X1  g0543(.A(new_n676), .B(KEYINPUT91), .ZN(new_n744));
  INV_X1    g0544(.A(G330), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(KEYINPUT95), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT95), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n679), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n216), .A2(G20), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n208), .B1(new_n750), .B2(G45), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n704), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n753), .B1(new_n744), .B2(new_n745), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n747), .A2(new_n749), .A3(new_n754), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n755), .A2(KEYINPUT96), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n221), .B1(G20), .B2(new_n370), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n209), .A2(new_n375), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n486), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n451), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT32), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n209), .A2(G190), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G179), .A2(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n394), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n762), .A2(new_n203), .B1(new_n763), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n768), .B1(new_n763), .B2(new_n767), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n486), .A2(G179), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n764), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n354), .B1(new_n771), .B2(new_n296), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n770), .A2(G20), .A3(G190), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n772), .B1(G87), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n759), .A2(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n451), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n760), .A2(G190), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n777), .A2(G50), .B1(new_n778), .B2(G77), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n209), .B1(new_n765), .B2(G190), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n554), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n776), .A2(G190), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n781), .B1(new_n782), .B2(G68), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n769), .A2(new_n775), .A3(new_n779), .A4(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G303), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n773), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G283), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n319), .B1(new_n771), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n766), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n786), .B(new_n788), .C1(G329), .C2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n761), .A2(G322), .ZN(new_n791));
  XNOR2_X1  g0591(.A(KEYINPUT33), .B(G317), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n777), .A2(G326), .B1(new_n782), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n780), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n778), .A2(G311), .B1(G294), .B2(new_n794), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n790), .A2(new_n791), .A3(new_n793), .A4(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n758), .B1(new_n784), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G13), .A2(G33), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(G20), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n757), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n212), .A2(new_n265), .ZN(new_n803));
  INV_X1    g0603(.A(G45), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n803), .B1(new_n804), .B2(new_n224), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(new_n250), .B2(new_n804), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n699), .A2(new_n319), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n807), .A2(G355), .B1(new_n311), .B2(new_n699), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n802), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n753), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n797), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n800), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n678), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n755), .A2(KEYINPUT96), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n756), .A2(new_n813), .A3(new_n814), .ZN(G396));
  NAND2_X1  g0615(.A1(new_n672), .A2(new_n380), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT99), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n816), .B(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n374), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n376), .B1(new_n371), .B2(new_n372), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n382), .B(new_n818), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n816), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n373), .A2(new_n374), .A3(new_n376), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n716), .B(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n740), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n826), .A2(new_n827), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n810), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n828), .B1(new_n830), .B2(KEYINPUT100), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(KEYINPUT100), .B2(new_n830), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n757), .A2(new_n798), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n753), .B1(G77), .B2(new_n834), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT97), .Z(new_n836));
  AOI22_X1  g0636(.A1(new_n777), .A2(G137), .B1(new_n778), .B2(G159), .ZN(new_n837));
  INV_X1    g0637(.A(G143), .ZN(new_n838));
  INV_X1    g0638(.A(new_n782), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n837), .B1(new_n838), .B2(new_n762), .C1(new_n461), .C2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT34), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n771), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(G68), .ZN(new_n844));
  INV_X1    g0644(.A(G132), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n844), .B1(new_n466), .B2(new_n773), .C1(new_n845), .C2(new_n766), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n265), .B(new_n846), .C1(G58), .C2(new_n794), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n840), .A2(new_n841), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n777), .A2(G303), .B1(new_n782), .B2(G283), .ZN(new_n850));
  INV_X1    g0650(.A(new_n778), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n850), .B1(new_n311), .B2(new_n851), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT98), .Z(new_n853));
  AOI21_X1  g0653(.A(new_n781), .B1(new_n761), .B2(G294), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n774), .A2(G107), .B1(new_n789), .B2(G311), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n354), .B1(new_n843), .B2(G87), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n842), .A2(new_n849), .B1(new_n853), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n836), .B1(new_n858), .B2(new_n757), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n824), .B2(new_n799), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n832), .A2(new_n860), .ZN(G384));
  NOR3_X1   g0661(.A1(new_n223), .A2(new_n228), .A3(new_n397), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT102), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n862), .A2(new_n863), .B1(G68), .B2(new_n201), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n863), .B2(new_n862), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n865), .A2(G1), .A3(new_n216), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT103), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT36), .ZN(new_n868));
  INV_X1    g0668(.A(new_n595), .ZN(new_n869));
  OAI211_X1 g0669(.A(G116), .B(new_n222), .C1(new_n869), .C2(KEYINPUT35), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n870), .A2(KEYINPUT101), .B1(KEYINPUT35), .B2(new_n869), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(KEYINPUT101), .B2(new_n870), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n867), .B1(new_n868), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n868), .B2(new_n872), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT39), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n442), .B1(new_n444), .B2(new_n445), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n413), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n389), .B1(new_n412), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n670), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n441), .A2(new_n450), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n880), .B1(new_n661), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n454), .B1(new_n878), .B2(new_n879), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n878), .A2(new_n440), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT37), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n448), .A2(new_n439), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n448), .A2(new_n670), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n886), .A2(new_n887), .A3(new_n888), .A4(new_n454), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n882), .A2(KEYINPUT38), .A3(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n887), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n458), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n886), .A2(new_n887), .A3(new_n454), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT37), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n889), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT38), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n875), .B1(new_n891), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT38), .B1(new_n882), .B2(new_n890), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n882), .A2(KEYINPUT38), .A3(new_n890), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n900), .A2(KEYINPUT39), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n528), .A2(new_n672), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n898), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n881), .A2(new_n879), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n657), .A2(new_n690), .A3(new_n824), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n659), .A2(new_n690), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n514), .A2(new_n518), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n513), .B(new_n672), .C1(new_n909), .C2(new_n527), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n513), .A2(new_n672), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n528), .A2(new_n519), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n908), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n914), .A2(KEYINPUT104), .ZN(new_n915));
  INV_X1    g0715(.A(new_n913), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n906), .B2(new_n907), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT104), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n917), .A2(new_n918), .B1(new_n891), .B2(new_n899), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n904), .B(new_n905), .C1(new_n915), .C2(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n530), .B(new_n715), .C1(KEYINPUT29), .C2(new_n716), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n921), .A2(new_n664), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n920), .B(new_n922), .Z(new_n923));
  OAI21_X1  g0723(.A(KEYINPUT105), .B1(new_n891), .B2(new_n897), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n528), .A2(new_n519), .A3(new_n911), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n911), .B1(new_n528), .B2(new_n519), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n824), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n733), .A2(KEYINPUT31), .A3(new_n672), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT31), .B1(new_n733), .B2(new_n672), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n927), .B1(new_n930), .B2(new_n718), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT105), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n458), .A2(new_n892), .B1(new_n895), .B2(new_n889), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n901), .B(new_n932), .C1(new_n933), .C2(KEYINPUT38), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n924), .A2(new_n931), .A3(KEYINPUT40), .A4(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n733), .A2(KEYINPUT31), .A3(new_n672), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n718), .A2(new_n736), .A3(new_n936), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n910), .A2(new_n912), .B1(new_n821), .B2(new_n823), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n937), .B(new_n938), .C1(new_n891), .C2(new_n899), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT40), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n935), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n530), .A2(new_n937), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n944), .A2(G330), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n923), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n208), .B2(new_n750), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n923), .A2(new_n946), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n874), .B1(new_n948), .B2(new_n949), .ZN(G367));
  INV_X1    g0750(.A(KEYINPUT42), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n633), .A2(new_n602), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n601), .B2(new_n672), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n641), .A2(new_n672), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n694), .A2(new_n951), .A3(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT106), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n957), .B(new_n958), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n954), .A2(new_n710), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n672), .B1(new_n960), .B2(new_n602), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n694), .A2(new_n956), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n961), .B1(new_n962), .B2(KEYINPUT42), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n690), .A2(new_n636), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n656), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(new_n654), .B2(new_n964), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n959), .A2(new_n963), .B1(KEYINPUT43), .B2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT43), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n956), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n689), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n959), .A2(new_n969), .A3(new_n966), .A4(new_n963), .ZN(new_n974));
  AND3_X1   g0774(.A1(new_n971), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n973), .B1(new_n971), .B2(new_n974), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n703), .B(KEYINPUT41), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n573), .B(new_n690), .C1(new_n685), .C2(new_n686), .ZN(new_n979));
  INV_X1    g0779(.A(new_n695), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n979), .A2(new_n980), .A3(new_n956), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(KEYINPUT107), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT107), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n696), .A2(new_n983), .A3(new_n956), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n982), .A2(new_n984), .A3(KEYINPUT45), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT44), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n696), .B2(new_n956), .ZN(new_n987));
  OAI211_X1 g0787(.A(KEYINPUT44), .B(new_n972), .C1(new_n694), .C2(new_n695), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n985), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(KEYINPUT45), .B1(new_n982), .B2(new_n984), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n688), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n687), .A2(new_n691), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n979), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n747), .A2(new_n749), .A3(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n746), .A2(new_n979), .A3(new_n993), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n995), .A2(new_n742), .A3(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n982), .A2(new_n984), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT45), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n1001), .A2(new_n689), .A3(new_n989), .A4(new_n985), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n992), .A2(new_n998), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n978), .B1(new_n1003), .B2(new_n742), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n977), .B1(new_n1004), .B2(new_n752), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n801), .B1(new_n212), .B2(new_n349), .C1(new_n245), .C2(new_n803), .ZN(new_n1006));
  AND2_X1   g0806(.A1(new_n1006), .A2(new_n753), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n771), .A2(new_n554), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n409), .B(new_n1008), .C1(G317), .C2(new_n789), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT108), .Z(new_n1010));
  NAND2_X1  g0810(.A1(new_n774), .A2(G116), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT46), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n778), .A2(G283), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n761), .A2(G303), .B1(new_n782), .B2(G294), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n777), .A2(G311), .B1(G107), .B2(new_n794), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n777), .A2(G143), .B1(G68), .B2(new_n794), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1017), .B1(new_n394), .B2(new_n839), .C1(new_n201), .C2(new_n851), .ZN(new_n1018));
  INV_X1    g0818(.A(G137), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n773), .A2(new_n203), .B1(new_n766), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(G150), .B2(new_n761), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n354), .B1(new_n771), .B2(new_n228), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT109), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1021), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n1010), .A2(new_n1016), .B1(new_n1018), .B2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1007), .B1(new_n1029), .B2(new_n758), .C1(new_n967), .C2(new_n812), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1005), .A2(new_n1030), .ZN(G387));
  NAND3_X1  g0831(.A1(new_n995), .A2(new_n752), .A3(new_n996), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n777), .A2(G322), .B1(new_n782), .B2(G311), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n761), .A2(G317), .B1(new_n778), .B2(G303), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1035), .A2(KEYINPUT48), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(KEYINPUT48), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n774), .A2(G294), .B1(new_n794), .B2(G283), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT49), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1041), .A2(KEYINPUT113), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(KEYINPUT113), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n843), .A2(G116), .B1(new_n789), .B2(G326), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1042), .A2(new_n1043), .A3(new_n265), .A4(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n773), .A2(new_n228), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1008), .B(new_n1046), .C1(G150), .C2(new_n789), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n777), .A2(G159), .B1(new_n778), .B2(G68), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n344), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n761), .A2(G50), .B1(new_n782), .B2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n349), .A2(new_n780), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1051), .A2(new_n265), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1047), .A2(new_n1048), .A3(new_n1050), .A4(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n758), .B1(new_n1045), .B2(new_n1053), .ZN(new_n1054));
  NOR3_X1   g0854(.A1(new_n685), .A2(new_n686), .A3(new_n812), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n807), .A2(new_n705), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(G107), .B2(new_n212), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n803), .B1(new_n242), .B2(G45), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n804), .B1(new_n204), .B2(new_n228), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n344), .A2(G50), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1059), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n705), .B(KEYINPUT111), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1062), .B(new_n1063), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1057), .B1(new_n1058), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n753), .B1(new_n1065), .B2(new_n802), .ZN(new_n1066));
  OR3_X1    g0866(.A1(new_n1054), .A2(new_n1055), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n997), .A2(new_n704), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n742), .B1(new_n995), .B2(new_n996), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1032), .B(new_n1067), .C1(new_n1068), .C2(new_n1069), .ZN(G393));
  NAND3_X1  g0870(.A1(new_n992), .A2(new_n752), .A3(new_n1002), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n801), .B1(new_n554), .B2(new_n212), .C1(new_n253), .C2(new_n803), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n753), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n794), .A2(G77), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1074), .B1(new_n851), .B2(new_n344), .C1(new_n201), .C2(new_n839), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n774), .A2(G68), .B1(new_n789), .B2(G143), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n1076), .A2(KEYINPUT114), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1076), .A2(KEYINPUT114), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n409), .B1(new_n315), .B2(new_n771), .ZN(new_n1079));
  OR4_X1    g0879(.A1(new_n1075), .A2(new_n1077), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(G150), .A2(new_n777), .B1(new_n761), .B2(G159), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT51), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(G311), .A2(new_n761), .B1(new_n777), .B2(G317), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT52), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G294), .A2(new_n778), .B1(new_n782), .B2(G303), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n354), .B1(new_n843), .B2(G107), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n774), .A2(G283), .B1(new_n789), .B2(G322), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n794), .A2(G116), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n1080), .A2(new_n1082), .B1(new_n1084), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1073), .B1(new_n1090), .B2(new_n757), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n956), .B2(new_n812), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1003), .A2(new_n704), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n998), .B1(new_n992), .B2(new_n1002), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1071), .B(new_n1092), .C1(new_n1093), .C2(new_n1094), .ZN(G390));
  NAND2_X1  g0895(.A1(new_n902), .A2(new_n898), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n798), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n810), .B1(new_n833), .B2(new_n344), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n777), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1074), .B1(new_n762), .B2(new_n311), .C1(new_n787), .C2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n319), .B1(new_n773), .B2(new_n315), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n844), .B1(new_n266), .B2(new_n766), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(G97), .A2(new_n778), .B1(new_n782), .B2(G107), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT117), .Z(new_n1105));
  AOI22_X1  g0905(.A1(G128), .A2(new_n777), .B1(new_n761), .B2(G132), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n1019), .B2(new_n839), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n773), .A2(new_n461), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT53), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1109), .B(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(KEYINPUT54), .B(G143), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n851), .A2(new_n1112), .B1(new_n394), .B2(new_n780), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n319), .B1(new_n789), .B2(G125), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n201), .B2(new_n771), .ZN(new_n1115));
  NOR3_X1   g0915(.A1(new_n1111), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1103), .A2(new_n1105), .B1(new_n1108), .B2(new_n1116), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1097), .B(new_n1098), .C1(new_n758), .C2(new_n1117), .ZN(new_n1118));
  AND3_X1   g0918(.A1(new_n937), .A2(G330), .A3(new_n938), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n903), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n914), .A2(new_n1120), .B1(new_n898), .B2(new_n902), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n924), .A2(new_n1120), .A3(new_n934), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT115), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n913), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n910), .A2(new_n912), .A3(KEYINPUT115), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n690), .B(new_n824), .C1(new_n711), .C2(new_n714), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1126), .B1(new_n1127), .B2(new_n907), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1122), .A2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1119), .B1(new_n1121), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1096), .B1(new_n917), .B2(new_n903), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n739), .A2(G330), .A3(new_n824), .A4(new_n913), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1131), .B(new_n1132), .C1(new_n1128), .C2(new_n1122), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1118), .B1(new_n1134), .B2(new_n751), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n745), .B1(new_n930), .B2(new_n718), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1136), .A2(new_n824), .B1(new_n1125), .B2(new_n1124), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1132), .A2(new_n907), .A3(new_n1127), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT116), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n739), .A2(G330), .A3(new_n824), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n916), .A2(new_n1141), .B1(new_n1136), .B2(new_n938), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n908), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1140), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n1141), .A2(new_n916), .ZN(new_n1145));
  OAI211_X1 g0945(.A(KEYINPUT116), .B(new_n908), .C1(new_n1145), .C2(new_n1119), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1139), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n530), .A2(new_n1136), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n922), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1148), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n703), .B1(new_n1152), .B2(new_n1134), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1154), .A2(new_n1133), .A3(new_n1130), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1135), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(G378));
  OAI21_X1  g0957(.A(new_n1151), .B1(new_n1134), .B2(new_n1147), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n745), .B1(new_n939), .B2(new_n940), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n935), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(KEYINPUT121), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT121), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1159), .A2(new_n935), .A3(new_n1162), .ZN(new_n1163));
  XOR2_X1   g0963(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1164));
  XNOR2_X1  g0964(.A(new_n485), .B(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n468), .A2(new_n670), .ZN(new_n1166));
  XOR2_X1   g0966(.A(new_n1166), .B(KEYINPUT120), .Z(new_n1167));
  XOR2_X1   g0967(.A(new_n1165), .B(new_n1167), .Z(new_n1168));
  NAND3_X1  g0968(.A1(new_n1161), .A2(new_n1163), .A3(new_n1168), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n1159), .A2(new_n1162), .A3(new_n935), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1168), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1169), .A2(new_n920), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n920), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1174));
  OAI211_X1 g0974(.A(KEYINPUT57), .B(new_n1158), .C1(new_n1173), .C2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n704), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(KEYINPUT122), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n920), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1162), .B1(new_n1159), .B2(new_n935), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1170), .A2(new_n1179), .A3(new_n1171), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1163), .A2(new_n1168), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1178), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1169), .A2(new_n920), .A3(new_n1172), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(KEYINPUT57), .B1(new_n1184), .B2(new_n1158), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT122), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1175), .A2(new_n1187), .A3(new_n704), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1177), .A2(new_n1186), .A3(new_n1188), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(G97), .A2(new_n782), .B1(new_n778), .B2(new_n348), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1190), .B1(new_n296), .B2(new_n762), .C1(new_n311), .C2(new_n1099), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n771), .A2(new_n203), .ZN(new_n1192));
  XOR2_X1   g0992(.A(new_n1192), .B(KEYINPUT118), .Z(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n265), .A2(new_n701), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1046), .B1(G283), .B2(new_n789), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n204), .B2(new_n780), .ZN(new_n1197));
  NOR4_X1   g0997(.A1(new_n1191), .A2(new_n1194), .A3(new_n1195), .A4(new_n1197), .ZN(new_n1198));
  XOR2_X1   g0998(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(G50), .B1(new_n263), .B2(new_n701), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1198), .A2(new_n1200), .B1(new_n1195), .B2(new_n1201), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n761), .A2(G128), .B1(new_n778), .B2(G137), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n777), .A2(G125), .B1(new_n782), .B2(G132), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n773), .A2(new_n1112), .B1(new_n780), .B2(new_n461), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n263), .B(new_n701), .C1(new_n771), .C2(new_n394), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G124), .B2(new_n789), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT59), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1211), .B1(new_n1207), .B2(new_n1212), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1202), .B1(new_n1209), .B2(new_n1213), .C1(new_n1200), .C2(new_n1198), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n757), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n810), .B1(new_n833), .B2(new_n201), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(new_n1168), .C2(new_n799), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1184), .B2(new_n752), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1189), .A2(new_n1219), .ZN(G375));
  INV_X1    g1020(.A(new_n978), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1152), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1126), .A2(new_n798), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n753), .B1(G68), .B2(new_n834), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n773), .A2(new_n394), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G128), .B2(new_n789), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n778), .A2(G150), .B1(G50), .B2(new_n794), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1227), .A2(new_n409), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n777), .A2(G132), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1230), .B1(new_n839), .B2(new_n1112), .C1(new_n762), .C2(new_n1019), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1193), .B(new_n1229), .C1(new_n1231), .C2(KEYINPUT124), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n1231), .A2(KEYINPUT124), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n773), .A2(new_n554), .B1(new_n766), .B2(new_n785), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT123), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n354), .B(new_n1051), .C1(G77), .C2(new_n843), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n761), .A2(G283), .B1(new_n782), .B2(G116), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n777), .A2(G294), .B1(new_n778), .B2(G107), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n1232), .A2(new_n1233), .B1(new_n1235), .B2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1225), .B1(new_n1240), .B2(new_n757), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1148), .A2(new_n752), .B1(new_n1224), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1223), .A2(new_n1242), .ZN(G381));
  INV_X1    g1043(.A(G390), .ZN(new_n1244));
  NOR4_X1   g1044(.A1(G381), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n1245), .A3(new_n1156), .ZN(new_n1246));
  OR3_X1    g1046(.A1(G375), .A2(new_n1246), .A3(G387), .ZN(G407));
  INV_X1    g1047(.A(new_n1219), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1185), .B1(new_n1176), .B2(KEYINPUT122), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1248), .B1(new_n1249), .B2(new_n1188), .ZN(new_n1250));
  INV_X1    g1050(.A(G343), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(G213), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1250), .A2(new_n1156), .A3(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(G407), .A2(G213), .A3(new_n1254), .ZN(new_n1255));
  XOR2_X1   g1055(.A(new_n1255), .B(KEYINPUT125), .Z(G409));
  INV_X1    g1056(.A(KEYINPUT60), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1222), .B1(new_n1154), .B2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1147), .A2(new_n1150), .A3(KEYINPUT60), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1258), .A2(new_n704), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1242), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1261), .A2(new_n832), .A3(new_n860), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1260), .A2(G384), .A3(new_n1242), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n1156), .B(new_n1248), .C1(new_n1249), .C2(new_n1188), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1184), .A2(new_n1158), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1218), .B1(new_n1268), .B2(new_n1221), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n751), .B1(new_n1184), .B2(KEYINPUT126), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1270), .B1(KEYINPUT126), .B2(new_n1184), .ZN(new_n1271));
  AOI21_X1  g1071(.A(G378), .B1(new_n1269), .B2(new_n1271), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1252), .B(new_n1265), .C1(new_n1266), .C2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(KEYINPUT62), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT61), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1253), .A2(G2897), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1262), .A2(new_n1263), .A3(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1276), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1272), .B1(new_n1250), .B2(G378), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1279), .B1(new_n1280), .B2(new_n1253), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1189), .A2(G378), .A3(new_n1219), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1156), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT62), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1285), .A2(new_n1286), .A3(new_n1252), .A4(new_n1265), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1274), .A2(new_n1275), .A3(new_n1281), .A4(new_n1287), .ZN(new_n1288));
  XOR2_X1   g1088(.A(G393), .B(G396), .Z(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1005), .A2(new_n1030), .A3(G390), .ZN(new_n1291));
  AOI21_X1  g1091(.A(G390), .B1(new_n1005), .B2(new_n1030), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1290), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(G387), .A2(new_n1244), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1005), .A2(new_n1030), .A3(G390), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1294), .A2(new_n1289), .A3(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT127), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1293), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1297), .B1(new_n1293), .B2(new_n1296), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1288), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1293), .A2(new_n1296), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT63), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1302), .B1(new_n1303), .B2(new_n1273), .ZN(new_n1304));
  OR2_X1    g1104(.A1(new_n1273), .A2(new_n1303), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1285), .A2(new_n1252), .ZN(new_n1306));
  AOI21_X1  g1106(.A(KEYINPUT61), .B1(new_n1306), .B2(new_n1279), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1304), .A2(new_n1305), .A3(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1301), .A2(new_n1308), .ZN(G405));
  NOR2_X1   g1109(.A1(new_n1250), .A2(G378), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1310), .A2(new_n1266), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1311), .A2(new_n1264), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1311), .A2(new_n1264), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1313), .A2(new_n1296), .A3(new_n1293), .A4(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1314), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1302), .B1(new_n1316), .B2(new_n1312), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1315), .A2(new_n1317), .ZN(G402));
endmodule


