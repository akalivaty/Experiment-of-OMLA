//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 1 1 0 0 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(new_n187), .B(KEYINPUT70), .Z(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT11), .ZN(new_n190));
  INV_X1    g004(.A(G134), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G137), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(G137), .ZN(new_n193));
  INV_X1    g007(.A(G137), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(KEYINPUT11), .A3(G134), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n192), .A2(new_n193), .A3(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G131), .ZN(new_n197));
  INV_X1    g011(.A(G131), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n192), .A2(new_n195), .A3(new_n198), .A4(new_n193), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(G146), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G143), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n201), .A2(KEYINPUT65), .A3(G146), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n202), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  AND2_X1   g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n204), .A2(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n201), .A2(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(KEYINPUT0), .A2(G128), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n207), .A2(new_n208), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n200), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n205), .A2(new_n206), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT1), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n218), .A2(new_n219), .A3(G128), .A4(new_n209), .ZN(new_n220));
  OAI21_X1  g034(.A(G128), .B1(new_n202), .B2(new_n219), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n211), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n193), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n191), .A2(G137), .ZN(new_n225));
  OAI21_X1  g039(.A(G131), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n223), .A2(new_n199), .A3(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n200), .A2(new_n214), .A3(KEYINPUT66), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n217), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n227), .A2(KEYINPUT30), .A3(new_n215), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT2), .B(G113), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n235));
  XNOR2_X1  g049(.A(G116), .B(G119), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G119), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G116), .ZN(new_n239));
  INV_X1    g053(.A(G116), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G119), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT67), .B1(new_n242), .B2(new_n233), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n237), .A2(new_n243), .B1(new_n242), .B2(new_n233), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n231), .A2(new_n232), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n227), .A2(new_n215), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(new_n245), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(G237), .A2(G953), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G210), .ZN(new_n251));
  INV_X1    g065(.A(G101), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n254));
  XOR2_X1   g068(.A(new_n253), .B(new_n254), .Z(new_n255));
  NAND3_X1  g069(.A1(new_n246), .A2(new_n249), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT31), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n246), .A2(KEYINPUT31), .A3(new_n249), .A4(new_n255), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n255), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT28), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n229), .A2(new_n245), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n248), .B1(new_n263), .B2(KEYINPUT68), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n229), .A2(new_n265), .A3(new_n245), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n262), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n248), .A2(KEYINPUT28), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n261), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n260), .A2(new_n269), .A3(KEYINPUT69), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT69), .B1(new_n260), .B2(new_n269), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n189), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT32), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI211_X1 g088(.A(KEYINPUT32), .B(new_n189), .C1(new_n270), .C2(new_n271), .ZN(new_n275));
  INV_X1    g089(.A(G472), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n263), .A2(KEYINPUT68), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(new_n249), .A3(new_n266), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT28), .ZN(new_n279));
  INV_X1    g093(.A(new_n268), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(new_n280), .A3(new_n255), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT29), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n246), .A2(new_n249), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n261), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n281), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n244), .B1(new_n227), .B2(new_n215), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n286), .B(KEYINPUT71), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n249), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n268), .B1(new_n288), .B2(KEYINPUT28), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n261), .A2(new_n282), .ZN(new_n290));
  AOI21_X1  g104(.A(G902), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n276), .B1(new_n285), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n274), .A2(new_n275), .A3(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G125), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n295), .A2(KEYINPUT16), .A3(G140), .ZN(new_n296));
  OR2_X1    g110(.A1(G125), .A2(G140), .ZN(new_n297));
  NAND2_X1  g111(.A1(G125), .A2(G140), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n296), .B1(new_n299), .B2(KEYINPUT16), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G146), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n238), .A2(G128), .ZN(new_n302));
  INV_X1    g116(.A(G128), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G119), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT24), .B(G110), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT23), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n308), .B1(new_n238), .B2(G128), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n303), .A2(KEYINPUT23), .A3(G119), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n302), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n307), .B1(new_n311), .B2(G110), .ZN(new_n312));
  AND2_X1   g126(.A1(G125), .A2(G140), .ZN(new_n313));
  NOR2_X1   g127(.A1(G125), .A2(G140), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT73), .ZN(new_n315));
  NOR3_X1   g129(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT73), .B1(new_n297), .B2(new_n298), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n204), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n301), .A2(new_n312), .A3(new_n318), .ZN(new_n319));
  XOR2_X1   g133(.A(new_n319), .B(KEYINPUT74), .Z(new_n320));
  XNOR2_X1  g134(.A(new_n300), .B(new_n204), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n311), .A2(G110), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n305), .A2(new_n306), .ZN(new_n323));
  OR3_X1    g137(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT22), .B(G137), .ZN(new_n326));
  INV_X1    g140(.A(G221), .ZN(new_n327));
  INV_X1    g141(.A(G234), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n327), .A2(new_n328), .A3(G953), .ZN(new_n329));
  XOR2_X1   g143(.A(new_n326), .B(new_n329), .Z(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n320), .A2(new_n324), .A3(new_n330), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OR3_X1    g148(.A1(new_n334), .A2(KEYINPUT25), .A3(G902), .ZN(new_n335));
  OAI21_X1  g149(.A(G217), .B1(new_n328), .B2(G902), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n336), .B(KEYINPUT72), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT25), .B1(new_n334), .B2(G902), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n335), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n337), .A2(G902), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n340), .B(KEYINPUT75), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n332), .A2(new_n333), .A3(new_n341), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G475), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n250), .A2(G214), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n201), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n250), .A2(G143), .A3(G214), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n198), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G237), .ZN(new_n349));
  INV_X1    g163(.A(G953), .ZN(new_n350));
  AND4_X1   g164(.A1(G143), .A2(new_n349), .A3(new_n350), .A4(G214), .ZN(new_n351));
  AOI21_X1  g165(.A(G143), .B1(new_n250), .B2(G214), .ZN(new_n352));
  OAI21_X1  g166(.A(G131), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT17), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n348), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  OR2_X1    g169(.A1(new_n353), .A2(new_n354), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n321), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  OAI211_X1 g171(.A(KEYINPUT18), .B(G131), .C1(new_n351), .C2(new_n352), .ZN(new_n358));
  NAND2_X1  g172(.A1(KEYINPUT18), .A2(G131), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n346), .A2(new_n347), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n297), .A2(KEYINPUT73), .A3(new_n298), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n315), .B1(new_n313), .B2(new_n314), .ZN(new_n362));
  AOI21_X1  g176(.A(G146), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n299), .A2(new_n204), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n358), .B(new_n360), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT84), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n365), .A2(new_n366), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n357), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT87), .ZN(new_n370));
  XNOR2_X1  g184(.A(G113), .B(G122), .ZN(new_n371));
  XNOR2_X1  g185(.A(KEYINPUT86), .B(G104), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n371), .B(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n364), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n318), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n376), .A2(KEYINPUT84), .A3(new_n360), .A4(new_n358), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n365), .A2(new_n366), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT87), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(new_n357), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n370), .A2(new_n374), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT88), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT88), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n370), .A2(new_n384), .A3(new_n374), .A4(new_n381), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n379), .A2(new_n373), .A3(new_n357), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n383), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G902), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n344), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(KEYINPUT19), .B1(new_n361), .B2(new_n362), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT19), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n299), .A2(new_n391), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n390), .A2(G146), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n301), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT85), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n348), .A2(new_n353), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n391), .B1(new_n316), .B2(new_n317), .ZN(new_n397));
  INV_X1    g211(.A(new_n392), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n204), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT85), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n400), .A3(new_n301), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n395), .A2(new_n396), .A3(new_n401), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n402), .A2(new_n379), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n386), .B1(new_n403), .B2(new_n373), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT20), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n404), .A2(new_n405), .A3(new_n344), .A4(new_n388), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n373), .B1(new_n402), .B2(new_n379), .ZN(new_n407));
  INV_X1    g221(.A(new_n386), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n344), .B(new_n388), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT20), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(G128), .B(G143), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT13), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n201), .A2(G128), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n413), .B(G134), .C1(KEYINPUT13), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n412), .A2(new_n191), .ZN(new_n416));
  INV_X1    g230(.A(G122), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n417), .A2(KEYINPUT89), .A3(G116), .ZN(new_n418));
  AOI21_X1  g232(.A(KEYINPUT89), .B1(new_n417), .B2(G116), .ZN(new_n419));
  OAI22_X1  g233(.A1(new_n418), .A2(new_n419), .B1(G116), .B2(new_n417), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n420), .A2(G107), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n420), .A2(G107), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n415), .B(new_n416), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT14), .B1(new_n418), .B2(new_n419), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n420), .A2(new_n424), .A3(G107), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n412), .B(new_n191), .ZN(new_n426));
  INV_X1    g240(.A(G107), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n427), .A2(KEYINPUT14), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n425), .B(new_n426), .C1(new_n420), .C2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n423), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(KEYINPUT9), .B(G234), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n432), .A2(G217), .A3(new_n350), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n423), .A2(new_n429), .A3(new_n433), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n388), .ZN(new_n438));
  INV_X1    g252(.A(G478), .ZN(new_n439));
  OR2_X1    g253(.A1(new_n439), .A2(KEYINPUT15), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n438), .B(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n389), .A2(new_n411), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n327), .B1(new_n432), .B2(new_n388), .ZN(new_n444));
  INV_X1    g258(.A(G469), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(new_n388), .ZN(new_n446));
  XNOR2_X1  g260(.A(G110), .B(G140), .ZN(new_n447));
  INV_X1    g261(.A(G227), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(G953), .ZN(new_n449));
  XOR2_X1   g263(.A(new_n447), .B(new_n449), .Z(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G104), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT3), .B1(new_n452), .B2(G107), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT3), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(new_n427), .A3(G104), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n452), .A2(G107), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n453), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G101), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n453), .A2(new_n455), .A3(new_n252), .A4(new_n456), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(KEYINPUT4), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT4), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n457), .A2(new_n461), .A3(G101), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n460), .A2(new_n214), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT77), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n220), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n207), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n221), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n207), .A2(KEYINPUT77), .A3(new_n219), .A4(G128), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n456), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n452), .A2(G107), .ZN(new_n471));
  OAI21_X1  g285(.A(G101), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n472), .A2(new_n459), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT10), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n463), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n200), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n223), .A2(new_n473), .A3(KEYINPUT10), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT78), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT78), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n223), .A2(new_n473), .A3(new_n480), .A4(KEYINPUT10), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n476), .A2(new_n477), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n477), .B1(new_n476), .B2(new_n482), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n451), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n223), .A2(new_n473), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n486), .B1(new_n473), .B2(new_n469), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(KEYINPUT79), .A2(KEYINPUT12), .ZN(new_n489));
  OR2_X1    g303(.A1(KEYINPUT79), .A2(KEYINPUT12), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n488), .A2(new_n200), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n476), .A2(new_n477), .A3(new_n482), .ZN(new_n492));
  OAI211_X1 g306(.A(KEYINPUT79), .B(KEYINPUT12), .C1(new_n487), .C2(new_n477), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n491), .A2(new_n492), .A3(new_n450), .A4(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(G902), .B1(new_n485), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n446), .B1(new_n495), .B2(new_n445), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n450), .B(KEYINPUT76), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n476), .A2(new_n482), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n200), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(new_n492), .A3(new_n450), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n499), .A2(G469), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n444), .B1(new_n496), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(G214), .B1(G237), .B2(G902), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n350), .A2(G952), .ZN(new_n507));
  NAND2_X1  g321(.A1(G234), .A2(G237), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XOR2_X1   g323(.A(KEYINPUT21), .B(G898), .Z(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(G902), .A3(G953), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(G210), .B1(G237), .B2(G902), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  OR2_X1    g329(.A1(new_n214), .A2(new_n295), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n220), .A2(new_n295), .A3(new_n222), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n350), .A2(G224), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n518), .B(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n237), .A2(new_n243), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n236), .A2(KEYINPUT5), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n522), .B(G113), .C1(KEYINPUT5), .C2(new_n239), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n521), .A2(new_n523), .A3(new_n473), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n460), .A2(new_n462), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n524), .B1(new_n525), .B2(new_n244), .ZN(new_n526));
  XNOR2_X1  g340(.A(G110), .B(G122), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(KEYINPUT80), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n528), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n524), .B(new_n530), .C1(new_n525), .C2(new_n244), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n529), .A2(KEYINPUT6), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT6), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n526), .A2(new_n533), .A3(new_n528), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n520), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n388), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n350), .A2(G224), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n518), .B(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n473), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT83), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n522), .A2(KEYINPUT81), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT81), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n236), .A2(new_n543), .A3(KEYINPUT5), .ZN(new_n544));
  OAI21_X1  g358(.A(G113), .B1(new_n239), .B2(KEYINPUT5), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT82), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT82), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n547), .B(G113), .C1(new_n239), .C2(KEYINPUT5), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n542), .A2(new_n544), .A3(new_n546), .A4(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n541), .B1(new_n549), .B2(new_n521), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n541), .A3(new_n521), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n540), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n521), .A2(new_n523), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT8), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n554), .A2(new_n540), .B1(new_n555), .B2(new_n530), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n531), .B1(new_n553), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n530), .A2(new_n555), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n539), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n515), .B1(new_n536), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n539), .ZN(new_n563));
  INV_X1    g377(.A(new_n531), .ZN(new_n564));
  INV_X1    g378(.A(new_n552), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n473), .B1(new_n565), .B2(new_n550), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n564), .B1(new_n566), .B2(new_n556), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n563), .B1(new_n567), .B2(new_n559), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n568), .A2(new_n388), .A3(new_n514), .A4(new_n535), .ZN(new_n569));
  AOI211_X1 g383(.A(new_n506), .B(new_n513), .C1(new_n562), .C2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n443), .A2(new_n504), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n294), .A2(new_n343), .A3(new_n572), .ZN(new_n573));
  XOR2_X1   g387(.A(KEYINPUT90), .B(G101), .Z(new_n574));
  XNOR2_X1  g388(.A(new_n573), .B(new_n574), .ZN(G3));
  NAND2_X1  g389(.A1(new_n260), .A2(new_n269), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT69), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n260), .A2(new_n269), .A3(KEYINPUT69), .ZN(new_n579));
  AOI21_X1  g393(.A(G902), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n343), .B(new_n272), .C1(new_n580), .C2(new_n276), .ZN(new_n581));
  INV_X1    g395(.A(new_n504), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT91), .ZN(new_n584));
  OR2_X1    g398(.A1(new_n569), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n562), .A2(new_n569), .A3(new_n584), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n585), .A2(new_n586), .A3(new_n505), .A4(new_n512), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n382), .A2(KEYINPUT88), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n385), .A2(new_n386), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n388), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n590), .A2(G475), .B1(new_n410), .B2(new_n406), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT33), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n435), .A2(new_n592), .A3(new_n436), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n592), .B1(new_n435), .B2(new_n436), .ZN(new_n595));
  OAI211_X1 g409(.A(G478), .B(new_n388), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT92), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n595), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n593), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n600), .A2(KEYINPUT92), .A3(G478), .A4(new_n388), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n438), .A2(new_n439), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n598), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n587), .A2(new_n591), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n583), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT34), .B(G104), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G6));
  NAND2_X1  g422(.A1(new_n406), .A2(new_n410), .ZN(new_n609));
  OR2_X1    g423(.A1(new_n609), .A2(KEYINPUT93), .ZN(new_n610));
  INV_X1    g424(.A(new_n389), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(KEYINPUT93), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n610), .A2(new_n611), .A3(new_n442), .A4(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(new_n587), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n583), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT35), .B(G107), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G9));
  OAI21_X1  g431(.A(new_n272), .B1(new_n580), .B2(new_n276), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n325), .B(KEYINPUT94), .ZN(new_n620));
  OR3_X1    g434(.A1(new_n620), .A2(KEYINPUT36), .A3(new_n331), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n620), .B1(KEYINPUT36), .B2(new_n331), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n622), .A3(new_n341), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n339), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n619), .A2(new_n572), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT37), .B(G110), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G12));
  AND2_X1   g441(.A1(new_n623), .A2(new_n339), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n585), .A2(new_n586), .A3(new_n505), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n509), .B1(new_n511), .B2(G900), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n613), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n294), .A2(new_n630), .A3(new_n504), .A4(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT95), .B(G128), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G30));
  XOR2_X1   g450(.A(new_n631), .B(KEYINPUT39), .Z(new_n637));
  NOR2_X1   g451(.A1(new_n582), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT40), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n562), .A2(new_n569), .ZN(new_n641));
  XOR2_X1   g455(.A(new_n641), .B(KEYINPUT38), .Z(new_n642));
  NOR2_X1   g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n591), .A2(new_n441), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n628), .A2(new_n644), .A3(new_n505), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT98), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n288), .A2(new_n261), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(G472), .A3(new_n256), .ZN(new_n648));
  NAND2_X1  g462(.A1(G472), .A2(G902), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT96), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n274), .A2(new_n275), .A3(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT97), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n274), .A2(KEYINPUT97), .A3(new_n275), .A4(new_n651), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n643), .A2(new_n646), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G143), .ZN(G45));
  AND2_X1   g471(.A1(new_n385), .A2(new_n386), .ZN(new_n658));
  AOI21_X1  g472(.A(G902), .B1(new_n658), .B2(new_n383), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n609), .B1(new_n659), .B2(new_n344), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n660), .A2(new_n603), .A3(new_n631), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n294), .A2(new_n630), .A3(new_n504), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G146), .ZN(G48));
  INV_X1    g478(.A(new_n494), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n450), .B1(new_n501), .B2(new_n492), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(G469), .B1(new_n667), .B2(G902), .ZN(new_n668));
  INV_X1    g482(.A(new_n444), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n495), .A2(new_n445), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT99), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n668), .A2(KEYINPUT99), .A3(new_n669), .A4(new_n670), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n294), .A2(new_n605), .A3(new_n675), .A4(new_n343), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT41), .B(G113), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G15));
  NAND4_X1  g492(.A1(new_n294), .A2(new_n614), .A3(new_n675), .A4(new_n343), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G116), .ZN(G18));
  NOR4_X1   g494(.A1(new_n671), .A2(new_n660), .A3(new_n442), .A4(new_n513), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n294), .A2(new_n630), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G119), .ZN(G21));
  AOI21_X1  g497(.A(new_n587), .B1(new_n673), .B2(new_n674), .ZN(new_n684));
  OR2_X1    g498(.A1(new_n289), .A2(new_n255), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n188), .B1(new_n685), .B2(new_n260), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n388), .B1(new_n270), .B2(new_n271), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT100), .B(G472), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n684), .A2(new_n343), .A3(new_n644), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G122), .ZN(G24));
  NOR2_X1   g505(.A1(new_n629), .A2(new_n671), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n689), .A2(new_n692), .A3(new_n624), .A4(new_n662), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G125), .ZN(G27));
  INV_X1    g508(.A(KEYINPUT101), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n502), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n502), .A2(new_n695), .ZN(new_n697));
  OAI211_X1 g511(.A(G469), .B(new_n499), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n444), .B1(new_n698), .B2(new_n496), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n662), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n562), .A2(new_n569), .A3(new_n505), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n700), .A2(KEYINPUT42), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n292), .B1(new_n272), .B2(new_n273), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n578), .A2(new_n579), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT102), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n705), .A2(new_n706), .A3(KEYINPUT32), .A4(new_n189), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n275), .A2(KEYINPUT102), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n704), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n709), .A2(KEYINPUT103), .A3(new_n343), .ZN(new_n710));
  AOI21_X1  g524(.A(KEYINPUT103), .B1(new_n709), .B2(new_n343), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n703), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT42), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n294), .A2(new_n343), .A3(new_n699), .A4(new_n702), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n713), .B1(new_n714), .B2(new_n661), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G131), .ZN(G33));
  NAND2_X1  g531(.A1(new_n339), .A2(new_n342), .ZN(new_n718));
  AOI211_X1 g532(.A(new_n718), .B(new_n701), .C1(new_n704), .C2(new_n275), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n719), .A2(KEYINPUT104), .A3(new_n633), .A4(new_n699), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n721));
  INV_X1    g535(.A(new_n633), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n721), .B1(new_n714), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G134), .ZN(G36));
  NAND2_X1  g539(.A1(new_n591), .A2(new_n603), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n728), .A2(KEYINPUT44), .A3(new_n618), .A4(new_n624), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n637), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n728), .A2(new_n618), .A3(new_n624), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT44), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n701), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI211_X1 g549(.A(KEYINPUT45), .B(new_n499), .C1(new_n696), .C2(new_n697), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n499), .A2(new_n502), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n736), .A2(G469), .A3(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n446), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(KEYINPUT46), .A3(new_n741), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n742), .A2(KEYINPUT105), .A3(new_n670), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT105), .B1(new_n742), .B2(new_n670), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT46), .B1(new_n740), .B2(new_n741), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n444), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n731), .A2(new_n732), .A3(new_n735), .A4(new_n747), .ZN(new_n748));
  XOR2_X1   g562(.A(KEYINPUT107), .B(G137), .Z(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(G39));
  XNOR2_X1  g564(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n747), .A2(new_n751), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n294), .A2(new_n343), .A3(new_n661), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n752), .A2(new_n702), .A3(new_n753), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G140), .ZN(G42));
  NAND2_X1  g570(.A1(new_n654), .A2(new_n655), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n671), .A2(new_n509), .A3(new_n701), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n757), .A2(new_n343), .A3(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n660), .A3(new_n603), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n689), .A2(new_n343), .ZN(new_n761));
  INV_X1    g575(.A(new_n509), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n761), .A2(new_n762), .A3(new_n728), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n692), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n760), .A2(new_n507), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT113), .ZN(new_n766));
  INV_X1    g580(.A(new_n671), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n763), .A2(new_n506), .A3(new_n642), .A4(new_n767), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n768), .B(KEYINPUT50), .Z(new_n769));
  AND2_X1   g583(.A1(new_n728), .A2(new_n758), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n624), .A3(new_n689), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n759), .A2(new_n591), .A3(new_n604), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n769), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n668), .A2(new_n670), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n669), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n776), .B1(new_n752), .B2(new_n753), .ZN(new_n777));
  INV_X1    g591(.A(new_n763), .ZN(new_n778));
  OR3_X1    g592(.A1(new_n777), .A2(new_n701), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n773), .A2(new_n774), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n769), .A2(new_n771), .A3(new_n772), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n777), .A2(new_n701), .A3(new_n778), .ZN(new_n782));
  OAI21_X1  g596(.A(KEYINPUT51), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n766), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n676), .A2(new_n679), .A3(new_n682), .A4(new_n690), .ZN(new_n786));
  AOI211_X1 g600(.A(new_n785), .B(new_n786), .C1(new_n712), .C2(new_n715), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n624), .A2(new_n632), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n629), .A2(new_n591), .A3(new_n441), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n652), .A2(new_n699), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n634), .A2(new_n663), .A3(new_n790), .A4(new_n693), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n582), .B1(new_n704), .B2(new_n275), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n794), .B(new_n630), .C1(new_n633), .C2(new_n662), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n795), .A2(KEYINPUT52), .A3(new_n693), .A4(new_n790), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n787), .A2(new_n797), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n442), .A2(new_n632), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n294), .A2(new_n504), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n700), .A2(new_n689), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n624), .A2(new_n702), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  AOI211_X1 g620(.A(new_n718), .B(new_n571), .C1(new_n704), .C2(new_n275), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT110), .B1(new_n660), .B2(new_n603), .ZN(new_n808));
  OAI211_X1 g622(.A(KEYINPUT110), .B(new_n603), .C1(new_n389), .C2(new_n411), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n570), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT111), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT110), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n813), .B1(new_n591), .B2(new_n604), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n809), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT111), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n816), .A3(new_n570), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n807), .B1(new_n818), .B2(new_n583), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n591), .A2(new_n442), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n641), .A2(new_n505), .A3(new_n512), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n619), .A2(new_n343), .A3(new_n504), .A4(new_n822), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n823), .A2(new_n625), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n806), .A2(new_n819), .A3(new_n824), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n720), .A2(new_n723), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n786), .B1(new_n712), .B2(new_n715), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n816), .B1(new_n815), .B2(new_n570), .ZN(new_n829));
  AOI211_X1 g643(.A(KEYINPUT111), .B(new_n821), .C1(new_n814), .C2(new_n809), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n583), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n573), .A3(new_n625), .A4(new_n823), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n804), .B1(new_n801), .B2(new_n802), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n828), .A2(new_n797), .A3(new_n724), .A4(new_n834), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n798), .A2(new_n827), .B1(new_n785), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n835), .A2(new_n785), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT112), .B1(new_n825), .B2(new_n826), .ZN(new_n840));
  INV_X1    g654(.A(new_n832), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n841), .A2(new_n842), .A3(new_n724), .A4(new_n806), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n840), .A2(new_n787), .A3(new_n797), .A4(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n839), .A2(new_n844), .A3(new_n837), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n710), .A2(new_n711), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n770), .ZN(new_n848));
  XOR2_X1   g662(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n849));
  XNOR2_X1  g663(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n784), .A2(new_n838), .A3(new_n845), .A4(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n851), .B1(G952), .B2(G953), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT49), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n642), .B(new_n343), .C1(KEYINPUT109), .C2(new_n853), .ZN(new_n854));
  NOR4_X1   g668(.A1(new_n854), .A2(new_n444), .A3(new_n506), .A4(new_n726), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(KEYINPUT109), .ZN(new_n856));
  XOR2_X1   g670(.A(new_n775), .B(new_n856), .Z(new_n857));
  NAND3_X1  g671(.A1(new_n855), .A2(new_n757), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n852), .A2(new_n858), .ZN(G75));
  AOI21_X1  g673(.A(new_n388), .B1(new_n839), .B2(new_n844), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT56), .B1(new_n860), .B2(G210), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT115), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n532), .A2(new_n534), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n863), .B(new_n520), .Z(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT55), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  OR3_X1    g680(.A1(new_n861), .A2(new_n862), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n350), .A2(G952), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n868), .B1(new_n861), .B2(new_n862), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n866), .B1(new_n861), .B2(new_n862), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n867), .A2(new_n869), .A3(new_n870), .ZN(G51));
  INV_X1    g685(.A(KEYINPUT116), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n446), .B(KEYINPUT57), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n839), .A2(new_n844), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT54), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n874), .B1(new_n876), .B2(new_n845), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n872), .B1(new_n877), .B2(new_n667), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n860), .A2(G469), .A3(new_n739), .A4(new_n736), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n839), .A2(new_n844), .A3(new_n837), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n837), .B1(new_n839), .B2(new_n844), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n873), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n667), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n882), .A2(KEYINPUT116), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n878), .A2(new_n879), .A3(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n868), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n885), .A2(new_n886), .ZN(G54));
  NAND3_X1  g701(.A1(new_n860), .A2(KEYINPUT58), .A3(G475), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(new_n404), .Z(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(new_n868), .ZN(G60));
  OAI21_X1  g704(.A(new_n845), .B1(new_n836), .B2(new_n837), .ZN(new_n891));
  NAND2_X1  g705(.A1(G478), .A2(G902), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT59), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n600), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n600), .B(new_n893), .C1(new_n880), .C2(new_n881), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n895), .A2(KEYINPUT117), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(KEYINPUT117), .ZN(new_n897));
  AOI211_X1 g711(.A(new_n868), .B(new_n894), .C1(new_n896), .C2(new_n897), .ZN(G63));
  AND2_X1   g712(.A1(new_n621), .A2(new_n622), .ZN(new_n899));
  NAND2_X1  g713(.A1(G217), .A2(G902), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT60), .Z(new_n901));
  NAND3_X1  g715(.A1(new_n875), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n875), .A2(new_n901), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n334), .B(KEYINPUT119), .Z(new_n904));
  OAI211_X1 g718(.A(new_n886), .B(new_n902), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n905), .A2(KEYINPUT118), .A3(KEYINPUT61), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT61), .B1(new_n905), .B2(KEYINPUT118), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(G66));
  OR2_X1    g722(.A1(new_n832), .A2(new_n786), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n350), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n510), .A2(G224), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(G953), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n910), .A2(KEYINPUT120), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n913), .B1(KEYINPUT120), .B2(new_n912), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n863), .B1(G898), .B2(new_n350), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT121), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n914), .B(new_n916), .ZN(G69));
  NOR2_X1   g731(.A1(new_n350), .A2(G900), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n918), .B1(new_n448), .B2(G953), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT124), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n231), .A2(new_n232), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n390), .A2(new_n392), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n922), .B(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT123), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n795), .A2(new_n693), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n656), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n656), .A2(new_n926), .A3(new_n929), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n814), .A2(new_n809), .A3(new_n820), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n719), .A2(new_n638), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n755), .A2(new_n748), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n925), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n932), .A2(new_n933), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n748), .A2(new_n936), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n939), .A2(new_n940), .A3(KEYINPUT123), .A4(new_n755), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n924), .B1(new_n942), .B2(new_n350), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n755), .A2(new_n716), .A3(new_n724), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n748), .A2(new_n926), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(KEYINPUT125), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n748), .A2(new_n948), .A3(new_n926), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n945), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n847), .A2(new_n732), .A3(new_n747), .A4(new_n789), .ZN(new_n951));
  AOI21_X1  g765(.A(G953), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n924), .B1(new_n952), .B2(new_n918), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n921), .B1(new_n944), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n924), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n947), .A2(new_n949), .ZN(new_n956));
  INV_X1    g770(.A(new_n945), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n956), .A2(new_n957), .A3(new_n951), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n350), .ZN(new_n959));
  INV_X1    g773(.A(new_n918), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n955), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n961), .A2(new_n943), .A3(new_n920), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n954), .A2(new_n962), .ZN(G72));
  XOR2_X1   g777(.A(new_n649), .B(KEYINPUT63), .Z(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n958), .B2(new_n909), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n283), .B(KEYINPUT126), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n965), .A2(new_n261), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n836), .B1(new_n256), .B2(new_n284), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n868), .B1(new_n968), .B2(new_n964), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n964), .B1(new_n942), .B2(new_n909), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n966), .A2(new_n261), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT127), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n971), .A2(KEYINPUT127), .A3(new_n972), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n970), .B1(new_n975), .B2(new_n976), .ZN(G57));
endmodule


