

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U321 ( .A(n459), .B(n458), .ZN(n568) );
  XNOR2_X1 U322 ( .A(n457), .B(KEYINPUT103), .ZN(n458) );
  NOR2_X1 U323 ( .A1(n432), .A2(n540), .ZN(n569) );
  XOR2_X1 U324 ( .A(KEYINPUT38), .B(n472), .Z(n495) );
  XOR2_X1 U325 ( .A(n443), .B(n367), .Z(n289) );
  XOR2_X1 U326 ( .A(n394), .B(n371), .Z(n290) );
  XNOR2_X1 U327 ( .A(n368), .B(n289), .ZN(n374) );
  XNOR2_X1 U328 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U329 ( .A(n374), .B(n373), .ZN(n375) );
  INV_X1 U330 ( .A(n561), .ZN(n547) );
  XNOR2_X1 U331 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U332 ( .A(n573), .B(KEYINPUT41), .ZN(n561) );
  INV_X1 U333 ( .A(G43GAT), .ZN(n477) );
  INV_X1 U334 ( .A(G29GAT), .ZN(n473) );
  XNOR2_X1 U335 ( .A(n450), .B(G190GAT), .ZN(n451) );
  XNOR2_X1 U336 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U337 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XNOR2_X1 U338 ( .A(n480), .B(n479), .ZN(G1330GAT) );
  XNOR2_X1 U339 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n291) );
  XNOR2_X1 U340 ( .A(n291), .B(KEYINPUT2), .ZN(n417) );
  XOR2_X1 U341 ( .A(G50GAT), .B(G162GAT), .Z(n339) );
  XOR2_X1 U342 ( .A(n417), .B(n339), .Z(n297) );
  XOR2_X1 U343 ( .A(G141GAT), .B(G22GAT), .Z(n344) );
  XNOR2_X1 U344 ( .A(G106GAT), .B(G78GAT), .ZN(n292) );
  XNOR2_X1 U345 ( .A(n292), .B(G148GAT), .ZN(n367) );
  XOR2_X1 U346 ( .A(n367), .B(KEYINPUT96), .Z(n294) );
  NAND2_X1 U347 ( .A1(G228GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U348 ( .A(n294), .B(n293), .ZN(n295) );
  XNOR2_X1 U349 ( .A(n344), .B(n295), .ZN(n296) );
  XNOR2_X1 U350 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U351 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n299) );
  XNOR2_X1 U352 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n298) );
  XNOR2_X1 U353 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U354 ( .A(n301), .B(n300), .Z(n312) );
  XOR2_X1 U355 ( .A(G204GAT), .B(G211GAT), .Z(n303) );
  XNOR2_X1 U356 ( .A(G197GAT), .B(KEYINPUT93), .ZN(n302) );
  XNOR2_X1 U357 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U358 ( .A(KEYINPUT21), .B(KEYINPUT91), .Z(n305) );
  XNOR2_X1 U359 ( .A(G218GAT), .B(KEYINPUT92), .ZN(n304) );
  XNOR2_X1 U360 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U361 ( .A(n307), .B(n306), .Z(n313) );
  XOR2_X1 U362 ( .A(KEYINPUT22), .B(KEYINPUT94), .Z(n309) );
  XNOR2_X1 U363 ( .A(KEYINPUT95), .B(KEYINPUT97), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U365 ( .A(n313), .B(n310), .ZN(n311) );
  XNOR2_X1 U366 ( .A(n312), .B(n311), .ZN(n462) );
  XOR2_X1 U367 ( .A(G92GAT), .B(G64GAT), .Z(n371) );
  XOR2_X1 U368 ( .A(n313), .B(n371), .Z(n315) );
  NAND2_X1 U369 ( .A1(G226GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U370 ( .A(n315), .B(n314), .ZN(n322) );
  XOR2_X1 U371 ( .A(G176GAT), .B(G183GAT), .Z(n317) );
  XNOR2_X1 U372 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n316) );
  XNOR2_X1 U373 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U374 ( .A(KEYINPUT86), .B(KEYINPUT17), .Z(n319) );
  XNOR2_X1 U375 ( .A(G190GAT), .B(KEYINPUT19), .ZN(n318) );
  XNOR2_X1 U376 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U377 ( .A(n321), .B(n320), .Z(n437) );
  XOR2_X1 U378 ( .A(n322), .B(n437), .Z(n324) );
  XNOR2_X1 U379 ( .A(G36GAT), .B(G8GAT), .ZN(n323) );
  XOR2_X1 U380 ( .A(n324), .B(n323), .Z(n515) );
  INV_X1 U381 ( .A(n515), .ZN(n501) );
  XOR2_X1 U382 ( .A(KEYINPUT47), .B(KEYINPUT113), .Z(n400) );
  XOR2_X1 U383 ( .A(G92GAT), .B(G106GAT), .Z(n326) );
  XNOR2_X1 U384 ( .A(G190GAT), .B(G99GAT), .ZN(n325) );
  XNOR2_X1 U385 ( .A(n326), .B(n325), .ZN(n343) );
  XOR2_X1 U386 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n328) );
  NAND2_X1 U387 ( .A1(G232GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U388 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U389 ( .A(n329), .B(KEYINPUT66), .Z(n334) );
  XOR2_X1 U390 ( .A(G29GAT), .B(G36GAT), .Z(n331) );
  XNOR2_X1 U391 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n330) );
  XNOR2_X1 U392 ( .A(n331), .B(n330), .ZN(n348) );
  XNOR2_X1 U393 ( .A(G85GAT), .B(KEYINPUT76), .ZN(n332) );
  XNOR2_X1 U394 ( .A(n332), .B(KEYINPUT77), .ZN(n363) );
  XNOR2_X1 U395 ( .A(n348), .B(n363), .ZN(n333) );
  XNOR2_X1 U396 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U397 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n336) );
  XNOR2_X1 U398 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n335) );
  XNOR2_X1 U399 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U400 ( .A(n338), .B(n337), .Z(n341) );
  XOR2_X1 U401 ( .A(G43GAT), .B(G134GAT), .Z(n442) );
  XNOR2_X1 U402 ( .A(n442), .B(n339), .ZN(n340) );
  XNOR2_X1 U403 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U404 ( .A(n343), .B(n342), .Z(n534) );
  INV_X1 U405 ( .A(n534), .ZN(n555) );
  XOR2_X1 U406 ( .A(G113GAT), .B(G15GAT), .Z(n438) );
  XNOR2_X1 U407 ( .A(n344), .B(n438), .ZN(n347) );
  XOR2_X1 U408 ( .A(G1GAT), .B(KEYINPUT69), .Z(n346) );
  XNOR2_X1 U409 ( .A(G8GAT), .B(KEYINPUT70), .ZN(n345) );
  XNOR2_X1 U410 ( .A(n346), .B(n345), .ZN(n395) );
  XNOR2_X1 U411 ( .A(n347), .B(n395), .ZN(n352) );
  XOR2_X1 U412 ( .A(n348), .B(KEYINPUT29), .Z(n350) );
  NAND2_X1 U413 ( .A1(G229GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U414 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U415 ( .A(n352), .B(n351), .Z(n360) );
  XOR2_X1 U416 ( .A(G197GAT), .B(G50GAT), .Z(n354) );
  XNOR2_X1 U417 ( .A(G169GAT), .B(G43GAT), .ZN(n353) );
  XNOR2_X1 U418 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U419 ( .A(KEYINPUT72), .B(KEYINPUT71), .Z(n356) );
  XNOR2_X1 U420 ( .A(KEYINPUT68), .B(KEYINPUT30), .ZN(n355) );
  XNOR2_X1 U421 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U422 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U423 ( .A(n360), .B(n359), .Z(n543) );
  INV_X1 U424 ( .A(n543), .ZN(n570) );
  XOR2_X1 U425 ( .A(KEYINPUT31), .B(KEYINPUT78), .Z(n362) );
  XNOR2_X1 U426 ( .A(KEYINPUT32), .B(KEYINPUT75), .ZN(n361) );
  XNOR2_X1 U427 ( .A(n362), .B(n361), .ZN(n376) );
  XOR2_X1 U428 ( .A(n363), .B(KEYINPUT33), .Z(n365) );
  NAND2_X1 U429 ( .A1(G230GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U430 ( .A(n365), .B(n364), .ZN(n368) );
  XNOR2_X1 U431 ( .A(G99GAT), .B(G71GAT), .ZN(n366) );
  XNOR2_X1 U432 ( .A(n366), .B(G120GAT), .ZN(n443) );
  XOR2_X1 U433 ( .A(G57GAT), .B(KEYINPUT74), .Z(n370) );
  XNOR2_X1 U434 ( .A(KEYINPUT73), .B(KEYINPUT13), .ZN(n369) );
  XNOR2_X1 U435 ( .A(n370), .B(n369), .ZN(n394) );
  XNOR2_X1 U436 ( .A(G176GAT), .B(G204GAT), .ZN(n372) );
  XNOR2_X1 U437 ( .A(n290), .B(n372), .ZN(n373) );
  XOR2_X1 U438 ( .A(n376), .B(n375), .Z(n573) );
  NOR2_X1 U439 ( .A1(n570), .A2(n561), .ZN(n377) );
  XNOR2_X1 U440 ( .A(n377), .B(KEYINPUT46), .ZN(n378) );
  NOR2_X1 U441 ( .A1(n555), .A2(n378), .ZN(n398) );
  XOR2_X1 U442 ( .A(G155GAT), .B(G78GAT), .Z(n380) );
  XNOR2_X1 U443 ( .A(G22GAT), .B(G211GAT), .ZN(n379) );
  XNOR2_X1 U444 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U445 ( .A(G71GAT), .B(G127GAT), .Z(n382) );
  XNOR2_X1 U446 ( .A(G15GAT), .B(G183GAT), .ZN(n381) );
  XNOR2_X1 U447 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U448 ( .A(n384), .B(n383), .Z(n389) );
  XOR2_X1 U449 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n386) );
  NAND2_X1 U450 ( .A1(G231GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U451 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U452 ( .A(KEYINPUT12), .B(n387), .ZN(n388) );
  XNOR2_X1 U453 ( .A(n389), .B(n388), .ZN(n393) );
  XOR2_X1 U454 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n391) );
  XNOR2_X1 U455 ( .A(G64GAT), .B(KEYINPUT83), .ZN(n390) );
  XNOR2_X1 U456 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U457 ( .A(n393), .B(n392), .Z(n397) );
  XNOR2_X1 U458 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U459 ( .A(n397), .B(n396), .Z(n552) );
  INV_X1 U460 ( .A(n552), .ZN(n577) );
  NAND2_X1 U461 ( .A1(n398), .A2(n577), .ZN(n399) );
  XNOR2_X1 U462 ( .A(n400), .B(n399), .ZN(n407) );
  XOR2_X1 U463 ( .A(n555), .B(KEYINPUT36), .Z(n581) );
  NOR2_X1 U464 ( .A1(n577), .A2(n581), .ZN(n402) );
  XNOR2_X1 U465 ( .A(KEYINPUT45), .B(KEYINPUT65), .ZN(n401) );
  XNOR2_X1 U466 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U467 ( .A(KEYINPUT114), .B(n403), .Z(n404) );
  NAND2_X1 U468 ( .A1(n570), .A2(n404), .ZN(n405) );
  NOR2_X1 U469 ( .A1(n573), .A2(n405), .ZN(n406) );
  NOR2_X1 U470 ( .A1(n407), .A2(n406), .ZN(n408) );
  XNOR2_X1 U471 ( .A(n408), .B(KEYINPUT48), .ZN(n539) );
  NOR2_X1 U472 ( .A1(n501), .A2(n539), .ZN(n410) );
  XNOR2_X1 U473 ( .A(KEYINPUT123), .B(KEYINPUT54), .ZN(n409) );
  XNOR2_X1 U474 ( .A(n410), .B(n409), .ZN(n432) );
  XOR2_X1 U475 ( .A(KEYINPUT0), .B(G127GAT), .Z(n441) );
  XOR2_X1 U476 ( .A(G85GAT), .B(G162GAT), .Z(n412) );
  XNOR2_X1 U477 ( .A(G29GAT), .B(G134GAT), .ZN(n411) );
  XNOR2_X1 U478 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U479 ( .A(n441), .B(n413), .Z(n415) );
  NAND2_X1 U480 ( .A1(G225GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U481 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U482 ( .A(n416), .B(KEYINPUT5), .Z(n419) );
  XNOR2_X1 U483 ( .A(n417), .B(KEYINPUT98), .ZN(n418) );
  XNOR2_X1 U484 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U485 ( .A(G148GAT), .B(G120GAT), .Z(n421) );
  XNOR2_X1 U486 ( .A(G141GAT), .B(G113GAT), .ZN(n420) );
  XNOR2_X1 U487 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U488 ( .A(n423), .B(n422), .Z(n431) );
  XOR2_X1 U489 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n425) );
  XNOR2_X1 U490 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n424) );
  XNOR2_X1 U491 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U492 ( .A(KEYINPUT99), .B(KEYINPUT4), .Z(n427) );
  XNOR2_X1 U493 ( .A(G1GAT), .B(G57GAT), .ZN(n426) );
  XNOR2_X1 U494 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U495 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U496 ( .A(n431), .B(n430), .Z(n498) );
  INV_X1 U497 ( .A(n498), .ZN(n540) );
  NAND2_X1 U498 ( .A1(n462), .A2(n569), .ZN(n433) );
  XNOR2_X1 U499 ( .A(KEYINPUT55), .B(n433), .ZN(n449) );
  XOR2_X1 U500 ( .A(KEYINPUT87), .B(KEYINPUT84), .Z(n435) );
  NAND2_X1 U501 ( .A1(G227GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U502 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U503 ( .A(KEYINPUT20), .B(n436), .ZN(n448) );
  XOR2_X1 U504 ( .A(KEYINPUT64), .B(KEYINPUT85), .Z(n440) );
  XNOR2_X1 U505 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U506 ( .A(n440), .B(n439), .Z(n446) );
  XNOR2_X1 U507 ( .A(n442), .B(n441), .ZN(n444) );
  XOR2_X1 U508 ( .A(n448), .B(n447), .Z(n503) );
  INV_X1 U509 ( .A(n503), .ZN(n525) );
  NAND2_X1 U510 ( .A1(n449), .A2(n525), .ZN(n564) );
  NOR2_X1 U511 ( .A1(n564), .A2(n534), .ZN(n452) );
  XNOR2_X1 U512 ( .A(KEYINPUT58), .B(KEYINPUT125), .ZN(n450) );
  XOR2_X1 U513 ( .A(n515), .B(KEYINPUT102), .Z(n453) );
  XOR2_X1 U514 ( .A(n453), .B(KEYINPUT27), .Z(n460) );
  XNOR2_X1 U515 ( .A(n462), .B(KEYINPUT67), .ZN(n454) );
  XOR2_X1 U516 ( .A(n454), .B(KEYINPUT28), .Z(n506) );
  AND2_X1 U517 ( .A1(n460), .A2(n506), .ZN(n455) );
  NAND2_X1 U518 ( .A1(n540), .A2(n455), .ZN(n523) );
  XOR2_X1 U519 ( .A(KEYINPUT88), .B(n503), .Z(n456) );
  NOR2_X1 U520 ( .A1(n523), .A2(n456), .ZN(n469) );
  NOR2_X1 U521 ( .A1(n525), .A2(n462), .ZN(n459) );
  INV_X1 U522 ( .A(KEYINPUT26), .ZN(n457) );
  NAND2_X1 U523 ( .A1(n568), .A2(n460), .ZN(n538) );
  NAND2_X1 U524 ( .A1(n525), .A2(n515), .ZN(n461) );
  NAND2_X1 U525 ( .A1(n462), .A2(n461), .ZN(n463) );
  XOR2_X1 U526 ( .A(KEYINPUT25), .B(n463), .Z(n464) );
  NAND2_X1 U527 ( .A1(n538), .A2(n464), .ZN(n465) );
  NAND2_X1 U528 ( .A1(n465), .A2(n498), .ZN(n467) );
  INV_X1 U529 ( .A(KEYINPUT104), .ZN(n466) );
  XNOR2_X1 U530 ( .A(n467), .B(n466), .ZN(n468) );
  NOR2_X1 U531 ( .A1(n469), .A2(n468), .ZN(n483) );
  NOR2_X1 U532 ( .A1(n483), .A2(n581), .ZN(n470) );
  NAND2_X1 U533 ( .A1(n470), .A2(n577), .ZN(n471) );
  XNOR2_X1 U534 ( .A(n471), .B(KEYINPUT37), .ZN(n510) );
  NOR2_X1 U535 ( .A1(n570), .A2(n573), .ZN(n484) );
  NAND2_X1 U536 ( .A1(n510), .A2(n484), .ZN(n472) );
  NAND2_X1 U537 ( .A1(n540), .A2(n495), .ZN(n476) );
  XOR2_X1 U538 ( .A(KEYINPUT39), .B(KEYINPUT107), .Z(n474) );
  XNOR2_X1 U539 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U540 ( .A(n476), .B(n475), .ZN(G1328GAT) );
  NAND2_X1 U541 ( .A1(n525), .A2(n495), .ZN(n480) );
  XOR2_X1 U542 ( .A(KEYINPUT108), .B(KEYINPUT40), .Z(n478) );
  NOR2_X1 U543 ( .A1(n577), .A2(n555), .ZN(n481) );
  XOR2_X1 U544 ( .A(KEYINPUT16), .B(n481), .Z(n482) );
  NOR2_X1 U545 ( .A1(n483), .A2(n482), .ZN(n497) );
  NAND2_X1 U546 ( .A1(n484), .A2(n497), .ZN(n491) );
  NOR2_X1 U547 ( .A1(n498), .A2(n491), .ZN(n486) );
  XNOR2_X1 U548 ( .A(KEYINPUT105), .B(KEYINPUT34), .ZN(n485) );
  XNOR2_X1 U549 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U550 ( .A(G1GAT), .B(n487), .ZN(G1324GAT) );
  NOR2_X1 U551 ( .A1(n501), .A2(n491), .ZN(n488) );
  XOR2_X1 U552 ( .A(G8GAT), .B(n488), .Z(G1325GAT) );
  NOR2_X1 U553 ( .A1(n503), .A2(n491), .ZN(n490) );
  XNOR2_X1 U554 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n489) );
  XNOR2_X1 U555 ( .A(n490), .B(n489), .ZN(G1326GAT) );
  NOR2_X1 U556 ( .A1(n506), .A2(n491), .ZN(n492) );
  XOR2_X1 U557 ( .A(KEYINPUT106), .B(n492), .Z(n493) );
  XNOR2_X1 U558 ( .A(G22GAT), .B(n493), .ZN(G1327GAT) );
  NAND2_X1 U559 ( .A1(n495), .A2(n515), .ZN(n494) );
  XNOR2_X1 U560 ( .A(n494), .B(G36GAT), .ZN(G1329GAT) );
  INV_X1 U561 ( .A(n506), .ZN(n519) );
  NAND2_X1 U562 ( .A1(n495), .A2(n519), .ZN(n496) );
  XNOR2_X1 U563 ( .A(n496), .B(G50GAT), .ZN(G1331GAT) );
  NOR2_X1 U564 ( .A1(n543), .A2(n561), .ZN(n511) );
  NAND2_X1 U565 ( .A1(n511), .A2(n497), .ZN(n505) );
  NOR2_X1 U566 ( .A1(n498), .A2(n505), .ZN(n499) );
  XOR2_X1 U567 ( .A(G57GAT), .B(n499), .Z(n500) );
  XNOR2_X1 U568 ( .A(KEYINPUT42), .B(n500), .ZN(G1332GAT) );
  NOR2_X1 U569 ( .A1(n501), .A2(n505), .ZN(n502) );
  XOR2_X1 U570 ( .A(G64GAT), .B(n502), .Z(G1333GAT) );
  NOR2_X1 U571 ( .A1(n503), .A2(n505), .ZN(n504) );
  XOR2_X1 U572 ( .A(G71GAT), .B(n504), .Z(G1334GAT) );
  NOR2_X1 U573 ( .A1(n506), .A2(n505), .ZN(n508) );
  XNOR2_X1 U574 ( .A(KEYINPUT43), .B(KEYINPUT109), .ZN(n507) );
  XNOR2_X1 U575 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U576 ( .A(G78GAT), .B(n509), .Z(G1335GAT) );
  XOR2_X1 U577 ( .A(G85GAT), .B(KEYINPUT111), .Z(n514) );
  NAND2_X1 U578 ( .A1(n511), .A2(n510), .ZN(n512) );
  XOR2_X1 U579 ( .A(KEYINPUT110), .B(n512), .Z(n520) );
  NAND2_X1 U580 ( .A1(n540), .A2(n520), .ZN(n513) );
  XNOR2_X1 U581 ( .A(n514), .B(n513), .ZN(G1336GAT) );
  NAND2_X1 U582 ( .A1(n520), .A2(n515), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n516), .B(KEYINPUT112), .ZN(n517) );
  XNOR2_X1 U584 ( .A(G92GAT), .B(n517), .ZN(G1337GAT) );
  NAND2_X1 U585 ( .A1(n520), .A2(n525), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n518), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U587 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n521), .B(KEYINPUT44), .ZN(n522) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n522), .ZN(G1339GAT) );
  NOR2_X1 U590 ( .A1(n539), .A2(n523), .ZN(n524) );
  NAND2_X1 U591 ( .A1(n525), .A2(n524), .ZN(n533) );
  NOR2_X1 U592 ( .A1(n570), .A2(n533), .ZN(n526) );
  XOR2_X1 U593 ( .A(G113GAT), .B(n526), .Z(G1340GAT) );
  NOR2_X1 U594 ( .A1(n561), .A2(n533), .ZN(n528) );
  XNOR2_X1 U595 ( .A(KEYINPUT115), .B(KEYINPUT49), .ZN(n527) );
  XNOR2_X1 U596 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U597 ( .A(G120GAT), .B(n529), .Z(G1341GAT) );
  NOR2_X1 U598 ( .A1(n577), .A2(n533), .ZN(n531) );
  XNOR2_X1 U599 ( .A(KEYINPUT116), .B(KEYINPUT50), .ZN(n530) );
  XNOR2_X1 U600 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U601 ( .A(G127GAT), .B(n532), .Z(G1342GAT) );
  NOR2_X1 U602 ( .A1(n534), .A2(n533), .ZN(n536) );
  XNOR2_X1 U603 ( .A(KEYINPUT117), .B(KEYINPUT51), .ZN(n535) );
  XNOR2_X1 U604 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U605 ( .A(G134GAT), .B(n537), .Z(G1343GAT) );
  NOR2_X1 U606 ( .A1(n539), .A2(n538), .ZN(n541) );
  NAND2_X1 U607 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U608 ( .A(KEYINPUT118), .B(n542), .Z(n556) );
  NAND2_X1 U609 ( .A1(n556), .A2(n543), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n544), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n546) );
  XNOR2_X1 U612 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n551) );
  XOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT52), .Z(n549) );
  NAND2_X1 U615 ( .A1(n547), .A2(n556), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U617 ( .A(n551), .B(n550), .Z(G1345GAT) );
  NAND2_X1 U618 ( .A1(n556), .A2(n552), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n553), .B(KEYINPUT122), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G155GAT), .B(n554), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n557), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U623 ( .A1(n570), .A2(n564), .ZN(n558) );
  XOR2_X1 U624 ( .A(G169GAT), .B(n558), .Z(G1348GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT124), .B(KEYINPUT56), .Z(n560) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n563) );
  NOR2_X1 U628 ( .A1(n561), .A2(n564), .ZN(n562) );
  XOR2_X1 U629 ( .A(n563), .B(n562), .Z(G1349GAT) );
  NOR2_X1 U630 ( .A1(n577), .A2(n564), .ZN(n565) );
  XOR2_X1 U631 ( .A(G183GAT), .B(n565), .Z(G1350GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT59), .B(KEYINPUT126), .Z(n567) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(n572) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n580) );
  NOR2_X1 U636 ( .A1(n570), .A2(n580), .ZN(n571) );
  XOR2_X1 U637 ( .A(n572), .B(n571), .Z(G1352GAT) );
  XOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT61), .Z(n576) );
  INV_X1 U639 ( .A(n580), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n580), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1354GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U646 ( .A(KEYINPUT62), .B(n582), .Z(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

