//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 1 0 1 0 1 0 1 0 0 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT0), .Z(new_n208));
  AOI22_X1  g0008(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n209));
  INV_X1    g0009(.A(G50), .ZN(new_n210));
  INV_X1    g0010(.A(G226), .ZN(new_n211));
  INV_X1    g0011(.A(G77), .ZN(new_n212));
  INV_X1    g0012(.A(G244), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n214), .B1(G97), .B2(G257), .ZN(new_n215));
  XNOR2_X1  g0015(.A(KEYINPUT65), .B(G68), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G58), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n215), .B(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n205), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(G58), .A2(G68), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT64), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n208), .B(new_n225), .C1(new_n228), .C2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT66), .B(G264), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G270), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(KEYINPUT69), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n227), .A2(G1), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n251), .B1(new_n252), .B2(new_n210), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n226), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n252), .A2(G13), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G20), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(KEYINPUT69), .A3(G50), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n253), .A2(new_n256), .A3(new_n257), .A4(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G13), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n210), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  OR2_X1    g0065(.A1(new_n265), .A2(KEYINPUT70), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(KEYINPUT70), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n227), .B1(new_n229), .B2(new_n210), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G20), .A2(G33), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n268), .B1(G150), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT8), .ZN(new_n271));
  OR3_X1    g0071(.A1(new_n271), .A2(new_n218), .A3(KEYINPUT68), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n271), .B1(new_n218), .B2(KEYINPUT68), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n227), .A2(G33), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n270), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n266), .A2(new_n267), .B1(new_n276), .B2(new_n255), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(KEYINPUT9), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT3), .B(G33), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G222), .ZN(new_n282));
  INV_X1    g0082(.A(G223), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n280), .B(new_n282), .C1(new_n283), .C2(new_n281), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n284), .B(new_n285), .C1(G77), .C2(new_n280), .ZN(new_n286));
  INV_X1    g0086(.A(G33), .ZN(new_n287));
  INV_X1    g0087(.A(G41), .ZN(new_n288));
  OAI211_X1 g0088(.A(G1), .B(G13), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n258), .B1(G41), .B2(G45), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n211), .A2(KEYINPUT67), .ZN(new_n293));
  OR2_X1    g0093(.A1(new_n211), .A2(KEYINPUT67), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G274), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n286), .A2(new_n295), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n277), .A2(KEYINPUT9), .B1(G190), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT10), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n299), .A2(G200), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n279), .A2(new_n301), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n300), .A2(G190), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n276), .A2(new_n255), .ZN(new_n306));
  INV_X1    g0106(.A(new_n267), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n265), .A2(KEYINPUT70), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT9), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n303), .B(new_n305), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT10), .B1(new_n311), .B2(new_n278), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n304), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G179), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n300), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G169), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n299), .A2(new_n316), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n309), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT14), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n292), .A2(G238), .ZN(new_n322));
  NOR2_X1   g0122(.A1(G226), .A2(G1698), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n323), .B1(new_n219), .B2(G1698), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n324), .A2(new_n280), .B1(G33), .B2(G97), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n322), .B(new_n298), .C1(new_n289), .C2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT13), .ZN(new_n327));
  OR2_X1    g0127(.A1(new_n325), .A2(new_n289), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT13), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n328), .A2(new_n329), .A3(new_n298), .A4(new_n322), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n321), .B1(new_n331), .B2(G169), .ZN(new_n332));
  AOI211_X1 g0132(.A(KEYINPUT14), .B(new_n316), .C1(new_n327), .C2(new_n330), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n331), .A2(new_n314), .ZN(new_n334));
  NOR3_X1   g0134(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n216), .A2(new_n227), .ZN(new_n336));
  INV_X1    g0136(.A(new_n269), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n337), .A2(new_n210), .B1(new_n275), .B2(new_n212), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n255), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n339), .B(KEYINPUT11), .ZN(new_n340));
  INV_X1    g0140(.A(G68), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT12), .B1(new_n263), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n257), .A2(KEYINPUT72), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT72), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n252), .A2(new_n344), .A3(G13), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT12), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n216), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n342), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  NOR3_X1   g0149(.A1(new_n346), .A2(new_n255), .A3(new_n252), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT74), .ZN(new_n351));
  AND3_X1   g0151(.A1(new_n350), .A2(new_n351), .A3(G68), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n351), .B1(new_n350), .B2(G68), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n340), .B(new_n349), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n335), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n331), .A2(G200), .ZN(new_n357));
  INV_X1    g0157(.A(G190), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n355), .B(new_n357), .C1(new_n358), .C2(new_n331), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G238), .A2(G1698), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n280), .B(new_n361), .C1(new_n219), .C2(G1698), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n362), .B(new_n285), .C1(G107), .C2(new_n280), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n363), .B(new_n298), .C1(new_n213), .C2(new_n291), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(G200), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT8), .B(G58), .ZN(new_n366));
  OAI22_X1  g0166(.A1(new_n366), .A2(new_n337), .B1(new_n227), .B2(new_n212), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT71), .ZN(new_n368));
  XNOR2_X1  g0168(.A(KEYINPUT15), .B(G87), .ZN(new_n369));
  OR2_X1    g0169(.A1(new_n369), .A2(new_n275), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT71), .ZN(new_n371));
  OAI221_X1 g0171(.A(new_n371), .B1(new_n227), .B2(new_n212), .C1(new_n366), .C2(new_n337), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n368), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n255), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n346), .A2(new_n255), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n375), .A2(G77), .A3(new_n259), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n346), .A2(new_n212), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n374), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT73), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n374), .A2(new_n376), .A3(KEYINPUT73), .A4(new_n377), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n364), .A2(new_n358), .ZN(new_n382));
  AND4_X1   g0182(.A1(new_n365), .A2(new_n380), .A3(new_n381), .A4(new_n382), .ZN(new_n383));
  NOR4_X1   g0183(.A1(new_n320), .A2(new_n356), .A3(new_n360), .A4(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT76), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n341), .A2(KEYINPUT65), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT65), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G68), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n388), .A3(G58), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n227), .B1(new_n389), .B2(new_n230), .ZN(new_n390));
  INV_X1    g0190(.A(G159), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n337), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n385), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT3), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(G33), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n287), .A2(KEYINPUT3), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT7), .B1(new_n397), .B2(new_n227), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT7), .ZN(new_n399));
  AOI211_X1 g0199(.A(new_n399), .B(G20), .C1(new_n395), .C2(new_n396), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n216), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n392), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n229), .B1(new_n216), .B2(G58), .ZN(new_n403));
  OAI211_X1 g0203(.A(KEYINPUT76), .B(new_n402), .C1(new_n403), .C2(new_n227), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n393), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT16), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT75), .B1(new_n287), .B2(KEYINPUT3), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT75), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n409), .A2(new_n394), .A3(G33), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n396), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n412), .A2(new_n399), .A3(new_n227), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n394), .A2(G33), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(new_n408), .B2(new_n410), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT7), .B1(new_n415), .B2(G20), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n413), .A2(G68), .A3(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n417), .A2(KEYINPUT16), .A3(new_n393), .A4(new_n404), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n407), .A2(new_n418), .A3(new_n255), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT77), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT77), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n407), .A2(new_n418), .A3(new_n421), .A4(new_n255), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n283), .A2(new_n281), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n211), .A2(G1698), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n411), .A2(new_n396), .A3(new_n424), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G87), .ZN(new_n427));
  XOR2_X1   g0227(.A(new_n427), .B(KEYINPUT78), .Z(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n297), .B1(new_n429), .B2(new_n285), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n291), .A2(new_n219), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(G190), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n256), .A2(new_n259), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n274), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n435), .B1(new_n274), .B2(new_n263), .ZN(new_n436));
  INV_X1    g0236(.A(G200), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n289), .B1(new_n426), .B2(new_n428), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n438), .A2(new_n297), .A3(new_n431), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n433), .B(new_n436), .C1(new_n437), .C2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT17), .B1(new_n423), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT17), .ZN(new_n443));
  AOI211_X1 g0243(.A(new_n443), .B(new_n440), .C1(new_n420), .C2(new_n422), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n423), .A2(new_n436), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n439), .A2(G179), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n439), .A2(new_n316), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n446), .A2(KEYINPUT18), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT18), .ZN(new_n452));
  INV_X1    g0252(.A(new_n436), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n453), .B1(new_n420), .B2(new_n422), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n452), .B1(new_n454), .B2(new_n449), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n380), .A2(new_n381), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n364), .A2(new_n316), .ZN(new_n458));
  OR2_X1    g0258(.A1(new_n364), .A2(G179), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n384), .A2(new_n445), .A3(new_n456), .A4(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n213), .A2(G1698), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n463), .A2(new_n395), .A3(new_n396), .A4(KEYINPUT4), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT81), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n280), .A2(KEYINPUT81), .A3(KEYINPUT4), .A4(new_n463), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g0268(.A1(G250), .A2(G1698), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n395), .A2(new_n396), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G283), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n409), .B1(new_n394), .B2(G33), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n287), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n396), .B(new_n463), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT4), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n468), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n285), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n258), .B(G45), .C1(new_n288), .C2(KEYINPUT5), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n288), .A2(KEYINPUT5), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT82), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(G274), .B1(new_n482), .B2(KEYINPUT82), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n285), .B1(new_n481), .B2(new_n482), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n486), .B1(G257), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n479), .A2(G190), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n289), .B1(new_n468), .B2(new_n477), .ZN(new_n490));
  OR2_X1    g0290(.A1(new_n484), .A2(new_n485), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n487), .A2(G257), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(G200), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(G97), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n263), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(KEYINPUT79), .B1(new_n287), .B2(G1), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT79), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n499), .A2(new_n258), .A3(G33), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n501), .A2(new_n256), .A3(new_n257), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(new_n496), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(G107), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n399), .B1(new_n280), .B2(G20), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n397), .A2(KEYINPUT7), .A3(new_n227), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n269), .A2(G77), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT6), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n496), .A2(new_n505), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n511), .B1(new_n512), .B2(new_n202), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n505), .A2(KEYINPUT6), .A3(G97), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n227), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR3_X1   g0315(.A1(new_n508), .A2(new_n510), .A3(new_n515), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n497), .B(new_n504), .C1(new_n516), .C2(new_n256), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT80), .ZN(new_n518));
  OAI21_X1  g0318(.A(G107), .B1(new_n398), .B2(new_n400), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n513), .A2(new_n514), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G20), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(new_n509), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n503), .B1(new_n522), .B2(new_n255), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT80), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n524), .A3(new_n497), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n495), .B1(new_n518), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n466), .A2(new_n467), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT4), .B1(new_n415), .B2(new_n463), .ZN(new_n528));
  NOR3_X1   g0328(.A1(new_n527), .A2(new_n528), .A3(new_n472), .ZN(new_n529));
  OAI211_X1 g0329(.A(G179), .B(new_n488), .C1(new_n529), .C2(new_n289), .ZN(new_n530));
  OAI21_X1  g0330(.A(G169), .B1(new_n490), .B2(new_n493), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n530), .A2(new_n531), .B1(new_n523), .B2(new_n497), .ZN(new_n532));
  OAI21_X1  g0332(.A(KEYINPUT83), .B1(new_n526), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n518), .A2(new_n525), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n489), .A2(new_n494), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT83), .ZN(new_n537));
  INV_X1    g0337(.A(new_n532), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n533), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(G45), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n222), .B1(new_n541), .B2(G1), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n258), .A2(new_n296), .A3(G45), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n289), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(G238), .A2(G1698), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(new_n213), .B2(G1698), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n411), .A2(new_n547), .A3(new_n396), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G116), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n545), .B1(new_n550), .B2(new_n285), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n314), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n415), .A2(new_n547), .B1(G33), .B2(G116), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n544), .B1(new_n553), .B2(new_n289), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n316), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n411), .A2(new_n227), .A3(G68), .A4(new_n396), .ZN(new_n556));
  NAND2_X1  g0356(.A1(G33), .A2(G97), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT19), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n227), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(G87), .B2(new_n203), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n558), .B1(new_n557), .B2(G20), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n556), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n255), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n346), .A2(new_n369), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n502), .A2(new_n369), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n552), .B(new_n555), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n554), .A2(G200), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n562), .A2(new_n255), .B1(new_n346), .B2(new_n369), .ZN(new_n569));
  INV_X1    g0369(.A(new_n502), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G87), .ZN(new_n571));
  OAI211_X1 g0371(.A(G190), .B(new_n544), .C1(new_n553), .C2(new_n289), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n568), .A2(new_n569), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT22), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n574), .A2(new_n221), .A3(G20), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n415), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n395), .A2(new_n396), .A3(new_n227), .A4(G87), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n574), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n505), .A2(G20), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT23), .ZN(new_n580));
  XNOR2_X1  g0380(.A(new_n579), .B(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n227), .A2(G33), .A3(G116), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n576), .A2(new_n578), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT24), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n415), .A2(new_n575), .B1(new_n577), .B2(new_n574), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n586), .A2(KEYINPUT24), .A3(new_n581), .A4(new_n582), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n587), .A3(new_n255), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n222), .A2(new_n281), .ZN(new_n589));
  INV_X1    g0389(.A(G257), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G1698), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n411), .A2(new_n396), .A3(new_n589), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(G33), .A2(G294), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n285), .ZN(new_n595));
  INV_X1    g0395(.A(new_n482), .ZN(new_n596));
  OAI211_X1 g0396(.A(G264), .B(new_n289), .C1(new_n596), .C2(new_n480), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n595), .A2(G190), .A3(new_n491), .A4(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n570), .A2(G107), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n257), .A2(G107), .ZN(new_n600));
  XNOR2_X1  g0400(.A(new_n600), .B(KEYINPUT25), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n588), .A2(new_n598), .A3(new_n599), .A4(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n289), .B1(new_n592), .B2(new_n593), .ZN(new_n603));
  INV_X1    g0403(.A(new_n597), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n603), .A2(new_n486), .A3(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n605), .A2(new_n437), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n567), .B(new_n573), .C1(new_n602), .C2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT21), .ZN(new_n608));
  INV_X1    g0408(.A(G116), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n263), .A2(new_n344), .ZN(new_n610));
  NOR3_X1   g0410(.A1(new_n259), .A2(KEYINPUT72), .A3(new_n262), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n609), .B1(new_n498), .B2(new_n500), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n343), .A2(new_n613), .A3(new_n256), .A4(new_n345), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n609), .A2(G20), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n255), .A2(new_n615), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n471), .B(new_n227), .C1(G33), .C2(new_n496), .ZN(new_n617));
  AOI21_X1  g0417(.A(KEYINPUT20), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AND4_X1   g0418(.A1(KEYINPUT20), .A2(new_n617), .A3(new_n255), .A4(new_n615), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n612), .B(new_n614), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G169), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n590), .A2(new_n281), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n281), .A2(G264), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n411), .A2(new_n396), .A3(new_n622), .A4(new_n623), .ZN(new_n624));
  XNOR2_X1  g0424(.A(KEYINPUT84), .B(G303), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n397), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n289), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  OAI211_X1 g0427(.A(G270), .B(new_n289), .C1(new_n596), .C2(new_n480), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n627), .A2(new_n486), .A3(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n608), .B1(new_n621), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n624), .A2(new_n626), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n486), .B1(new_n632), .B2(new_n285), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n628), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n634), .A2(KEYINPUT21), .A3(G169), .A4(new_n620), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n630), .A2(G179), .A3(new_n620), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n631), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n633), .A2(G190), .A3(new_n628), .ZN(new_n638));
  INV_X1    g0438(.A(new_n620), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n638), .B(new_n639), .C1(new_n437), .C2(new_n630), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n637), .A2(KEYINPUT85), .A3(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n640), .A2(new_n631), .A3(new_n635), .A4(new_n636), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT85), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n607), .B1(new_n641), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n588), .A2(new_n599), .A3(new_n601), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n604), .B1(new_n594), .B2(new_n285), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n491), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n316), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n605), .A2(new_n314), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n646), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  AND4_X1   g0451(.A1(new_n462), .A2(new_n540), .A3(new_n645), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n652), .B(KEYINPUT86), .ZN(G372));
  INV_X1    g0453(.A(new_n456), .ZN(new_n654));
  INV_X1    g0454(.A(new_n460), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n356), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n656), .A2(new_n360), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n654), .B1(new_n657), .B2(new_n445), .ZN(new_n658));
  INV_X1    g0458(.A(new_n313), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n319), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n637), .A2(new_n651), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT87), .ZN(new_n663));
  NOR4_X1   g0463(.A1(new_n526), .A2(new_n607), .A3(new_n663), .A4(new_n532), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n665));
  INV_X1    g0465(.A(new_n607), .ZN(new_n666));
  AOI21_X1  g0466(.A(KEYINPUT87), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n662), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT88), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n532), .A2(new_n567), .A3(new_n573), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT26), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n567), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n530), .A2(new_n531), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n518), .A2(new_n674), .A3(new_n525), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n567), .A2(new_n573), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n675), .A2(KEYINPUT26), .A3(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  OAI211_X1 g0478(.A(KEYINPUT88), .B(new_n662), .C1(new_n664), .C2(new_n667), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n670), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n661), .B1(new_n681), .B2(new_n461), .ZN(G369));
  NOR2_X1   g0482(.A1(new_n262), .A2(G20), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n258), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G213), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G343), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n639), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n641), .B2(new_n644), .ZN(new_n692));
  INV_X1    g0492(.A(new_n691), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n637), .A2(new_n693), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT89), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n651), .A2(new_n689), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n646), .A2(new_n689), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n606), .B2(new_n602), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n697), .B1(new_n699), .B2(new_n651), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT90), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n696), .A2(G330), .A3(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n637), .A2(new_n689), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n697), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n705), .ZN(G399));
  INV_X1    g0506(.A(new_n232), .ZN(new_n707));
  INV_X1    g0507(.A(new_n206), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G41), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G1), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n202), .A2(new_n221), .A3(new_n609), .ZN(new_n712));
  OAI22_X1  g0512(.A1(new_n707), .A2(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  OAI21_X1  g0514(.A(KEYINPUT26), .B1(new_n675), .B2(new_n676), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n715), .B(new_n567), .C1(KEYINPUT26), .C2(new_n671), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n665), .A2(new_n662), .A3(new_n666), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT29), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n718), .A2(new_n719), .A3(new_n689), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n680), .A2(new_n690), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n720), .B1(new_n721), .B2(new_n719), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n490), .A2(new_n493), .ZN(new_n723));
  NOR4_X1   g0523(.A1(new_n723), .A2(new_n630), .A3(new_n605), .A4(G179), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n490), .A2(new_n314), .A3(new_n493), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT30), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n554), .A2(new_n603), .A3(new_n604), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n725), .A2(new_n726), .A3(new_n630), .A4(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n633), .A2(new_n647), .A3(new_n628), .A4(new_n551), .ZN(new_n729));
  OAI21_X1  g0529(.A(KEYINPUT30), .B1(new_n530), .B2(new_n729), .ZN(new_n730));
  AOI22_X1  g0530(.A1(new_n554), .A2(new_n724), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT91), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT31), .ZN(new_n733));
  NOR4_X1   g0533(.A1(new_n731), .A2(new_n732), .A3(new_n733), .A4(new_n690), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n728), .A2(new_n730), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n605), .B1(new_n479), .B2(new_n488), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n736), .A2(new_n314), .A3(new_n634), .A4(new_n554), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n733), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(KEYINPUT91), .B1(new_n738), .B2(new_n689), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n734), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n729), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n726), .B1(new_n741), .B2(new_n725), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n530), .A2(new_n729), .A3(KEYINPUT30), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n737), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT92), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n690), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n731), .A2(KEYINPUT92), .ZN(new_n747));
  AOI21_X1  g0547(.A(KEYINPUT31), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(KEYINPUT93), .B1(new_n740), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n744), .A2(KEYINPUT31), .A3(new_n689), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n732), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n738), .A2(KEYINPUT91), .A3(new_n689), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n689), .B1(new_n731), .B2(KEYINPUT92), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n744), .A2(new_n745), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n733), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT93), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n753), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n540), .A2(new_n645), .A3(new_n651), .A4(new_n690), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n749), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n722), .B1(G330), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n714), .B1(new_n761), .B2(G1), .ZN(G364));
  AOI21_X1  g0562(.A(new_n711), .B1(G45), .B2(new_n683), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n696), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G13), .A2(G33), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n764), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n226), .B1(G20), .B2(new_n316), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n437), .A2(G179), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n771), .A2(G20), .A3(G190), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n221), .ZN(new_n773));
  NAND3_X1  g0573(.A1(G20), .A2(G179), .A3(G190), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G200), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n773), .B1(G58), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n771), .A2(G20), .A3(new_n358), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n505), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G179), .A2(G200), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n227), .B1(new_n779), .B2(G190), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n496), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n778), .A2(new_n781), .A3(new_n397), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n227), .A2(new_n314), .A3(G190), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G200), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n774), .A2(new_n437), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n785), .A2(G68), .B1(G50), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n776), .A2(new_n782), .A3(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n779), .A2(G20), .A3(new_n358), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G159), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT95), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT32), .Z(new_n793));
  AND2_X1   g0593(.A1(new_n783), .A2(new_n437), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n794), .A2(KEYINPUT94), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(KEYINPUT94), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n788), .B(new_n793), .C1(G77), .C2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n772), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n797), .A2(G311), .B1(G303), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n786), .B(KEYINPUT96), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G326), .ZN(new_n803));
  INV_X1    g0603(.A(G317), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n784), .B1(KEYINPUT33), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(KEYINPUT33), .B2(new_n804), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n800), .A2(new_n803), .A3(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G283), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n777), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n775), .ZN(new_n810));
  INV_X1    g0610(.A(G322), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n280), .B1(new_n790), .B2(G329), .ZN(new_n813));
  INV_X1    g0613(.A(G294), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n814), .B2(new_n780), .ZN(new_n815));
  NOR4_X1   g0615(.A1(new_n807), .A2(new_n809), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n770), .B1(new_n798), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(G355), .A2(new_n280), .A3(new_n206), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n415), .A2(new_n708), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n707), .B2(G45), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n249), .A2(new_n541), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n818), .B1(G116), .B2(new_n206), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n768), .A2(new_n770), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n769), .A2(new_n817), .A3(new_n824), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT97), .Z(new_n826));
  NOR2_X1   g0626(.A1(new_n696), .A2(G330), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n696), .A2(G330), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n764), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n826), .B1(new_n827), .B2(new_n829), .ZN(G396));
  INV_X1    g0630(.A(KEYINPUT98), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n460), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n457), .A2(KEYINPUT98), .A3(new_n458), .A4(new_n459), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n383), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n680), .A2(new_n690), .A3(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n760), .A2(G330), .ZN(new_n837));
  INV_X1    g0637(.A(new_n834), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n690), .B1(new_n380), .B2(new_n381), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n838), .A2(new_n839), .B1(new_n460), .B2(new_n690), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(new_n680), .B2(new_n690), .ZN(new_n841));
  OR3_X1    g0641(.A1(new_n836), .A2(new_n837), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n837), .B1(new_n836), .B2(new_n841), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n842), .A2(new_n764), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n780), .A2(new_n218), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n785), .A2(G150), .B1(G143), .B2(new_n775), .ZN(new_n846));
  INV_X1    g0646(.A(new_n797), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n846), .B1(new_n847), .B2(new_n391), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(G137), .B2(new_n786), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT34), .Z(new_n850));
  INV_X1    g0650(.A(new_n777), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(G68), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n412), .B1(G132), .B2(new_n790), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n850), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n845), .B(new_n854), .C1(G50), .C2(new_n799), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n851), .A2(G87), .ZN(new_n856));
  INV_X1    g0656(.A(G311), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n397), .B1(new_n789), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(new_n797), .B2(G116), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n799), .A2(G107), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n784), .A2(new_n808), .B1(new_n810), .B2(new_n814), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n781), .B(new_n861), .C1(G303), .C2(new_n786), .ZN(new_n862));
  AND4_X1   g0662(.A1(new_n856), .A2(new_n859), .A3(new_n860), .A4(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n770), .B1(new_n855), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n770), .A2(new_n766), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n212), .ZN(new_n866));
  OR2_X1    g0666(.A1(new_n840), .A2(new_n767), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n864), .A2(new_n763), .A3(new_n866), .A4(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n844), .A2(new_n868), .ZN(G384));
  NAND3_X1  g0669(.A1(new_n832), .A2(new_n690), .A3(new_n833), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n835), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n446), .A2(new_n450), .ZN(new_n873));
  INV_X1    g0673(.A(new_n687), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n446), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n423), .A2(new_n441), .ZN(new_n876));
  XOR2_X1   g0676(.A(KEYINPUT100), .B(KEYINPUT37), .Z(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n873), .A2(new_n875), .A3(new_n876), .A4(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n417), .A2(new_n393), .A3(new_n404), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n406), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(new_n255), .A3(new_n418), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n449), .A2(new_n687), .B1(new_n882), .B2(new_n436), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n440), .B1(new_n420), .B2(new_n422), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT37), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT99), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g0687(.A(KEYINPUT99), .B(KEYINPUT37), .C1(new_n883), .C2(new_n884), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n879), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n882), .A2(new_n436), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n874), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n456), .B2(new_n445), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n872), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT18), .B1(new_n446), .B2(new_n450), .ZN(new_n894));
  NOR3_X1   g0694(.A1(new_n454), .A2(new_n452), .A3(new_n449), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n445), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n891), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n879), .A2(new_n887), .A3(new_n888), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n898), .A2(KEYINPUT38), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n893), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n354), .A2(new_n689), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n359), .B(new_n902), .C1(new_n335), .C2(new_n355), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n332), .A2(new_n333), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n354), .B(new_n689), .C1(new_n904), .C2(new_n334), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n871), .A2(new_n901), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT39), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n898), .A2(KEYINPUT38), .A3(new_n899), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n454), .A2(new_n687), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n896), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n876), .B1(new_n454), .B2(new_n449), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n877), .B1(new_n912), .B2(new_n910), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n879), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT38), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n908), .B1(new_n909), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n356), .A2(new_n690), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n893), .A2(KEYINPUT39), .A3(new_n900), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n916), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n654), .A2(new_n687), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n907), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT101), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n660), .B1(new_n722), .B2(new_n462), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n923), .B(new_n924), .ZN(new_n925));
  AOI211_X1 g0725(.A(new_n383), .B(new_n839), .C1(new_n832), .C2(new_n833), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n460), .A2(new_n690), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n906), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n754), .A2(new_n755), .A3(new_n733), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n929), .A2(new_n748), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n928), .B1(new_n930), .B2(new_n759), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n931), .B(KEYINPUT40), .C1(new_n909), .C2(new_n915), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n746), .A2(KEYINPUT31), .A3(new_n747), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n759), .A2(new_n933), .A3(new_n756), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(new_n840), .A3(new_n906), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(new_n893), .B2(new_n900), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n932), .B(G330), .C1(new_n936), .C2(KEYINPUT40), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n934), .A2(G330), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n461), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT38), .B1(new_n898), .B2(new_n899), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n931), .B1(new_n909), .B2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT40), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(new_n934), .A3(new_n932), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n938), .A2(new_n940), .B1(new_n945), .B2(new_n461), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n925), .B(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n258), .B2(new_n683), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n609), .B1(new_n520), .B2(KEYINPUT35), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n949), .B(new_n228), .C1(KEYINPUT35), .C2(new_n520), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT36), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n232), .A2(G77), .A3(new_n389), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(G50), .B2(new_n341), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(G1), .A3(new_n262), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n948), .A2(new_n951), .A3(new_n954), .ZN(G367));
  AND3_X1   g0755(.A1(new_n696), .A2(G330), .A3(new_n702), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n665), .B1(new_n534), .B2(new_n690), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n675), .A2(new_n690), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n569), .A2(new_n571), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n689), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n567), .A2(new_n962), .A3(new_n573), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n567), .B2(new_n962), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT102), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n960), .B(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n702), .A2(new_n665), .A3(new_n704), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT42), .ZN(new_n970));
  INV_X1    g0770(.A(new_n959), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n538), .B1(new_n971), .B2(new_n651), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n972), .A2(new_n690), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n968), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n967), .B(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n709), .B(KEYINPUT41), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n702), .B1(new_n696), .B2(G330), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n956), .A2(new_n978), .B1(new_n637), .B2(new_n689), .ZN(new_n979));
  INV_X1    g0779(.A(new_n702), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n828), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n981), .A2(new_n703), .A3(new_n704), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  OR3_X1    g0783(.A1(new_n705), .A2(KEYINPUT44), .A3(new_n959), .ZN(new_n984));
  OAI21_X1  g0784(.A(KEYINPUT44), .B1(new_n705), .B2(new_n959), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n705), .A2(new_n959), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT45), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(KEYINPUT45), .B1(new_n705), .B2(new_n959), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n986), .B(new_n703), .C1(new_n989), .C2(new_n990), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n985), .B(new_n984), .C1(new_n989), .C2(new_n990), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n956), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n983), .A2(new_n991), .A3(new_n761), .A4(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n977), .B1(new_n994), .B2(new_n761), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n258), .B1(new_n683), .B2(G45), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n975), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n780), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(G68), .ZN(new_n1000));
  INV_X1    g0800(.A(G150), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n810), .A2(new_n1001), .B1(new_n777), .B2(new_n212), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n797), .A2(G50), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n802), .A2(G143), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n397), .B1(new_n790), .B2(G137), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n799), .A2(G58), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n1002), .B(new_n1007), .C1(G159), .C2(new_n785), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n415), .B1(new_n785), .B2(G294), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n851), .A2(G97), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n799), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n999), .A2(G107), .B1(new_n625), .B2(new_n775), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT46), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n772), .B2(new_n609), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n1015), .A2(KEYINPUT103), .B1(G317), .B2(new_n790), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n847), .B2(new_n808), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1013), .B(new_n1017), .C1(G311), .C2(new_n802), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1015), .A2(KEYINPUT103), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n1000), .A2(new_n1008), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT47), .Z(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n770), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n768), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n964), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n819), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n823), .B1(new_n206), .B2(new_n369), .C1(new_n241), .C2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1022), .A2(new_n763), .A3(new_n1024), .A4(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n998), .A2(new_n1027), .ZN(G387));
  NAND2_X1  g0828(.A1(new_n983), .A2(new_n997), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n366), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n210), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT50), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n341), .A2(new_n212), .ZN(new_n1033));
  NOR4_X1   g0833(.A1(new_n1032), .A2(G45), .A3(new_n1033), .A4(new_n712), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n819), .B1(new_n237), .B2(new_n541), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n280), .A2(new_n712), .A3(new_n206), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n206), .A2(G107), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n823), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n780), .A2(new_n369), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n797), .B2(G68), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n799), .A2(G77), .B1(G50), .B2(new_n775), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n786), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1041), .B(new_n1042), .C1(new_n391), .C2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n415), .B1(new_n274), .B2(new_n784), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1010), .B1(new_n1001), .B2(new_n789), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT104), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n797), .A2(new_n625), .B1(G311), .B2(new_n785), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n804), .B2(new_n810), .C1(new_n801), .C2(new_n811), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT48), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n808), .B2(new_n780), .C1(new_n814), .C2(new_n772), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT49), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n412), .B1(new_n609), .B2(new_n777), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G326), .B2(new_n790), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1048), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n770), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n763), .B(new_n1039), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1058), .A2(KEYINPUT105), .B1(new_n980), .B2(new_n768), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(KEYINPUT105), .B2(new_n1058), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n983), .A2(new_n761), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n709), .B(KEYINPUT106), .Z(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n983), .A2(new_n761), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1029), .B(new_n1060), .C1(new_n1064), .C2(new_n1065), .ZN(G393));
  NAND2_X1  g0866(.A1(new_n991), .A2(new_n993), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1067), .A2(new_n996), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n823), .B1(new_n246), .B2(new_n1025), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G97), .B2(new_n708), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n856), .B1(new_n210), .B2(new_n784), .C1(new_n212), .C2(new_n780), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n412), .B(new_n1072), .C1(new_n216), .C2(new_n799), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n797), .A2(new_n1030), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n790), .A2(G143), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(G150), .A2(new_n786), .B1(new_n775), .B2(G159), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT51), .Z(new_n1077));
  NAND4_X1  g0877(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .A4(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(G311), .A2(new_n775), .B1(new_n786), .B2(G317), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT52), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(G294), .B2(new_n797), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n772), .A2(new_n808), .B1(new_n789), .B2(new_n811), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT107), .Z(new_n1083));
  AOI211_X1 g0883(.A(new_n280), .B(new_n778), .C1(new_n625), .C2(new_n785), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1081), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n780), .A2(new_n609), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1078), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n764), .B(new_n1071), .C1(new_n1087), .C2(new_n770), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT108), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n1023), .B2(new_n959), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n761), .A2(new_n983), .B1(new_n991), .B2(new_n993), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT109), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n1063), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n994), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1069), .B(new_n1090), .C1(new_n1094), .C2(new_n1095), .ZN(G390));
  NAND2_X1  g0896(.A1(new_n916), .A2(new_n919), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n906), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n835), .B2(new_n870), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1097), .B1(new_n1099), .B2(new_n918), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n690), .B(new_n834), .C1(new_n716), .C2(new_n717), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n870), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n906), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1103), .B(new_n917), .C1(new_n909), .C2(new_n915), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(KEYINPUT110), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n913), .A2(new_n879), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n875), .B1(new_n456), .B2(new_n445), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n872), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n918), .B1(new_n1108), .B2(new_n900), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT110), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(new_n1110), .A3(new_n1103), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1105), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n760), .A2(G330), .A3(new_n840), .A4(new_n906), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n1100), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n939), .A2(new_n928), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(new_n1100), .B2(new_n1112), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n934), .A2(G330), .A3(new_n840), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n1098), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(KEYINPUT111), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1102), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT111), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1119), .A2(new_n1123), .A3(new_n1098), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1121), .A2(new_n1113), .A3(new_n1122), .A4(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n758), .A2(new_n759), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n757), .B1(new_n753), .B2(new_n756), .ZN(new_n1127));
  OAI211_X1 g0927(.A(G330), .B(new_n840), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1115), .B1(new_n1128), .B2(new_n1098), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n871), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1125), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n660), .B(new_n940), .C1(new_n722), .C2(new_n462), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1131), .A2(KEYINPUT112), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(KEYINPUT112), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1118), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1100), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n1100), .A2(new_n1112), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1137), .B1(new_n1138), .B2(new_n1116), .ZN(new_n1139));
  AND4_X1   g0939(.A1(new_n1122), .A2(new_n1121), .A3(new_n1113), .A4(new_n1124), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1128), .A2(new_n1098), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1141), .A2(new_n1116), .B1(new_n835), .B2(new_n870), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1132), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT112), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1139), .A2(new_n1145), .A3(new_n1133), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1136), .A2(new_n1146), .A3(new_n1063), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n274), .A2(new_n865), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n767), .B1(new_n916), .B2(new_n919), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n847), .A2(new_n496), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n852), .B1(new_n212), .B2(new_n780), .C1(new_n1043), .C2(new_n808), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n397), .B1(new_n789), .B2(new_n814), .ZN(new_n1152));
  NOR4_X1   g0952(.A1(new_n1150), .A2(new_n1151), .A3(new_n773), .A4(new_n1152), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n1153), .B1(new_n505), .B2(new_n784), .C1(new_n609), .C2(new_n810), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n777), .A2(new_n210), .ZN(new_n1155));
  OR3_X1    g0955(.A1(new_n772), .A2(KEYINPUT53), .A3(new_n1001), .ZN(new_n1156));
  OAI21_X1  g0956(.A(KEYINPUT53), .B1(new_n772), .B2(new_n1001), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n790), .A2(G125), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1156), .A2(new_n280), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1155), .B(new_n1159), .C1(G132), .C2(new_n775), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n786), .A2(G128), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n999), .A2(G159), .ZN(new_n1162));
  XOR2_X1   g0962(.A(KEYINPUT54), .B(G143), .Z(new_n1163));
  AOI22_X1  g0963(.A1(new_n797), .A2(new_n1163), .B1(G137), .B2(new_n785), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .A4(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1057), .B1(new_n1154), .B2(new_n1165), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n1149), .A2(new_n764), .A3(new_n1166), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1118), .A2(new_n997), .B1(new_n1148), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1147), .A2(new_n1168), .ZN(G378));
  INV_X1    g0969(.A(new_n865), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n763), .B1(G50), .B2(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT115), .ZN(new_n1172));
  AOI211_X1 g0972(.A(G41), .B(new_n415), .C1(G283), .C2(new_n790), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1173), .B1(new_n218), .B2(new_n777), .C1(new_n212), .C2(new_n772), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n785), .A2(G97), .B1(G116), .B2(new_n786), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1000), .B(new_n1175), .C1(new_n847), .C2(new_n369), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1174), .B(new_n1176), .C1(G107), .C2(new_n775), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT114), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT58), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n287), .A2(new_n288), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT113), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1181), .B(new_n210), .C1(new_n415), .C2(G41), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n797), .A2(G137), .B1(G150), .B2(new_n999), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n785), .A2(G132), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n775), .A2(G128), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n799), .A2(new_n1163), .B1(G125), .B2(new_n786), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .A4(new_n1186), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT59), .Z(new_n1188));
  NAND2_X1  g0988(.A1(new_n790), .A2(G124), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1181), .B1(G159), .B2(new_n851), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n1179), .A2(new_n1182), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n320), .A2(KEYINPUT55), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT55), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n313), .A2(new_n1194), .A3(new_n319), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1196), .A2(new_n309), .A3(new_n874), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1193), .B(new_n1195), .C1(new_n277), .C2(new_n687), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1199), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1172), .B1(new_n1057), .B2(new_n1192), .C1(new_n1202), .C2(new_n767), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT117), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT118), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1202), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n937), .A2(new_n1206), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n944), .A2(new_n1202), .A3(G330), .A4(new_n932), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1209), .A2(new_n922), .ZN(new_n1210));
  AND2_X1   g1010(.A1(new_n920), .A2(new_n921), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1208), .A2(new_n1207), .B1(new_n1211), .B2(new_n907), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1205), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1209), .A2(new_n922), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1207), .A2(new_n1211), .A3(new_n907), .A4(new_n1208), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1214), .A2(KEYINPUT118), .A3(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1213), .A2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1204), .B1(new_n1217), .B2(new_n997), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT119), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1132), .B(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1136), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(KEYINPUT57), .B1(new_n1222), .B2(new_n1217), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1145), .A2(new_n1133), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1220), .B1(new_n1224), .B2(new_n1118), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1214), .A2(KEYINPUT120), .A3(new_n1215), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT120), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1212), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1226), .A2(KEYINPUT57), .A3(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1063), .B1(new_n1225), .B2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1218), .B1(new_n1223), .B2(new_n1230), .ZN(G375));
  NOR2_X1   g1031(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1224), .A2(new_n977), .A3(new_n1232), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n415), .B1(new_n772), .B2(new_n391), .C1(new_n218), .C2(new_n777), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(new_n797), .B2(G150), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1163), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n1236), .A2(new_n784), .B1(new_n210), .B2(new_n780), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G137), .B2(new_n775), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n790), .A2(G128), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n786), .A2(G132), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1235), .A2(new_n1238), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n777), .A2(new_n212), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1242), .B(new_n1040), .C1(new_n797), .C2(G107), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n775), .A2(G283), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n799), .A2(G97), .B1(new_n790), .B2(G303), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT122), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n280), .B1(new_n786), .B2(G294), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1243), .A2(new_n1244), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n784), .A2(new_n609), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1241), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n764), .B1(new_n1250), .B2(new_n770), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(G68), .B2(new_n1170), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1252), .B(KEYINPUT123), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n906), .A2(new_n767), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1254), .B(KEYINPUT121), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1131), .A2(new_n997), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1233), .A2(new_n1257), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT124), .ZN(G381));
  NOR3_X1   g1059(.A1(G381), .A2(G396), .A3(G393), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1222), .A2(new_n1261), .A3(KEYINPUT57), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1136), .A2(new_n1221), .B1(new_n1213), .B2(new_n1216), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1262), .B(new_n1063), .C1(new_n1263), .C2(KEYINPUT57), .ZN(new_n1264));
  INV_X1    g1064(.A(G378), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1264), .A2(new_n1265), .A3(new_n1218), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1092), .B1(new_n1061), .B2(new_n1067), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n994), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1062), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1068), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1271), .A2(new_n998), .A3(new_n1027), .A4(new_n1090), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1266), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(G384), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1260), .A2(new_n1273), .A3(new_n1274), .ZN(G407));
  INV_X1    g1075(.A(G213), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1276), .A2(G343), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(KEYINPUT125), .B1(new_n1266), .B2(new_n1278), .ZN(new_n1279));
  OR3_X1    g1079(.A1(new_n1266), .A2(KEYINPUT125), .A3(new_n1278), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(G407), .A2(G213), .A3(new_n1279), .A4(new_n1280), .ZN(G409));
  NAND2_X1  g1081(.A1(G375), .A2(G378), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1232), .A2(KEYINPUT60), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1063), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1232), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1145), .A2(KEYINPUT60), .A3(new_n1133), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1284), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1274), .B1(new_n1287), .B2(new_n1257), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1285), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1284), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1291), .A2(G384), .A3(new_n1256), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1288), .A2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1204), .B1(new_n1263), .B2(new_n976), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1226), .A2(new_n997), .A3(new_n1228), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1147), .A2(new_n1168), .A3(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1277), .B1(new_n1294), .B2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1282), .A2(new_n1293), .A3(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT62), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1299), .A2(KEYINPUT126), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1282), .A2(new_n1297), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1277), .A2(G2897), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1288), .A2(new_n1292), .A3(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1303), .B1(new_n1288), .B2(new_n1292), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1302), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT61), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1282), .A2(new_n1297), .A3(new_n1293), .A4(new_n1309), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1301), .A2(new_n1307), .A3(new_n1308), .A4(new_n1310), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(G393), .B(G396), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(G390), .A2(G387), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1312), .B1(new_n1272), .B2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1272), .A2(new_n1313), .A3(new_n1312), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1315), .A2(KEYINPUT127), .A3(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(KEYINPUT127), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1311), .A2(new_n1319), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1282), .A2(new_n1297), .A3(KEYINPUT63), .A4(new_n1293), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1272), .A2(new_n1313), .A3(new_n1312), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1322), .A2(new_n1314), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1321), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1298), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT63), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1326), .B1(new_n1302), .B2(new_n1306), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1324), .B(new_n1308), .C1(new_n1325), .C2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1320), .A2(new_n1328), .ZN(G405));
  NAND2_X1  g1129(.A1(new_n1266), .A2(new_n1282), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1330), .A2(new_n1293), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1288), .A2(new_n1292), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1332), .B1(new_n1266), .B2(new_n1282), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1331), .A2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1319), .A2(new_n1334), .ZN(new_n1335));
  OAI22_X1  g1135(.A1(new_n1317), .A2(new_n1318), .B1(new_n1331), .B2(new_n1333), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(G402));
endmodule


