

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770;

  INV_X2 U383 ( .A(G953), .ZN(n742) );
  XNOR2_X2 U384 ( .A(n538), .B(KEYINPUT103), .ZN(n539) );
  NAND2_X2 U385 ( .A1(n540), .A2(n539), .ZN(n543) );
  AND2_X2 U386 ( .A1(n519), .A2(n518), .ZN(n540) );
  NAND2_X2 U387 ( .A1(n456), .A2(n601), .ZN(n458) );
  XNOR2_X2 U388 ( .A(n495), .B(n396), .ZN(n388) );
  AND2_X1 U389 ( .A1(n372), .A2(n385), .ZN(n371) );
  NAND2_X1 U390 ( .A1(n371), .A2(n387), .ZN(n370) );
  AND2_X1 U391 ( .A1(n382), .A2(n514), .ZN(n377) );
  NAND2_X2 U392 ( .A1(n511), .A2(n509), .ZN(n510) );
  XNOR2_X1 U393 ( .A(n522), .B(KEYINPUT31), .ZN(n720) );
  XNOR2_X1 U394 ( .A(n433), .B(G469), .ZN(n565) );
  XNOR2_X1 U395 ( .A(n754), .B(n383), .ZN(n443) );
  XNOR2_X1 U396 ( .A(KEYINPUT67), .B(G101), .ZN(n383) );
  BUF_X1 U397 ( .A(G116), .Z(n364) );
  BUF_X1 U398 ( .A(n664), .Z(n362) );
  BUF_X1 U399 ( .A(n590), .Z(n363) );
  XNOR2_X2 U400 ( .A(KEYINPUT10), .B(n413), .ZN(n755) );
  INV_X1 U401 ( .A(n732), .ZN(n365) );
  INV_X1 U402 ( .A(n732), .ZN(n726) );
  BUF_X1 U403 ( .A(n388), .Z(n366) );
  XOR2_X2 U404 ( .A(G116), .B(G122), .Z(n489) );
  XNOR2_X2 U405 ( .A(n450), .B(n749), .ZN(n697) );
  XNOR2_X2 U406 ( .A(n458), .B(n457), .ZN(n590) );
  XNOR2_X2 U407 ( .A(n440), .B(n439), .ZN(n749) );
  XNOR2_X1 U408 ( .A(n370), .B(n599), .ZN(n610) );
  NAND2_X1 U409 ( .A1(n515), .A2(n381), .ZN(n376) );
  INV_X1 U410 ( .A(KEYINPUT86), .ZN(n381) );
  NOR2_X1 U411 ( .A1(n588), .A2(n598), .ZN(n372) );
  XNOR2_X1 U412 ( .A(n587), .B(n386), .ZN(n385) );
  OR2_X1 U413 ( .A1(n727), .A2(G902), .ZN(n433) );
  XNOR2_X1 U414 ( .A(n584), .B(n583), .ZN(n607) );
  NAND2_X1 U415 ( .A1(n368), .A2(n506), .ZN(n375) );
  NOR2_X1 U416 ( .A1(n690), .A2(G902), .ZN(n484) );
  INV_X1 U417 ( .A(KEYINPUT46), .ZN(n386) );
  NAND2_X1 U418 ( .A1(n516), .A2(n379), .ZN(n378) );
  NAND2_X1 U419 ( .A1(G234), .A2(G237), .ZN(n460) );
  INV_X1 U420 ( .A(G237), .ZN(n451) );
  XNOR2_X1 U421 ( .A(KEYINPUT85), .B(KEYINPUT48), .ZN(n599) );
  NOR2_X1 U422 ( .A1(G953), .A2(G237), .ZN(n470) );
  XNOR2_X1 U423 ( .A(n388), .B(n443), .ZN(n432) );
  NOR2_X1 U424 ( .A1(n375), .A2(n625), .ZN(n600) );
  XNOR2_X1 U425 ( .A(n478), .B(n374), .ZN(n373) );
  XNOR2_X1 U426 ( .A(n481), .B(n477), .ZN(n374) );
  AND2_X1 U427 ( .A1(n684), .A2(G953), .ZN(n740) );
  XNOR2_X1 U428 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n579) );
  XNOR2_X1 U429 ( .A(n389), .B(n369), .ZN(n585) );
  OR2_X1 U430 ( .A1(n593), .A2(n594), .ZN(n387) );
  XNOR2_X1 U431 ( .A(n375), .B(KEYINPUT112), .ZN(n591) );
  BUF_X1 U432 ( .A(n517), .Z(n695) );
  INV_X1 U433 ( .A(n705), .ZN(n717) );
  OR2_X1 U434 ( .A1(n530), .A2(n529), .ZN(n705) );
  XOR2_X1 U435 ( .A(n452), .B(KEYINPUT92), .Z(n367) );
  AND2_X1 U436 ( .A1(n717), .A2(n589), .ZN(n368) );
  XNOR2_X1 U437 ( .A(KEYINPUT110), .B(KEYINPUT40), .ZN(n369) );
  XNOR2_X1 U438 ( .A(n373), .B(n482), .ZN(n690) );
  NAND2_X1 U439 ( .A1(n377), .A2(n376), .ZN(n380) );
  NAND2_X1 U440 ( .A1(n664), .A2(n663), .ZN(n382) );
  NAND2_X1 U441 ( .A1(n380), .A2(n378), .ZN(n519) );
  INV_X1 U442 ( .A(n382), .ZN(n379) );
  XNOR2_X1 U443 ( .A(n500), .B(n499), .ZN(n517) );
  XNOR2_X2 U444 ( .A(KEYINPUT4), .B(G146), .ZN(n754) );
  INV_X1 U445 ( .A(n456), .ZN(n554) );
  XNOR2_X2 U446 ( .A(n384), .B(n367), .ZN(n456) );
  NAND2_X1 U447 ( .A1(n697), .A2(n670), .ZN(n384) );
  INV_X1 U448 ( .A(n387), .ZN(n723) );
  XNOR2_X1 U449 ( .A(n366), .B(n756), .ZN(n761) );
  INV_X1 U450 ( .A(n585), .ZN(n767) );
  NAND2_X1 U451 ( .A1(n607), .A2(n717), .ZN(n389) );
  XNOR2_X2 U452 ( .A(n441), .B(G134), .ZN(n495) );
  XNOR2_X2 U453 ( .A(n424), .B(n423), .ZN(n624) );
  AND2_X1 U454 ( .A1(n514), .A2(KEYINPUT86), .ZN(n390) );
  OR2_X1 U455 ( .A1(n550), .A2(n462), .ZN(n391) );
  INV_X1 U456 ( .A(n523), .ZN(n466) );
  XNOR2_X1 U457 ( .A(n417), .B(n416), .ZN(n418) );
  INV_X1 U458 ( .A(KEYINPUT101), .ZN(n490) );
  NOR2_X1 U459 ( .A1(n614), .A2(n613), .ZN(n617) );
  NAND2_X1 U460 ( .A1(n463), .A2(n391), .ZN(n465) );
  XNOR2_X1 U461 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U462 ( .A(n493), .B(n492), .ZN(n494) );
  INV_X1 U463 ( .A(KEYINPUT39), .ZN(n583) );
  XNOR2_X1 U464 ( .A(n727), .B(n728), .ZN(n729) );
  XNOR2_X1 U465 ( .A(n730), .B(n729), .ZN(n731) );
  XNOR2_X1 U466 ( .A(n580), .B(n579), .ZN(n769) );
  XNOR2_X2 U467 ( .A(KEYINPUT64), .B(G143), .ZN(n393) );
  INV_X1 U468 ( .A(G128), .ZN(n392) );
  XNOR2_X2 U469 ( .A(n393), .B(n392), .ZN(n441) );
  XNOR2_X1 U470 ( .A(G137), .B(G131), .ZN(n395) );
  INV_X1 U471 ( .A(KEYINPUT70), .ZN(n394) );
  XNOR2_X1 U472 ( .A(n395), .B(n394), .ZN(n396) );
  NAND2_X1 U473 ( .A1(n470), .A2(G210), .ZN(n397) );
  XNOR2_X1 U474 ( .A(n397), .B(KEYINPUT5), .ZN(n399) );
  XNOR2_X1 U475 ( .A(n364), .B(KEYINPUT73), .ZN(n398) );
  XNOR2_X1 U476 ( .A(n399), .B(n398), .ZN(n402) );
  XNOR2_X1 U477 ( .A(G119), .B(G113), .ZN(n401) );
  XNOR2_X2 U478 ( .A(KEYINPUT90), .B(KEYINPUT3), .ZN(n400) );
  XNOR2_X1 U479 ( .A(n401), .B(n400), .ZN(n437) );
  XNOR2_X1 U480 ( .A(n402), .B(n437), .ZN(n403) );
  XNOR2_X1 U481 ( .A(n432), .B(n403), .ZN(n681) );
  OR2_X2 U482 ( .A1(n681), .A2(G902), .ZN(n404) );
  INV_X1 U483 ( .A(G472), .ZN(n679) );
  XNOR2_X2 U484 ( .A(n404), .B(n679), .ZN(n620) );
  XNOR2_X1 U485 ( .A(n620), .B(KEYINPUT6), .ZN(n506) );
  XNOR2_X1 U486 ( .A(G119), .B(G137), .ZN(n405) );
  XOR2_X1 U487 ( .A(n405), .B(KEYINPUT23), .Z(n409) );
  XOR2_X1 U488 ( .A(KEYINPUT77), .B(KEYINPUT24), .Z(n407) );
  XNOR2_X1 U489 ( .A(G110), .B(G128), .ZN(n406) );
  XNOR2_X1 U490 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U491 ( .A(n409), .B(n408), .ZN(n412) );
  NAND2_X1 U492 ( .A1(G234), .A2(n742), .ZN(n410) );
  XOR2_X1 U493 ( .A(KEYINPUT8), .B(n410), .Z(n486) );
  NAND2_X1 U494 ( .A1(G221), .A2(n486), .ZN(n411) );
  XNOR2_X1 U495 ( .A(n412), .B(n411), .ZN(n414) );
  XOR2_X1 U496 ( .A(G125), .B(G140), .Z(n413) );
  XOR2_X1 U497 ( .A(G146), .B(n755), .Z(n482) );
  XOR2_X1 U498 ( .A(n414), .B(n482), .Z(n737) );
  OR2_X1 U499 ( .A1(G902), .A2(n737), .ZN(n419) );
  XNOR2_X1 U500 ( .A(KEYINPUT15), .B(G902), .ZN(n670) );
  NAND2_X1 U501 ( .A1(G234), .A2(n670), .ZN(n415) );
  XNOR2_X1 U502 ( .A(KEYINPUT20), .B(n415), .ZN(n420) );
  AND2_X1 U503 ( .A1(n420), .A2(G217), .ZN(n417) );
  XNOR2_X1 U504 ( .A(KEYINPUT25), .B(KEYINPUT76), .ZN(n416) );
  XNOR2_X2 U505 ( .A(n419), .B(n418), .ZN(n507) );
  NAND2_X1 U506 ( .A1(n420), .A2(G221), .ZN(n422) );
  INV_X1 U507 ( .A(KEYINPUT21), .ZN(n421) );
  XNOR2_X1 U508 ( .A(n422), .B(n421), .ZN(n618) );
  NAND2_X1 U509 ( .A1(n507), .A2(n618), .ZN(n424) );
  INV_X1 U510 ( .A(KEYINPUT68), .ZN(n423) );
  AND2_X1 U511 ( .A1(n506), .A2(n624), .ZN(n434) );
  XNOR2_X1 U512 ( .A(G110), .B(G107), .ZN(n425) );
  XNOR2_X1 U513 ( .A(n425), .B(KEYINPUT89), .ZN(n427) );
  XNOR2_X1 U514 ( .A(G104), .B(KEYINPUT74), .ZN(n426) );
  XNOR2_X1 U515 ( .A(n427), .B(n426), .ZN(n439) );
  XOR2_X1 U516 ( .A(G140), .B(KEYINPUT78), .Z(n429) );
  NAND2_X1 U517 ( .A1(G227), .A2(n742), .ZN(n428) );
  XNOR2_X1 U518 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U519 ( .A(n439), .B(n430), .ZN(n431) );
  XNOR2_X1 U520 ( .A(n432), .B(n431), .ZN(n727) );
  XNOR2_X2 U521 ( .A(n565), .B(KEYINPUT1), .ZN(n625) );
  NAND2_X1 U522 ( .A1(n434), .A2(n625), .ZN(n436) );
  XNOR2_X1 U523 ( .A(KEYINPUT71), .B(KEYINPUT33), .ZN(n435) );
  XNOR2_X2 U524 ( .A(n436), .B(n435), .ZN(n636) );
  INV_X1 U525 ( .A(n636), .ZN(n467) );
  XNOR2_X1 U526 ( .A(n489), .B(KEYINPUT16), .ZN(n438) );
  XNOR2_X1 U527 ( .A(n438), .B(n437), .ZN(n440) );
  INV_X1 U528 ( .A(n441), .ZN(n442) );
  XNOR2_X1 U529 ( .A(n443), .B(n442), .ZN(n449) );
  XOR2_X1 U530 ( .A(KEYINPUT18), .B(KEYINPUT91), .Z(n445) );
  NAND2_X1 U531 ( .A1(G224), .A2(n742), .ZN(n444) );
  XNOR2_X1 U532 ( .A(n445), .B(n444), .ZN(n447) );
  XNOR2_X1 U533 ( .A(KEYINPUT17), .B(G125), .ZN(n446) );
  XNOR2_X1 U534 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U535 ( .A(n449), .B(n448), .ZN(n450) );
  INV_X1 U536 ( .A(G902), .ZN(n496) );
  NAND2_X1 U537 ( .A1(n496), .A2(n451), .ZN(n453) );
  NAND2_X1 U538 ( .A1(n453), .A2(G210), .ZN(n452) );
  NAND2_X1 U539 ( .A1(n453), .A2(G214), .ZN(n455) );
  INV_X1 U540 ( .A(KEYINPUT93), .ZN(n454) );
  XNOR2_X1 U541 ( .A(n455), .B(n454), .ZN(n601) );
  INV_X1 U542 ( .A(n601), .ZN(n637) );
  INV_X1 U543 ( .A(KEYINPUT87), .ZN(n457) );
  XNOR2_X1 U544 ( .A(KEYINPUT75), .B(KEYINPUT19), .ZN(n459) );
  XNOR2_X1 U545 ( .A(n590), .B(n459), .ZN(n567) );
  INV_X1 U546 ( .A(n567), .ZN(n463) );
  XNOR2_X1 U547 ( .A(n460), .B(KEYINPUT14), .ZN(n461) );
  AND2_X1 U548 ( .A1(n461), .A2(G952), .ZN(n651) );
  AND2_X1 U549 ( .A1(n651), .A2(n742), .ZN(n550) );
  OR2_X1 U550 ( .A1(n742), .A2(G898), .ZN(n750) );
  NAND2_X1 U551 ( .A1(G902), .A2(n461), .ZN(n546) );
  NOR2_X1 U552 ( .A1(n750), .A2(n546), .ZN(n462) );
  XNOR2_X1 U553 ( .A(KEYINPUT66), .B(KEYINPUT0), .ZN(n464) );
  XNOR2_X2 U554 ( .A(n465), .B(n464), .ZN(n523) );
  NAND2_X1 U555 ( .A1(n467), .A2(n466), .ZN(n469) );
  INV_X1 U556 ( .A(KEYINPUT34), .ZN(n468) );
  XNOR2_X1 U557 ( .A(n469), .B(n468), .ZN(n498) );
  XOR2_X1 U558 ( .A(G122), .B(G143), .Z(n472) );
  NAND2_X1 U559 ( .A1(n470), .A2(G214), .ZN(n471) );
  XNOR2_X1 U560 ( .A(n472), .B(n471), .ZN(n476) );
  XOR2_X1 U561 ( .A(KEYINPUT12), .B(KEYINPUT99), .Z(n474) );
  XNOR2_X1 U562 ( .A(G131), .B(KEYINPUT98), .ZN(n473) );
  XNOR2_X1 U563 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U564 ( .A(n476), .B(n475), .Z(n478) );
  XNOR2_X1 U565 ( .A(G113), .B(G104), .ZN(n477) );
  XOR2_X1 U566 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n480) );
  XNOR2_X1 U567 ( .A(KEYINPUT11), .B(KEYINPUT95), .ZN(n479) );
  XNOR2_X1 U568 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U569 ( .A(KEYINPUT13), .B(KEYINPUT100), .ZN(n483) );
  XNOR2_X1 U570 ( .A(n484), .B(n483), .ZN(n485) );
  INV_X1 U571 ( .A(G475), .ZN(n688) );
  XNOR2_X1 U572 ( .A(n485), .B(n688), .ZN(n530) );
  XOR2_X1 U573 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n488) );
  NAND2_X1 U574 ( .A1(G217), .A2(n486), .ZN(n487) );
  XNOR2_X1 U575 ( .A(n488), .B(n487), .ZN(n493) );
  XNOR2_X1 U576 ( .A(n489), .B(G107), .ZN(n491) );
  XNOR2_X1 U577 ( .A(n495), .B(n494), .ZN(n734) );
  NAND2_X1 U578 ( .A1(n734), .A2(n496), .ZN(n497) );
  INV_X1 U579 ( .A(G478), .ZN(n733) );
  XNOR2_X1 U580 ( .A(n497), .B(n733), .ZN(n528) );
  NOR2_X1 U581 ( .A1(n530), .A2(n528), .ZN(n555) );
  NAND2_X1 U582 ( .A1(n498), .A2(n555), .ZN(n500) );
  XNOR2_X1 U583 ( .A(KEYINPUT84), .B(KEYINPUT35), .ZN(n499) );
  AND2_X1 U584 ( .A1(n528), .A2(n530), .ZN(n639) );
  NAND2_X1 U585 ( .A1(n639), .A2(n618), .ZN(n501) );
  OR2_X2 U586 ( .A1(n523), .A2(n501), .ZN(n504) );
  INV_X1 U587 ( .A(KEYINPUT72), .ZN(n502) );
  XNOR2_X1 U588 ( .A(n502), .B(KEYINPUT22), .ZN(n503) );
  XNOR2_X2 U589 ( .A(n504), .B(n503), .ZN(n511) );
  INV_X1 U590 ( .A(KEYINPUT88), .ZN(n505) );
  XNOR2_X1 U591 ( .A(n625), .B(n505), .ZN(n594) );
  INV_X1 U592 ( .A(n507), .ZN(n558) );
  OR2_X1 U593 ( .A1(n506), .A2(n507), .ZN(n508) );
  NOR2_X1 U594 ( .A1(n594), .A2(n508), .ZN(n509) );
  XNOR2_X2 U595 ( .A(n510), .B(KEYINPUT32), .ZN(n664) );
  XNOR2_X1 U596 ( .A(n620), .B(KEYINPUT104), .ZN(n544) );
  BUF_X1 U597 ( .A(n544), .Z(n562) );
  NAND2_X1 U598 ( .A1(n562), .A2(n558), .ZN(n512) );
  NOR2_X1 U599 ( .A1(n512), .A2(n625), .ZN(n513) );
  NAND2_X1 U600 ( .A1(n511), .A2(n513), .ZN(n663) );
  INV_X1 U601 ( .A(KEYINPUT44), .ZN(n514) );
  INV_X1 U602 ( .A(n517), .ZN(n515) );
  NAND2_X1 U603 ( .A1(n515), .A2(n390), .ZN(n516) );
  NAND2_X1 U604 ( .A1(n695), .A2(KEYINPUT44), .ZN(n518) );
  INV_X1 U605 ( .A(n624), .ZN(n520) );
  NOR2_X1 U606 ( .A1(n620), .A2(n520), .ZN(n521) );
  NAND2_X1 U607 ( .A1(n625), .A2(n521), .ZN(n630) );
  OR2_X1 U608 ( .A1(n523), .A2(n630), .ZN(n522) );
  INV_X1 U609 ( .A(n720), .ZN(n527) );
  NAND2_X1 U610 ( .A1(n565), .A2(n624), .ZN(n551) );
  OR2_X1 U611 ( .A1(n523), .A2(n551), .ZN(n525) );
  INV_X1 U612 ( .A(KEYINPUT94), .ZN(n524) );
  XNOR2_X1 U613 ( .A(n525), .B(n524), .ZN(n526) );
  NAND2_X1 U614 ( .A1(n526), .A2(n620), .ZN(n708) );
  NAND2_X1 U615 ( .A1(n527), .A2(n708), .ZN(n532) );
  INV_X1 U616 ( .A(n528), .ZN(n529) );
  AND2_X1 U617 ( .A1(n530), .A2(n529), .ZN(n719) );
  INV_X1 U618 ( .A(n719), .ZN(n709) );
  AND2_X1 U619 ( .A1(n709), .A2(n705), .ZN(n641) );
  XNOR2_X1 U620 ( .A(n641), .B(KEYINPUT80), .ZN(n569) );
  INV_X1 U621 ( .A(n569), .ZN(n531) );
  NAND2_X1 U622 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U623 ( .A(n533), .B(KEYINPUT102), .ZN(n537) );
  OR2_X1 U624 ( .A1(n506), .A2(n558), .ZN(n534) );
  NOR2_X1 U625 ( .A1(n625), .A2(n534), .ZN(n535) );
  AND2_X1 U626 ( .A1(n511), .A2(n535), .ZN(n703) );
  INV_X1 U627 ( .A(n703), .ZN(n536) );
  NAND2_X1 U628 ( .A1(n537), .A2(n536), .ZN(n538) );
  INV_X1 U629 ( .A(KEYINPUT83), .ZN(n541) );
  XNOR2_X1 U630 ( .A(n541), .B(KEYINPUT45), .ZN(n542) );
  XNOR2_X2 U631 ( .A(n543), .B(n542), .ZN(n741) );
  NOR2_X1 U632 ( .A1(n544), .A2(n637), .ZN(n545) );
  XNOR2_X1 U633 ( .A(n545), .B(KEYINPUT30), .ZN(n553) );
  NOR2_X1 U634 ( .A1(G900), .A2(n546), .ZN(n547) );
  NAND2_X1 U635 ( .A1(G953), .A2(n547), .ZN(n548) );
  XNOR2_X1 U636 ( .A(KEYINPUT105), .B(n548), .ZN(n549) );
  NOR2_X1 U637 ( .A1(n550), .A2(n549), .ZN(n560) );
  NOR2_X1 U638 ( .A1(n560), .A2(n551), .ZN(n552) );
  NAND2_X1 U639 ( .A1(n553), .A2(n552), .ZN(n582) );
  INV_X1 U640 ( .A(n554), .ZN(n604) );
  NAND2_X1 U641 ( .A1(n555), .A2(n604), .ZN(n556) );
  NOR2_X1 U642 ( .A1(n582), .A2(n556), .ZN(n557) );
  XNOR2_X1 U643 ( .A(n557), .B(KEYINPUT108), .ZN(n768) );
  NAND2_X1 U644 ( .A1(n558), .A2(n618), .ZN(n559) );
  NOR2_X1 U645 ( .A1(n560), .A2(n559), .ZN(n589) );
  INV_X1 U646 ( .A(n589), .ZN(n561) );
  NOR2_X1 U647 ( .A1(n562), .A2(n561), .ZN(n564) );
  XOR2_X1 U648 ( .A(KEYINPUT28), .B(KEYINPUT109), .Z(n563) );
  XNOR2_X1 U649 ( .A(n564), .B(n563), .ZN(n566) );
  NAND2_X1 U650 ( .A1(n566), .A2(n565), .ZN(n576) );
  NOR2_X1 U651 ( .A1(n576), .A2(n567), .ZN(n715) );
  INV_X1 U652 ( .A(n715), .ZN(n572) );
  INV_X1 U653 ( .A(KEYINPUT47), .ZN(n597) );
  XNOR2_X1 U654 ( .A(n597), .B(KEYINPUT69), .ZN(n568) );
  NOR2_X1 U655 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U656 ( .A1(n570), .A2(KEYINPUT79), .ZN(n571) );
  NOR2_X1 U657 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U658 ( .A1(n768), .A2(n573), .ZN(n575) );
  NAND2_X1 U659 ( .A1(KEYINPUT79), .A2(n597), .ZN(n574) );
  NAND2_X1 U660 ( .A1(n575), .A2(n574), .ZN(n588) );
  INV_X1 U661 ( .A(n576), .ZN(n578) );
  XNOR2_X1 U662 ( .A(n554), .B(KEYINPUT38), .ZN(n581) );
  AND2_X1 U663 ( .A1(n581), .A2(n601), .ZN(n643) );
  NAND2_X1 U664 ( .A1(n639), .A2(n643), .ZN(n577) );
  XNOR2_X1 U665 ( .A(n577), .B(KEYINPUT41), .ZN(n653) );
  NAND2_X1 U666 ( .A1(n578), .A2(n653), .ZN(n580) );
  INV_X1 U667 ( .A(n769), .ZN(n586) );
  INV_X1 U668 ( .A(n581), .ZN(n638) );
  NOR2_X2 U669 ( .A1(n582), .A2(n638), .ZN(n584) );
  NAND2_X1 U670 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U671 ( .A1(n591), .A2(n363), .ZN(n592) );
  XOR2_X1 U672 ( .A(KEYINPUT36), .B(n592), .Z(n593) );
  NOR2_X1 U673 ( .A1(n715), .A2(KEYINPUT79), .ZN(n595) );
  NOR2_X1 U674 ( .A1(n641), .A2(n595), .ZN(n596) );
  NOR2_X1 U675 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U676 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n603) );
  NAND2_X1 U677 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U678 ( .A(n603), .B(n602), .Z(n605) );
  NOR2_X1 U679 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U680 ( .A(n606), .B(KEYINPUT107), .ZN(n766) );
  AND2_X1 U681 ( .A1(n607), .A2(n719), .ZN(n725) );
  INV_X1 U682 ( .A(n725), .ZN(n608) );
  AND2_X1 U683 ( .A1(n766), .A2(n608), .ZN(n609) );
  AND2_X2 U684 ( .A1(n610), .A2(n609), .ZN(n615) );
  NAND2_X1 U685 ( .A1(n741), .A2(n615), .ZN(n675) );
  INV_X1 U686 ( .A(KEYINPUT2), .ZN(n665) );
  NOR2_X1 U687 ( .A1(n665), .A2(KEYINPUT81), .ZN(n611) );
  AND2_X1 U688 ( .A1(n675), .A2(n611), .ZN(n614) );
  XNOR2_X1 U689 ( .A(n741), .B(KEYINPUT81), .ZN(n612) );
  NOR2_X1 U690 ( .A1(n612), .A2(KEYINPUT2), .ZN(n613) );
  INV_X1 U691 ( .A(n615), .ZN(n760) );
  NOR2_X1 U692 ( .A1(n615), .A2(KEYINPUT2), .ZN(n616) );
  NOR2_X1 U693 ( .A1(n617), .A2(n616), .ZN(n658) );
  NOR2_X1 U694 ( .A1(n507), .A2(n618), .ZN(n619) );
  XOR2_X1 U695 ( .A(KEYINPUT49), .B(n619), .Z(n622) );
  INV_X1 U696 ( .A(n620), .ZN(n621) );
  NOR2_X1 U697 ( .A1(n622), .A2(n621), .ZN(n623) );
  XOR2_X1 U698 ( .A(n623), .B(KEYINPUT118), .Z(n628) );
  NOR2_X1 U699 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U700 ( .A(KEYINPUT50), .B(n626), .ZN(n627) );
  NOR2_X1 U701 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U702 ( .A(KEYINPUT119), .B(n629), .Z(n632) );
  INV_X1 U703 ( .A(n630), .ZN(n631) );
  NOR2_X1 U704 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U705 ( .A(KEYINPUT51), .B(n633), .ZN(n634) );
  NAND2_X1 U706 ( .A1(n634), .A2(n653), .ZN(n635) );
  XNOR2_X1 U707 ( .A(n635), .B(KEYINPUT120), .ZN(n648) );
  INV_X1 U708 ( .A(n636), .ZN(n654) );
  NAND2_X1 U709 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U710 ( .A1(n640), .A2(n639), .ZN(n645) );
  INV_X1 U711 ( .A(n641), .ZN(n642) );
  NAND2_X1 U712 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U713 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U714 ( .A1(n654), .A2(n646), .ZN(n647) );
  NAND2_X1 U715 ( .A1(n648), .A2(n647), .ZN(n650) );
  XNOR2_X1 U716 ( .A(KEYINPUT52), .B(KEYINPUT121), .ZN(n649) );
  XOR2_X1 U717 ( .A(n650), .B(n649), .Z(n652) );
  NAND2_X1 U718 ( .A1(n652), .A2(n651), .ZN(n656) );
  NAND2_X1 U719 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U720 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X2 U721 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U722 ( .A(n659), .B(KEYINPUT122), .ZN(n660) );
  NAND2_X1 U723 ( .A1(n660), .A2(n742), .ZN(n662) );
  INV_X1 U724 ( .A(KEYINPUT53), .ZN(n661) );
  XNOR2_X1 U725 ( .A(n662), .B(n661), .ZN(G75) );
  XNOR2_X1 U726 ( .A(n663), .B(G110), .ZN(G12) );
  XNOR2_X1 U727 ( .A(n362), .B(G119), .ZN(G21) );
  NAND2_X1 U728 ( .A1(KEYINPUT2), .A2(KEYINPUT82), .ZN(n667) );
  NOR2_X1 U729 ( .A1(n665), .A2(KEYINPUT82), .ZN(n666) );
  NAND2_X1 U730 ( .A1(n670), .A2(n666), .ZN(n669) );
  AND2_X1 U731 ( .A1(n667), .A2(n669), .ZN(n668) );
  NAND2_X1 U732 ( .A1(n675), .A2(n668), .ZN(n674) );
  INV_X1 U733 ( .A(n669), .ZN(n672) );
  INV_X1 U734 ( .A(n670), .ZN(n671) );
  OR2_X1 U735 ( .A1(n672), .A2(n671), .ZN(n673) );
  AND2_X2 U736 ( .A1(n674), .A2(n673), .ZN(n678) );
  INV_X1 U737 ( .A(n675), .ZN(n676) );
  NAND2_X1 U738 ( .A1(n676), .A2(KEYINPUT2), .ZN(n677) );
  NAND2_X2 U739 ( .A1(n678), .A2(n677), .ZN(n732) );
  NOR2_X1 U740 ( .A1(n732), .A2(n679), .ZN(n683) );
  XNOR2_X1 U741 ( .A(KEYINPUT113), .B(KEYINPUT62), .ZN(n680) );
  XNOR2_X1 U742 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U743 ( .A(n683), .B(n682), .ZN(n685) );
  INV_X1 U744 ( .A(G952), .ZN(n684) );
  NOR2_X1 U745 ( .A1(n685), .A2(n740), .ZN(n687) );
  XOR2_X1 U746 ( .A(KEYINPUT114), .B(KEYINPUT63), .Z(n686) );
  XNOR2_X1 U747 ( .A(n687), .B(n686), .ZN(G57) );
  NOR2_X1 U748 ( .A1(n732), .A2(n688), .ZN(n692) );
  XOR2_X1 U749 ( .A(KEYINPUT65), .B(KEYINPUT59), .Z(n689) );
  XNOR2_X1 U750 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U751 ( .A(n692), .B(n691), .ZN(n693) );
  NOR2_X1 U752 ( .A1(n693), .A2(n740), .ZN(n694) );
  XNOR2_X1 U753 ( .A(n694), .B(KEYINPUT60), .ZN(G60) );
  INV_X1 U754 ( .A(G122), .ZN(n696) );
  XNOR2_X1 U755 ( .A(n696), .B(n695), .ZN(G24) );
  NAND2_X1 U756 ( .A1(n365), .A2(G210), .ZN(n700) );
  XNOR2_X1 U757 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n698) );
  XNOR2_X1 U758 ( .A(n697), .B(n698), .ZN(n699) );
  XNOR2_X1 U759 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X2 U760 ( .A1(n701), .A2(n740), .ZN(n702) );
  XNOR2_X1 U761 ( .A(n702), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U762 ( .A(G101), .B(n703), .ZN(n704) );
  XNOR2_X1 U763 ( .A(n704), .B(KEYINPUT115), .ZN(G3) );
  NOR2_X1 U764 ( .A1(n708), .A2(n705), .ZN(n706) );
  XOR2_X1 U765 ( .A(KEYINPUT116), .B(n706), .Z(n707) );
  XNOR2_X1 U766 ( .A(G104), .B(n707), .ZN(G6) );
  XOR2_X1 U767 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n711) );
  NOR2_X1 U768 ( .A1(n708), .A2(n709), .ZN(n710) );
  XOR2_X1 U769 ( .A(n711), .B(n710), .Z(n712) );
  XNOR2_X1 U770 ( .A(G107), .B(n712), .ZN(G9) );
  XOR2_X1 U771 ( .A(G128), .B(KEYINPUT29), .Z(n714) );
  NAND2_X1 U772 ( .A1(n715), .A2(n719), .ZN(n713) );
  XNOR2_X1 U773 ( .A(n714), .B(n713), .ZN(G30) );
  NAND2_X1 U774 ( .A1(n715), .A2(n717), .ZN(n716) );
  XNOR2_X1 U775 ( .A(n716), .B(G146), .ZN(G48) );
  NAND2_X1 U776 ( .A1(n720), .A2(n717), .ZN(n718) );
  XNOR2_X1 U777 ( .A(n718), .B(G113), .ZN(G15) );
  XOR2_X1 U778 ( .A(n364), .B(KEYINPUT117), .Z(n722) );
  NAND2_X1 U779 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U780 ( .A(n722), .B(n721), .ZN(G18) );
  XNOR2_X1 U781 ( .A(n723), .B(G125), .ZN(n724) );
  XNOR2_X1 U782 ( .A(n724), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U783 ( .A(G134), .B(n725), .Z(G36) );
  NAND2_X1 U784 ( .A1(n726), .A2(G469), .ZN(n730) );
  XOR2_X1 U785 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n728) );
  NOR2_X1 U786 ( .A1(n740), .A2(n731), .ZN(G54) );
  NOR2_X1 U787 ( .A1(n732), .A2(n733), .ZN(n735) );
  XNOR2_X1 U788 ( .A(n735), .B(n734), .ZN(n736) );
  NOR2_X1 U789 ( .A1(n740), .A2(n736), .ZN(G63) );
  NAND2_X1 U790 ( .A1(n726), .A2(G217), .ZN(n738) );
  XNOR2_X1 U791 ( .A(n738), .B(n737), .ZN(n739) );
  NOR2_X1 U792 ( .A1(n740), .A2(n739), .ZN(G66) );
  NAND2_X1 U793 ( .A1(n741), .A2(n742), .ZN(n743) );
  XOR2_X1 U794 ( .A(KEYINPUT123), .B(n743), .Z(n747) );
  NAND2_X1 U795 ( .A1(G953), .A2(G224), .ZN(n744) );
  XNOR2_X1 U796 ( .A(KEYINPUT61), .B(n744), .ZN(n745) );
  NAND2_X1 U797 ( .A1(n745), .A2(G898), .ZN(n746) );
  NAND2_X1 U798 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U799 ( .A(n748), .B(KEYINPUT124), .ZN(n753) );
  XOR2_X1 U800 ( .A(n749), .B(G101), .Z(n751) );
  NAND2_X1 U801 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U802 ( .A(n753), .B(n752), .Z(G69) );
  XNOR2_X1 U803 ( .A(n755), .B(n754), .ZN(n756) );
  XNOR2_X1 U804 ( .A(n761), .B(KEYINPUT126), .ZN(n757) );
  XNOR2_X1 U805 ( .A(G227), .B(n757), .ZN(n758) );
  NAND2_X1 U806 ( .A1(n758), .A2(G900), .ZN(n759) );
  NAND2_X1 U807 ( .A1(n759), .A2(G953), .ZN(n765) );
  XOR2_X1 U808 ( .A(n761), .B(n760), .Z(n762) );
  NOR2_X1 U809 ( .A1(G953), .A2(n762), .ZN(n763) );
  XNOR2_X1 U810 ( .A(KEYINPUT125), .B(n763), .ZN(n764) );
  NAND2_X1 U811 ( .A1(n765), .A2(n764), .ZN(G72) );
  XNOR2_X1 U812 ( .A(G140), .B(n766), .ZN(G42) );
  XOR2_X1 U813 ( .A(n767), .B(G131), .Z(G33) );
  XOR2_X1 U814 ( .A(G143), .B(n768), .Z(G45) );
  XNOR2_X1 U815 ( .A(G137), .B(KEYINPUT127), .ZN(n770) );
  XNOR2_X1 U816 ( .A(n770), .B(n769), .ZN(G39) );
endmodule

