//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 0 1 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1296, new_n1297,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1369, new_n1370, new_n1371;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(new_n204), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT64), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n209), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT65), .Z(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  INV_X1    g0019(.A(G97), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT69), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G68), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT67), .B(G238), .ZN(new_n226));
  INV_X1    g0026(.A(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT68), .B(G77), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT66), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n231), .B1(new_n222), .B2(new_n223), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n206), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  OR2_X1    g0033(.A1(new_n233), .A2(KEYINPUT1), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n233), .A2(KEYINPUT1), .ZN(new_n235));
  AND3_X1   g0035(.A1(new_n216), .A2(new_n234), .A3(new_n235), .ZN(G361));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT70), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n240), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT71), .ZN(new_n247));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  XNOR2_X1  g0053(.A(KEYINPUT3), .B(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G232), .ZN(new_n257));
  INV_X1    g0057(.A(G107), .ZN(new_n258));
  OAI22_X1  g0058(.A1(new_n256), .A2(new_n257), .B1(new_n258), .B2(new_n254), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n254), .A2(G1698), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT73), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n260), .B(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n226), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n259), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(G1), .A2(G13), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G41), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  AND2_X1   g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  OAI21_X1  g0069(.A(G274), .B1(new_n269), .B2(new_n210), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT72), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G274), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n274), .B1(new_n265), .B2(new_n266), .ZN(new_n275));
  INV_X1    g0075(.A(new_n272), .ZN(new_n276));
  AOI21_X1  g0076(.A(KEYINPUT72), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n267), .A2(new_n272), .ZN(new_n278));
  OAI22_X1  g0078(.A1(new_n273), .A2(new_n277), .B1(new_n227), .B2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n268), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G190), .ZN(new_n281));
  INV_X1    g0081(.A(new_n228), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G20), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G20), .A2(G33), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n204), .A2(G33), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT15), .B(G87), .ZN(new_n288));
  OAI221_X1 g0088(.A(new_n283), .B1(new_n285), .B2(new_n286), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n210), .ZN(new_n291));
  INV_X1    g0091(.A(G13), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(G1), .ZN(new_n293));
  AOI21_X1  g0093(.A(KEYINPUT75), .B1(new_n293), .B2(G20), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n203), .A2(G13), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT75), .ZN(new_n296));
  NOR3_X1   g0096(.A1(new_n295), .A2(new_n296), .A3(new_n204), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n289), .A2(new_n291), .B1(new_n228), .B2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n291), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n300), .B(G77), .C1(G1), .C2(new_n204), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G200), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n281), .B(new_n303), .C1(new_n304), .C2(new_n280), .ZN(new_n305));
  INV_X1    g0105(.A(G179), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n280), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(new_n268), .B2(new_n279), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(new_n302), .A3(new_n309), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n271), .B1(new_n270), .B2(new_n272), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n275), .A2(KEYINPUT72), .A3(new_n276), .ZN(new_n313));
  INV_X1    g0113(.A(new_n278), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n312), .A2(new_n313), .B1(new_n314), .B2(G226), .ZN(new_n315));
  INV_X1    g0115(.A(G222), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n256), .A2(new_n316), .B1(new_n228), .B2(new_n254), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n317), .B1(new_n262), .B2(G223), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n315), .B1(new_n318), .B2(new_n267), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n319), .A2(G179), .ZN(new_n320));
  NOR2_X1   g0120(.A1(G50), .A2(G58), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n204), .B1(new_n321), .B2(new_n225), .ZN(new_n322));
  INV_X1    g0122(.A(G150), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n286), .A2(new_n287), .B1(new_n323), .B2(new_n285), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT74), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n322), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(new_n325), .B2(new_n324), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n291), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n295), .A2(new_n204), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(new_n291), .ZN(new_n330));
  INV_X1    g0130(.A(G50), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(new_n203), .B2(G20), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n330), .A2(new_n332), .B1(new_n331), .B2(new_n329), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n319), .A2(new_n308), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n320), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G190), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n319), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n338), .B(KEYINPUT76), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n334), .A2(KEYINPUT9), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n334), .A2(KEYINPUT9), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n340), .A2(new_n341), .B1(G200), .B2(new_n319), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT10), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n339), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n343), .B1(new_n339), .B2(new_n342), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n311), .B(new_n336), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n298), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT12), .B1(new_n347), .B2(G68), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n225), .A2(G20), .ZN(new_n349));
  OR3_X1    g0149(.A1(new_n349), .A2(new_n295), .A3(KEYINPUT12), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n225), .B1(new_n203), .B2(G20), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n348), .A2(new_n350), .B1(new_n300), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G77), .ZN(new_n353));
  OAI221_X1 g0153(.A(new_n349), .B1(new_n287), .B2(new_n353), .C1(new_n285), .C2(new_n331), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n291), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT11), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n354), .A2(KEYINPUT11), .A3(new_n291), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(KEYINPUT80), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT80), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n357), .A2(new_n361), .A3(new_n358), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n352), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT79), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n273), .B2(new_n277), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n312), .A2(KEYINPUT79), .A3(new_n313), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n314), .A2(G238), .ZN(new_n367));
  AND3_X1   g0167(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT13), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G33), .A2(G97), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT77), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT77), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n372), .A2(G33), .A3(G97), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G33), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT3), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT3), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G33), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n376), .A2(new_n378), .A3(G226), .A4(new_n255), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n376), .A2(new_n378), .A3(G232), .A4(G1698), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n374), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT78), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT78), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n374), .A2(new_n379), .A3(new_n380), .A4(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n269), .A2(new_n210), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n368), .A2(new_n369), .A3(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n267), .B1(new_n382), .B2(new_n384), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT13), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT14), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(new_n393), .A3(G169), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n388), .A2(G179), .A3(new_n391), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n393), .B1(new_n392), .B2(G169), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n363), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n392), .A2(G200), .ZN(new_n399));
  INV_X1    g0199(.A(new_n363), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n388), .A2(G190), .A3(new_n391), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n273), .A2(new_n277), .B1(new_n257), .B2(new_n278), .ZN(new_n404));
  MUX2_X1   g0204(.A(G223), .B(G226), .S(G1698), .Z(new_n405));
  INV_X1    g0205(.A(KEYINPUT81), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n377), .ZN(new_n407));
  NAND2_X1  g0207(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n407), .A2(G33), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n405), .A2(new_n409), .A3(new_n376), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G87), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n267), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NOR3_X1   g0212(.A1(new_n404), .A2(new_n412), .A3(G179), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n410), .A2(new_n411), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n386), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n312), .A2(new_n313), .B1(new_n314), .B2(G232), .ZN(new_n416));
  AOI21_X1  g0216(.A(G169), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT82), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n308), .B1(new_n404), .B2(new_n412), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n415), .A2(new_n416), .A3(new_n306), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT82), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n286), .B1(new_n203), .B2(G20), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n424), .A2(new_n330), .B1(new_n329), .B2(new_n286), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n291), .ZN(new_n427));
  INV_X1    g0227(.A(G58), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(new_n225), .ZN(new_n429));
  NOR2_X1   g0229(.A1(G58), .A2(G68), .ZN(new_n430));
  OAI21_X1  g0230(.A(G20), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n284), .A2(G159), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(G20), .B1(new_n409), .B2(new_n376), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT7), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n225), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n376), .ZN(new_n437));
  AND2_X1   g0237(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n438));
  NOR2_X1   g0238(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n437), .B1(new_n440), .B2(G33), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT7), .B1(new_n441), .B2(G20), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n433), .B1(new_n436), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n427), .B1(new_n443), .B2(KEYINPUT16), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT16), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n435), .A2(G20), .ZN(new_n446));
  AOI21_X1  g0246(.A(G33), .B1(new_n407), .B2(new_n408), .ZN(new_n447));
  INV_X1    g0247(.A(new_n378), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n435), .B1(new_n254), .B2(G20), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n225), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n445), .B1(new_n451), .B2(new_n433), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n426), .B1(new_n444), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT18), .B1(new_n423), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n433), .ZN(new_n455));
  NOR3_X1   g0255(.A1(new_n438), .A2(new_n439), .A3(new_n375), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n435), .B(new_n204), .C1(new_n456), .C2(new_n437), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G68), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n434), .A2(new_n435), .ZN(new_n459));
  OAI211_X1 g0259(.A(KEYINPUT16), .B(new_n455), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n460), .A2(new_n452), .A3(new_n291), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n425), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT18), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n462), .A2(new_n463), .A3(new_n418), .A4(new_n422), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n304), .B1(new_n404), .B2(new_n412), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n415), .A2(new_n416), .A3(new_n337), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n461), .A2(new_n467), .A3(new_n425), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT17), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n461), .A2(new_n467), .A3(KEYINPUT17), .A4(new_n425), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n454), .A2(new_n464), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n346), .A2(new_n403), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n329), .A2(new_n258), .ZN(new_n474));
  XOR2_X1   g0274(.A(new_n474), .B(KEYINPUT25), .Z(new_n475));
  OAI21_X1  g0275(.A(new_n330), .B1(G1), .B2(new_n375), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n475), .B1(new_n258), .B2(new_n476), .ZN(new_n477));
  AND2_X1   g0277(.A1(KEYINPUT22), .A2(G87), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n409), .A2(new_n204), .A3(new_n376), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G116), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(G20), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT23), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(new_n204), .B2(G107), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n258), .A2(KEYINPUT23), .A3(G20), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n376), .A2(new_n378), .ZN(new_n486));
  NOR3_X1   g0286(.A1(new_n486), .A2(G20), .A3(new_n218), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n479), .B(new_n485), .C1(new_n487), .C2(KEYINPUT22), .ZN(new_n488));
  XNOR2_X1  g0288(.A(new_n488), .B(KEYINPUT24), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n477), .B1(new_n489), .B2(new_n291), .ZN(new_n490));
  INV_X1    g0290(.A(G41), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n203), .B(G45), .C1(new_n491), .C2(KEYINPUT5), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT5), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n493), .A2(G41), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n267), .B(G264), .C1(new_n492), .C2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n492), .A2(KEYINPUT84), .ZN(new_n496));
  INV_X1    g0296(.A(G45), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(G1), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT84), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n493), .A2(G41), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n494), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n496), .A2(new_n501), .A3(new_n275), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G294), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(G250), .A2(G1698), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n506), .B1(new_n221), .B2(G1698), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n505), .B1(new_n441), .B2(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n495), .B(new_n503), .C1(new_n508), .C2(new_n267), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT92), .ZN(new_n510));
  INV_X1    g0310(.A(new_n495), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n507), .A2(new_n409), .A3(new_n376), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n504), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n511), .B1(new_n513), .B2(new_n386), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT92), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n514), .A2(new_n515), .A3(new_n503), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n510), .A2(G169), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n514), .A2(G179), .A3(new_n503), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT93), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n490), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n517), .A2(KEYINPUT93), .A3(new_n518), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n515), .B1(new_n514), .B2(new_n503), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n267), .B1(new_n512), .B2(new_n504), .ZN(new_n524));
  INV_X1    g0324(.A(new_n503), .ZN(new_n525));
  NOR4_X1   g0325(.A1(new_n524), .A2(new_n525), .A3(KEYINPUT92), .A4(new_n511), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n337), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n509), .A2(new_n304), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n521), .A2(new_n522), .B1(new_n529), .B2(new_n490), .ZN(new_n530));
  INV_X1    g0330(.A(new_n294), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n329), .A2(KEYINPUT75), .ZN(new_n532));
  INV_X1    g0332(.A(G116), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n533), .B1(new_n203), .B2(G33), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n427), .B(new_n535), .C1(new_n294), .C2(new_n297), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n290), .A2(new_n210), .B1(G20), .B2(new_n533), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G283), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n538), .B(new_n204), .C1(G33), .C2(new_n220), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT20), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n537), .A2(KEYINPUT20), .A3(new_n539), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n534), .B(new_n536), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  MUX2_X1   g0343(.A(G257), .B(G264), .S(G1698), .Z(new_n544));
  NAND3_X1  g0344(.A1(new_n544), .A2(new_n409), .A3(new_n376), .ZN(new_n545));
  XNOR2_X1  g0345(.A(KEYINPUT89), .B(G303), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n486), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n267), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n267), .B(G270), .C1(new_n492), .C2(new_n494), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n503), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(G200), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT90), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n543), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n548), .A2(new_n550), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(G190), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n552), .B1(new_n543), .B2(new_n551), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT21), .ZN(new_n559));
  OAI21_X1  g0359(.A(G169), .B1(new_n548), .B2(new_n550), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n559), .B1(new_n543), .B2(new_n560), .ZN(new_n561));
  OR2_X1    g0361(.A1(new_n548), .A2(new_n550), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n562), .A2(KEYINPUT21), .A3(G169), .A4(new_n542), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n554), .A2(G179), .A3(new_n542), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n561), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(KEYINPUT91), .B1(new_n558), .B2(new_n565), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n561), .A2(new_n563), .A3(new_n564), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n543), .A2(new_n551), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT90), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n569), .A2(new_n555), .A3(new_n553), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT91), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n567), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n409), .A2(new_n204), .A3(G68), .A4(new_n376), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT19), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n287), .B2(new_n220), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n371), .A2(new_n373), .ZN(new_n577));
  AOI21_X1  g0377(.A(G20), .B1(new_n577), .B2(KEYINPUT19), .ZN(new_n578));
  NOR3_X1   g0378(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n574), .B(new_n576), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n291), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n298), .A2(new_n288), .ZN(new_n582));
  AOI211_X1 g0382(.A(new_n291), .B(new_n329), .C1(new_n203), .C2(G33), .ZN(new_n583));
  INV_X1    g0383(.A(new_n288), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n581), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(G238), .A2(G1698), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n227), .B2(G1698), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n588), .A2(new_n409), .A3(new_n376), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n267), .B1(new_n589), .B2(new_n480), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n498), .A2(new_n274), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n219), .B1(new_n497), .B2(G1), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n267), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n308), .B1(new_n590), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n590), .A2(new_n594), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n306), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n586), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n580), .A2(new_n291), .B1(new_n298), .B2(new_n288), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n589), .A2(new_n480), .ZN(new_n600));
  OAI211_X1 g0400(.A(G190), .B(new_n593), .C1(new_n600), .C2(new_n267), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n583), .A2(G87), .ZN(new_n602));
  OAI21_X1  g0402(.A(G200), .B1(new_n590), .B2(new_n594), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n599), .A2(new_n601), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n598), .A2(KEYINPUT88), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT88), .B1(new_n598), .B2(new_n604), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT86), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n376), .A2(new_n378), .A3(G250), .A4(G1698), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT83), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT83), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n254), .A2(new_n611), .A3(G250), .A4(G1698), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n227), .A2(G1698), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n409), .A2(new_n376), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT4), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g0417(.A1(KEYINPUT4), .A2(G244), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n376), .A2(new_n378), .A3(new_n618), .A4(new_n255), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n538), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n613), .A2(new_n617), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n386), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n267), .B(G257), .C1(new_n492), .C2(new_n494), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n503), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n608), .B1(new_n627), .B2(G179), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n625), .B1(new_n622), .B2(new_n386), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n629), .A2(KEYINPUT86), .A3(new_n306), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n627), .A2(new_n308), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n258), .A2(KEYINPUT6), .A3(G97), .ZN(new_n632));
  XOR2_X1   g0432(.A(G97), .B(G107), .Z(new_n633));
  OAI21_X1  g0433(.A(new_n632), .B1(new_n633), .B2(KEYINPUT6), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n634), .A2(G20), .B1(G77), .B2(new_n284), .ZN(new_n635));
  INV_X1    g0435(.A(new_n446), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n375), .B1(new_n438), .B2(new_n439), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n636), .B1(new_n637), .B2(new_n378), .ZN(new_n638));
  AOI21_X1  g0438(.A(KEYINPUT7), .B1(new_n486), .B2(new_n204), .ZN(new_n639));
  OAI21_X1  g0439(.A(G107), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n427), .B1(new_n635), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n329), .A2(new_n220), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n642), .B1(new_n476), .B2(new_n220), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n628), .A2(new_n630), .A3(new_n631), .A4(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n620), .B1(new_n616), .B2(new_n615), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n267), .B1(new_n647), .B2(new_n613), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n304), .B1(new_n648), .B2(new_n625), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n623), .A2(new_n337), .A3(new_n626), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n651), .A2(KEYINPUT85), .A3(new_n644), .ZN(new_n652));
  AOI21_X1  g0452(.A(KEYINPUT85), .B1(new_n651), .B2(new_n644), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n646), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(KEYINPUT87), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT87), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n646), .B(new_n656), .C1(new_n652), .C2(new_n653), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n607), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  AND4_X1   g0458(.A1(new_n473), .A2(new_n530), .A3(new_n573), .A4(new_n658), .ZN(G372));
  INV_X1    g0459(.A(new_n336), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n454), .A2(new_n464), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n392), .A2(G169), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT14), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n664), .A2(new_n395), .A3(new_n394), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n307), .A2(new_n302), .A3(new_n309), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n665), .A2(new_n363), .B1(new_n666), .B2(new_n402), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT94), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n470), .B(new_n471), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n402), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n398), .B1(new_n670), .B2(new_n310), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(KEYINPUT94), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n662), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n344), .A2(new_n345), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n660), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n519), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n567), .B1(new_n676), .B2(new_n490), .ZN(new_n677));
  AOI21_X1  g0477(.A(G200), .B1(new_n623), .B2(new_n626), .ZN(new_n678));
  AOI211_X1 g0478(.A(G190), .B(new_n625), .C1(new_n622), .C2(new_n386), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n644), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT85), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n651), .A2(KEYINPUT85), .A3(new_n644), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n598), .A2(new_n604), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n685), .B1(new_n529), .B2(new_n490), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n677), .A2(new_n684), .A3(new_n646), .A4(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n598), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n646), .A2(new_n685), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT26), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(KEYINPUT26), .B1(new_n607), .B2(new_n646), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n687), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n473), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n675), .A2(new_n694), .ZN(G369));
  NAND2_X1  g0495(.A1(new_n293), .A2(new_n204), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n697));
  XOR2_X1   g0497(.A(new_n697), .B(KEYINPUT95), .Z(new_n698));
  INV_X1    g0498(.A(G213), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n699), .B1(new_n696), .B2(KEYINPUT27), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G343), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n567), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n676), .A2(new_n490), .ZN(new_n705));
  INV_X1    g0505(.A(new_n703), .ZN(new_n706));
  AOI22_X1  g0506(.A1(new_n530), .A2(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n543), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n573), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT96), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n709), .A2(new_n567), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n521), .A2(new_n522), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n529), .A2(new_n490), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n490), .A2(new_n706), .ZN(new_n718));
  OAI22_X1  g0518(.A1(new_n717), .A2(new_n718), .B1(new_n715), .B2(new_n706), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n708), .B1(new_n566), .B2(new_n572), .ZN(new_n720));
  OAI21_X1  g0520(.A(KEYINPUT96), .B1(new_n720), .B2(new_n712), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n714), .A2(new_n719), .A3(new_n721), .A4(G330), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n722), .A2(KEYINPUT97), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(KEYINPUT97), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n707), .B1(new_n723), .B2(new_n724), .ZN(G399));
  INV_X1    g0525(.A(KEYINPUT88), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n685), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n598), .A2(KEYINPUT88), .A3(new_n604), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n630), .ZN(new_n730));
  OAI22_X1  g0530(.A1(new_n629), .A2(G169), .B1(new_n641), .B2(new_n643), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT86), .B1(new_n629), .B2(new_n306), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n690), .B1(new_n729), .B2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n685), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n733), .A2(new_n690), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n598), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n703), .B1(new_n738), .B2(new_n687), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT99), .B1(new_n739), .B2(KEYINPUT29), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n684), .A2(new_n646), .A3(new_n686), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n565), .B1(new_n521), .B2(new_n522), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n733), .B(new_n690), .C1(new_n605), .C2(new_n606), .ZN(new_n744));
  OAI21_X1  g0544(.A(KEYINPUT26), .B1(new_n646), .B2(new_n685), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n744), .A2(new_n745), .A3(new_n598), .ZN(new_n746));
  OAI211_X1 g0546(.A(KEYINPUT29), .B(new_n706), .C1(new_n743), .C2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n693), .A2(new_n706), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT99), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT29), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n740), .A2(new_n747), .A3(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G330), .ZN(new_n753));
  AND3_X1   g0553(.A1(new_n530), .A2(new_n573), .A3(new_n706), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n658), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n562), .A2(new_n306), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n596), .A2(new_n514), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n756), .A2(new_n629), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(KEYINPUT98), .A2(KEYINPUT30), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n759), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n756), .A2(new_n629), .A3(new_n757), .A4(new_n761), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n554), .A2(new_n596), .A3(G179), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(new_n509), .A3(new_n627), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n760), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(new_n703), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n766), .A2(KEYINPUT31), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(KEYINPUT31), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n753), .B1(new_n755), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n752), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT100), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n752), .A2(KEYINPUT100), .A3(new_n771), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n774), .A2(new_n203), .A3(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n207), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(G41), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n579), .A2(new_n533), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n778), .A2(new_n779), .A3(new_n203), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n780), .B1(new_n214), .B2(new_n778), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT28), .Z(new_n782));
  NAND2_X1  g0582(.A1(new_n776), .A2(new_n782), .ZN(G364));
  NOR2_X1   g0583(.A1(new_n292), .A2(G20), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n203), .B1(new_n784), .B2(G45), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n778), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n714), .A2(new_n721), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G13), .A2(G33), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n777), .A2(new_n486), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n794), .A2(G355), .B1(new_n533), .B2(new_n777), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT101), .Z(new_n796));
  NOR2_X1   g0596(.A1(new_n249), .A2(new_n497), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n777), .A2(new_n441), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(G45), .B2(new_n213), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n796), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n210), .B1(G20), .B2(new_n308), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n792), .A2(new_n801), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT102), .Z(new_n803));
  NOR2_X1   g0603(.A1(new_n204), .A2(new_n306), .ZN(new_n804));
  NOR2_X1   g0604(.A1(G190), .A2(G200), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G311), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n805), .A2(G20), .A3(new_n306), .ZN(new_n808));
  INV_X1    g0608(.A(G329), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n806), .A2(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n804), .A2(G190), .A3(new_n304), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n254), .B(new_n810), .C1(G322), .C2(new_n812), .ZN(new_n813));
  NOR4_X1   g0613(.A1(new_n204), .A2(new_n304), .A3(G179), .A4(G190), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT104), .Z(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G283), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n804), .A2(G200), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(new_n337), .ZN(new_n818));
  NOR4_X1   g0618(.A1(new_n204), .A2(new_n337), .A3(new_n304), .A4(G179), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n818), .A2(G326), .B1(G303), .B2(new_n819), .ZN(new_n820));
  NOR3_X1   g0620(.A1(new_n337), .A2(G179), .A3(G200), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n204), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n804), .A2(new_n337), .A3(G200), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(KEYINPUT33), .B(G317), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G294), .A2(new_n823), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n813), .A2(new_n816), .A3(new_n820), .A4(new_n827), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n811), .B(KEYINPUT103), .Z(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(G58), .ZN(new_n831));
  INV_X1    g0631(.A(new_n808), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(G159), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(KEYINPUT32), .ZN(new_n834));
  INV_X1    g0634(.A(new_n806), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n486), .B1(new_n835), .B2(new_n282), .ZN(new_n836));
  INV_X1    g0636(.A(new_n819), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n837), .A2(new_n218), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(G68), .B2(new_n825), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n831), .A2(new_n834), .A3(new_n836), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n815), .A2(G107), .ZN(new_n841));
  AOI22_X1  g0641(.A1(G97), .A2(new_n823), .B1(new_n818), .B2(G50), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n841), .B(new_n842), .C1(KEYINPUT32), .C2(new_n833), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n828), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n800), .A2(new_n803), .B1(new_n801), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n788), .B1(new_n793), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n789), .A2(new_n753), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n714), .A2(G330), .A3(new_n721), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n787), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT105), .Z(G396));
  NAND2_X1  g0651(.A1(new_n703), .A2(new_n302), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n305), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n310), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n310), .A2(new_n703), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n748), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n855), .B1(new_n853), .B2(new_n310), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n693), .A2(new_n706), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n787), .B1(new_n771), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n771), .B2(new_n861), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n818), .A2(G137), .B1(new_n835), .B2(G159), .ZN(new_n864));
  INV_X1    g0664(.A(G143), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n864), .B1(new_n323), .B2(new_n824), .C1(new_n829), .C2(new_n865), .ZN(new_n866));
  XOR2_X1   g0666(.A(new_n866), .B(KEYINPUT106), .Z(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(KEYINPUT34), .ZN(new_n868));
  INV_X1    g0668(.A(new_n815), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n869), .A2(new_n225), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n441), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(G132), .B2(new_n832), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n823), .A2(G58), .B1(G50), .B2(new_n819), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n868), .A2(new_n871), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n867), .A2(KEYINPUT34), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n869), .A2(new_n218), .ZN(new_n877));
  INV_X1    g0677(.A(G294), .ZN(new_n878));
  OAI22_X1  g0678(.A1(new_n811), .A2(new_n878), .B1(new_n807), .B2(new_n808), .ZN(new_n879));
  AOI211_X1 g0679(.A(new_n254), .B(new_n879), .C1(G116), .C2(new_n835), .ZN(new_n880));
  AOI22_X1  g0680(.A1(G97), .A2(new_n823), .B1(new_n818), .B2(G303), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n825), .A2(G283), .B1(new_n819), .B2(G107), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  OAI22_X1  g0683(.A1(new_n875), .A2(new_n876), .B1(new_n877), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n801), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n801), .A2(new_n790), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n788), .B1(new_n353), .B2(new_n886), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n885), .B(new_n887), .C1(new_n791), .C2(new_n859), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n863), .A2(new_n888), .ZN(G384));
  OR2_X1    g0689(.A1(new_n634), .A2(KEYINPUT35), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n634), .A2(KEYINPUT35), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n890), .A2(G116), .A3(new_n212), .A4(new_n891), .ZN(new_n892));
  XOR2_X1   g0692(.A(new_n892), .B(KEYINPUT36), .Z(new_n893));
  OR3_X1    g0693(.A1(new_n228), .A2(new_n213), .A3(new_n429), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n331), .A2(G68), .ZN(new_n895));
  AOI211_X1 g0695(.A(new_n203), .B(G13), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n658), .A2(new_n754), .B1(new_n768), .B2(new_n767), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n363), .A2(new_n703), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT107), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n398), .A2(new_n402), .A3(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n899), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n665), .B2(new_n670), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n859), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT40), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n898), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n455), .B1(new_n458), .B2(new_n459), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n445), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n426), .B1(new_n444), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n910), .A2(new_n701), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n472), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n468), .B1(new_n910), .B2(new_n701), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n423), .A2(new_n910), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT37), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n462), .A2(new_n418), .A3(new_n422), .ZN(new_n916));
  INV_X1    g0716(.A(new_n701), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n462), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT37), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n916), .A2(new_n918), .A3(new_n919), .A4(new_n468), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n915), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n912), .A2(new_n921), .A3(KEYINPUT38), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n470), .A2(new_n471), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(KEYINPUT108), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT108), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n470), .A2(new_n925), .A3(new_n471), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n924), .A2(new_n454), .A3(new_n464), .A4(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n918), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n916), .A2(new_n468), .A3(new_n918), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT37), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n927), .A2(new_n928), .B1(new_n920), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n922), .B1(new_n931), .B2(KEYINPUT38), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n912), .A2(new_n921), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT38), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n922), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n857), .B1(new_n903), .B2(new_n901), .ZN(new_n937));
  INV_X1    g0737(.A(new_n657), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n656), .B1(new_n684), .B2(new_n646), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n729), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n530), .A2(new_n573), .A3(new_n706), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n769), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n936), .A2(new_n937), .A3(new_n942), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n907), .A2(new_n932), .B1(new_n943), .B2(new_n906), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n473), .A2(new_n942), .ZN(new_n946));
  OAI21_X1  g0746(.A(G330), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(new_n946), .B2(new_n945), .ZN(new_n948));
  AND3_X1   g0748(.A1(new_n912), .A2(new_n921), .A3(KEYINPUT38), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT38), .B1(new_n912), .B2(new_n921), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(KEYINPUT39), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n665), .A2(new_n363), .A3(new_n706), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n926), .A2(new_n454), .A3(new_n464), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n925), .B1(new_n470), .B2(new_n471), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n928), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n930), .A2(new_n920), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n949), .B1(new_n934), .B2(new_n959), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n952), .B(new_n954), .C1(KEYINPUT39), .C2(new_n960), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n901), .A2(new_n903), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(new_n860), .B2(new_n856), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n963), .A2(new_n936), .B1(new_n661), .B2(new_n701), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n740), .A2(new_n473), .A3(new_n747), .A4(new_n751), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n675), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n965), .B(new_n967), .Z(new_n968));
  OAI22_X1  g0768(.A1(new_n948), .A2(new_n968), .B1(new_n203), .B2(new_n784), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n948), .A2(new_n968), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n897), .B1(new_n969), .B2(new_n970), .ZN(G367));
  INV_X1    g0771(.A(new_n798), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n240), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n802), .B1(new_n207), .B2(new_n288), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n787), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n830), .A2(new_n546), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n819), .A2(G116), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT46), .ZN(new_n978));
  INV_X1    g0778(.A(new_n818), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n979), .A2(new_n807), .B1(new_n258), .B2(new_n822), .ZN(new_n980));
  INV_X1    g0780(.A(new_n814), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n981), .A2(new_n220), .B1(new_n824), .B2(new_n878), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(G283), .ZN(new_n984));
  INV_X1    g0784(.A(G317), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n806), .A2(new_n984), .B1(new_n808), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n986), .A2(new_n441), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n976), .A2(new_n978), .A3(new_n983), .A4(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n822), .A2(new_n225), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(G150), .B2(new_n812), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT111), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n825), .A2(G159), .B1(new_n835), .B2(G50), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n991), .A2(KEYINPUT110), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(KEYINPUT110), .B2(new_n991), .ZN(new_n995));
  INV_X1    g0795(.A(G137), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n254), .B1(new_n808), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(new_n818), .B2(G143), .ZN(new_n998));
  AOI22_X1  g0798(.A1(G58), .A2(new_n819), .B1(new_n282), .B2(new_n814), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n998), .B(new_n999), .C1(new_n993), .C2(new_n992), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n988), .B1(new_n995), .B2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g0801(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n1002));
  XNOR2_X1  g0802(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n975), .B1(new_n1003), .B2(new_n801), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n792), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n599), .A2(new_n602), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n703), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n735), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n688), .A2(new_n1006), .A3(new_n703), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1004), .B1(new_n1005), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n530), .A2(new_n704), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n719), .B2(new_n704), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(new_n848), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n705), .A2(new_n706), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1013), .A2(new_n1017), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n646), .B1(new_n644), .B2(new_n706), .C1(new_n652), .C2(new_n653), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n733), .A2(new_n703), .ZN(new_n1020));
  XOR2_X1   g0820(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n1021));
  NAND4_X1  g0821(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1021), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1023), .B1(new_n707), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n707), .A2(new_n1024), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT45), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(KEYINPUT45), .B1(new_n707), .B2(new_n1024), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1022), .B(new_n1025), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n723), .B2(new_n724), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n722), .A2(KEYINPUT97), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1026), .B(new_n1027), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n722), .A2(KEYINPUT97), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1031), .A2(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1016), .A2(new_n1037), .B1(new_n774), .B2(new_n775), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n778), .B(KEYINPUT41), .Z(new_n1039));
  OAI21_X1  g0839(.A(new_n785), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1024), .A2(new_n530), .A3(new_n704), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1041), .A2(KEYINPUT42), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n684), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n646), .B1(new_n1043), .B2(new_n715), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n1041), .A2(KEYINPUT42), .B1(new_n706), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1010), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT43), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1010), .A2(KEYINPUT43), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1046), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1042), .A2(new_n1045), .A3(new_n1048), .A4(new_n1047), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1032), .A2(new_n1034), .A3(new_n1024), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1012), .B1(new_n1040), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(G387));
  AND3_X1   g0859(.A1(new_n752), .A2(KEYINPUT100), .A3(new_n771), .ZN(new_n1060));
  AOI21_X1  g0860(.A(KEYINPUT100), .B1(new_n752), .B2(new_n771), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1016), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n774), .A2(new_n775), .A3(new_n1015), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1062), .A2(new_n1063), .A3(new_n778), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1016), .A2(new_n786), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n794), .A2(new_n779), .B1(new_n258), .B2(new_n777), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n244), .A2(new_n497), .ZN(new_n1067));
  AOI211_X1 g0867(.A(G45), .B(new_n779), .C1(G68), .C2(G77), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n286), .ZN(new_n1069));
  AOI21_X1  g0869(.A(KEYINPUT50), .B1(new_n1069), .B2(new_n331), .ZN(new_n1070));
  AND3_X1   g0870(.A1(new_n1069), .A2(KEYINPUT50), .A3(new_n331), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1068), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n798), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1066), .B1(new_n1067), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n788), .B1(new_n1074), .B2(new_n803), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(G159), .A2(new_n818), .B1(new_n825), .B2(new_n1069), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n228), .B2(new_n837), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n872), .B1(new_n823), .B2(new_n584), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n835), .A2(G68), .B1(new_n832), .B2(G150), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(new_n331), .C2(new_n811), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n1077), .B(new_n1080), .C1(G97), .C2(new_n815), .ZN(new_n1081));
  INV_X1    g0881(.A(G326), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n872), .B1(new_n1082), .B2(new_n808), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n818), .A2(G322), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n825), .A2(G311), .B1(new_n835), .B2(new_n546), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1084), .B(new_n1085), .C1(new_n829), .C2(new_n985), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT48), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n823), .A2(G283), .B1(G294), .B2(new_n819), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT49), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1083), .B(new_n1093), .C1(G116), .C2(new_n814), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1081), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n801), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n1075), .B1(new_n719), .B2(new_n1005), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n1065), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1064), .A2(new_n1099), .ZN(G393));
  INV_X1    g0900(.A(new_n778), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1015), .B1(new_n774), .B2(new_n775), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1101), .B1(new_n1102), .B2(new_n1037), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n1031), .A2(new_n1036), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1062), .A2(KEYINPUT115), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(KEYINPUT115), .B1(new_n1062), .B2(new_n1104), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1103), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1024), .A2(new_n1005), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT113), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n802), .B1(new_n220), .B2(new_n207), .C1(new_n972), .C2(new_n252), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n787), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(G150), .A2(new_n818), .B1(new_n812), .B2(G159), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT51), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n441), .B1(new_n865), .B2(new_n808), .C1(new_n286), .C2(new_n806), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n822), .A2(new_n353), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n1117), .B1(new_n225), .B2(new_n837), .C1(new_n331), .C2(new_n824), .ZN(new_n1118));
  NOR4_X1   g0918(.A1(new_n1114), .A2(new_n877), .A3(new_n1115), .A4(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  OR2_X1    g0920(.A1(new_n1120), .A2(KEYINPUT114), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n979), .A2(new_n985), .B1(new_n807), .B2(new_n811), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT52), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n486), .B1(new_n806), .B2(new_n878), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(G322), .B2(new_n832), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n837), .A2(new_n984), .B1(new_n533), .B2(new_n822), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n546), .B2(new_n825), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1123), .A2(new_n841), .A3(new_n1125), .A4(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1120), .A2(KEYINPUT114), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1121), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1112), .B1(new_n1130), .B2(new_n801), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1037), .A2(new_n786), .B1(new_n1110), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1108), .A2(new_n1132), .ZN(G390));
  NAND2_X1  g0933(.A1(new_n860), .A2(new_n856), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n904), .B1(new_n770), .B2(new_n859), .ZN(new_n1135));
  NOR4_X1   g0935(.A1(new_n898), .A2(new_n962), .A3(new_n753), .A4(new_n857), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n706), .B(new_n854), .C1(new_n743), .C2(new_n746), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n856), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT116), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1138), .A2(KEYINPUT116), .A3(new_n856), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n942), .A2(G330), .A3(new_n859), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n962), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n770), .A2(new_n859), .A3(new_n904), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1143), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1137), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n770), .A2(new_n473), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n966), .A2(new_n675), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1148), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT117), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n959), .A2(new_n934), .ZN(new_n1154));
  AOI21_X1  g0954(.A(KEYINPUT39), .B1(new_n1154), .B2(new_n922), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n935), .A2(KEYINPUT39), .A3(new_n922), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n1155), .A2(new_n1156), .B1(new_n963), .B2(new_n954), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1138), .A2(KEYINPUT116), .A3(new_n856), .ZN(new_n1158));
  AOI21_X1  g0958(.A(KEYINPUT116), .B1(new_n1138), .B2(new_n856), .ZN(new_n1159));
  NOR3_X1   g0959(.A1(new_n1158), .A2(new_n1159), .A3(new_n962), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n932), .A2(new_n953), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1157), .B(new_n1146), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1141), .A2(new_n904), .A3(new_n1142), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1161), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1146), .B1(new_n1166), .B2(new_n1157), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1152), .B(new_n1153), .C1(new_n1163), .C2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1157), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n1136), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1150), .B1(new_n1137), .B2(new_n1147), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1170), .B(new_n1162), .C1(new_n1171), .C2(KEYINPUT117), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1168), .A2(new_n778), .A3(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1170), .A2(new_n786), .A3(new_n1162), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n790), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n886), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n486), .B1(new_n808), .B2(new_n878), .C1(new_n811), .C2(new_n533), .ZN(new_n1177));
  NOR4_X1   g0977(.A1(new_n870), .A2(new_n838), .A3(new_n1177), .A4(new_n1116), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n818), .A2(G283), .B1(new_n835), .B2(G97), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n258), .B2(new_n824), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT119), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(KEYINPUT54), .B(G143), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n823), .A2(G159), .B1(new_n835), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n996), .B2(new_n824), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT118), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n819), .A2(G150), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT53), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n486), .B1(new_n812), .B2(G132), .ZN(new_n1189));
  INV_X1    g0989(.A(G125), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1189), .B1(new_n1190), .B2(new_n808), .ZN(new_n1191));
  INV_X1    g0991(.A(G128), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n979), .A2(new_n1192), .B1(new_n331), .B2(new_n981), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1188), .A2(new_n1191), .A3(new_n1193), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n1178), .A2(new_n1181), .B1(new_n1186), .B2(new_n1194), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n787), .B1(new_n1069), .B2(new_n1176), .C1(new_n1195), .C2(new_n1097), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT120), .Z(new_n1197));
  NAND2_X1  g0997(.A1(new_n1175), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1174), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1173), .A2(new_n1200), .ZN(G378));
  NAND4_X1  g1001(.A1(new_n932), .A2(KEYINPUT40), .A3(new_n942), .A4(new_n937), .ZN(new_n1202));
  NOR3_X1   g1002(.A1(new_n951), .A2(new_n898), .A3(new_n905), .ZN(new_n1203));
  OAI211_X1 g1003(.A(G330), .B(new_n1202), .C1(new_n1203), .C2(KEYINPUT40), .ZN(new_n1204));
  XOR2_X1   g1004(.A(KEYINPUT123), .B(KEYINPUT56), .Z(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n336), .B1(new_n344), .B2(new_n345), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n334), .A2(new_n917), .ZN(new_n1208));
  XOR2_X1   g1008(.A(new_n1208), .B(KEYINPUT55), .Z(new_n1209));
  AND2_X1   g1009(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1206), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1213), .A2(new_n1205), .A3(new_n1214), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1212), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1204), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n965), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1212), .A2(new_n1215), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n943), .A2(new_n906), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1219), .A2(new_n1220), .A3(G330), .A4(new_n1202), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1217), .A2(new_n1218), .A3(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1218), .B1(new_n1217), .B2(new_n1221), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1219), .A2(new_n790), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1176), .A2(G50), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n812), .A2(G107), .B1(G283), .B2(new_n832), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n288), .B2(new_n806), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n989), .B(new_n1228), .C1(new_n282), .C2(new_n819), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n979), .A2(new_n533), .B1(new_n428), .B2(new_n981), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(G97), .B2(new_n825), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n441), .A2(G41), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1229), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT58), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  AOI211_X1 g1035(.A(G50), .B(new_n1232), .C1(new_n375), .C2(new_n491), .ZN(new_n1236));
  XOR2_X1   g1036(.A(new_n1236), .B(KEYINPUT121), .Z(new_n1237));
  AND2_X1   g1037(.A1(new_n1235), .A2(new_n1237), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n811), .A2(new_n1192), .B1(new_n806), .B2(new_n996), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n825), .A2(G132), .B1(new_n819), .B2(new_n1183), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n1190), .B2(new_n979), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n1239), .B(new_n1241), .C1(G150), .C2(new_n823), .ZN(new_n1242));
  XOR2_X1   g1042(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n1243));
  NOR2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n814), .A2(G159), .ZN(new_n1246));
  AOI211_X1 g1046(.A(G33), .B(G41), .C1(new_n832), .C2(G124), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n1238), .B1(new_n1234), .B2(new_n1233), .C1(new_n1244), .C2(new_n1248), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n788), .B(new_n1226), .C1(new_n1249), .C2(new_n801), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1224), .A2(new_n786), .B1(new_n1225), .B2(new_n1250), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1163), .A2(new_n1167), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1150), .B1(new_n1252), .B2(new_n1148), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1219), .B1(new_n944), .B2(G330), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1204), .A2(new_n1216), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n965), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1217), .A2(new_n1218), .A3(new_n1221), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1256), .A2(KEYINPUT57), .A3(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n778), .B1(new_n1253), .B2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1170), .A2(new_n1162), .A3(new_n1148), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1151), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT57), .B1(new_n1224), .B2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1251), .B1(new_n1259), .B2(new_n1262), .ZN(G375));
  NAND2_X1  g1063(.A1(new_n1148), .A2(new_n786), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n787), .B1(G68), .B2(new_n1176), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n811), .A2(new_n984), .B1(new_n806), .B2(new_n258), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n254), .B(new_n1266), .C1(G303), .C2(new_n832), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n815), .A2(G77), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n584), .A2(new_n823), .B1(new_n825), .B2(G116), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n818), .A2(G294), .B1(G97), .B2(new_n819), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1267), .A2(new_n1268), .A3(new_n1269), .A4(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n830), .A2(G137), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n825), .A2(new_n1183), .B1(G58), .B2(new_n814), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(G50), .A2(new_n823), .B1(new_n818), .B2(G132), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n872), .B1(G150), .B2(new_n835), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1272), .A2(new_n1273), .A3(new_n1274), .A4(new_n1275), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n819), .A2(G159), .B1(new_n832), .B2(G128), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1277), .B(KEYINPUT124), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1271), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1265), .B1(new_n1279), .B2(new_n801), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n904), .B2(new_n791), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1264), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1039), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1137), .A2(new_n1150), .A3(new_n1147), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1152), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1283), .A2(new_n1286), .ZN(G381));
  NOR2_X1   g1087(.A1(G393), .A2(G396), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NOR4_X1   g1089(.A1(G390), .A2(new_n1289), .A3(G384), .A4(G381), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1101), .B1(new_n1291), .B2(new_n1252), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1199), .B1(new_n1292), .B2(new_n1168), .ZN(new_n1293));
  INV_X1    g1093(.A(G375), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1290), .A2(new_n1058), .A3(new_n1293), .A4(new_n1294), .ZN(G407));
  NAND2_X1  g1095(.A1(new_n702), .A2(G213), .ZN(new_n1296));
  OR3_X1    g1096(.A1(G375), .A2(G378), .A3(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(G407), .A2(new_n1297), .A3(G213), .ZN(G409));
  OR2_X1    g1098(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1299));
  OAI22_X1  g1099(.A1(new_n1104), .A2(new_n1015), .B1(new_n1061), .B2(new_n1060), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1284), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1299), .B1(new_n1301), .B2(new_n785), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1108), .B(new_n1132), .C1(new_n1302), .C2(new_n1012), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n778), .B1(new_n1062), .B2(new_n1104), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT115), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1305), .B1(new_n1102), .B2(new_n1037), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1304), .B1(new_n1306), .B2(new_n1105), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1132), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1058), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1303), .A2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT125), .B1(G390), .B2(new_n1058), .ZN(new_n1311));
  AND2_X1   g1111(.A1(G393), .A2(G396), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1312), .A2(new_n1288), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1310), .B1(new_n1311), .B2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1313), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1315), .A2(new_n1303), .A3(new_n1309), .A4(KEYINPUT125), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1314), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  OAI211_X1 g1118(.A(G378), .B(new_n1251), .C1(new_n1259), .C2(new_n1262), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1224), .A2(new_n1261), .A3(new_n1284), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1225), .A2(new_n1250), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1321), .B1(new_n1322), .B2(new_n785), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1293), .B1(new_n1320), .B2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1319), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n1296), .ZN(new_n1326));
  INV_X1    g1126(.A(G384), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1150), .A2(new_n1137), .A3(new_n1147), .A4(KEYINPUT60), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(new_n778), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1152), .A2(KEYINPUT60), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1329), .B1(new_n1330), .B2(new_n1285), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1327), .B1(new_n1331), .B2(new_n1282), .ZN(new_n1332));
  AND2_X1   g1132(.A1(new_n1328), .A2(new_n778), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT60), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1171), .A2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1285), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1333), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1337), .A2(G384), .A3(new_n1283), .ZN(new_n1338));
  INV_X1    g1138(.A(G2897), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1296), .A2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1340), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1332), .A2(new_n1338), .A3(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1341), .B1(new_n1332), .B2(new_n1338), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1326), .A2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT61), .ZN(new_n1347));
  AOI21_X1  g1147(.A(KEYINPUT126), .B1(new_n1346), .B2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1332), .A2(new_n1338), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1349), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1325), .A2(new_n1296), .A3(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(KEYINPUT62), .ZN(new_n1352));
  AOI22_X1  g1152(.A1(new_n1319), .A2(new_n1324), .B1(G213), .B2(new_n702), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT62), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1353), .A2(new_n1354), .A3(new_n1350), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1352), .A2(new_n1355), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1318), .B1(new_n1348), .B2(new_n1356), .ZN(new_n1357));
  AND4_X1   g1157(.A1(KEYINPUT63), .A2(new_n1325), .A3(new_n1296), .A4(new_n1350), .ZN(new_n1358));
  AOI21_X1  g1158(.A(KEYINPUT63), .B1(new_n1353), .B2(new_n1350), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1317), .B1(new_n1358), .B2(new_n1359), .ZN(new_n1360));
  INV_X1    g1160(.A(KEYINPUT126), .ZN(new_n1361));
  AND3_X1   g1161(.A1(new_n1314), .A2(new_n1316), .A3(new_n1361), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1349), .A2(new_n1340), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1363), .A2(new_n1342), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1347), .B1(new_n1353), .B2(new_n1364), .ZN(new_n1365));
  NOR2_X1   g1165(.A1(new_n1362), .A2(new_n1365), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1360), .A2(new_n1366), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1357), .A2(new_n1367), .ZN(G405));
  NAND2_X1  g1168(.A1(G375), .A2(new_n1293), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1369), .A2(new_n1319), .ZN(new_n1370));
  XNOR2_X1  g1170(.A(new_n1370), .B(new_n1350), .ZN(new_n1371));
  XNOR2_X1  g1171(.A(new_n1371), .B(new_n1318), .ZN(G402));
endmodule


