

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U552 ( .A(KEYINPUT99), .ZN(n740) );
  NOR2_X1 U553 ( .A1(G651), .A2(n643), .ZN(n650) );
  XNOR2_X1 U554 ( .A(KEYINPUT23), .B(KEYINPUT65), .ZN(n527) );
  XNOR2_X1 U555 ( .A(n528), .B(n527), .ZN(n531) );
  XOR2_X1 U556 ( .A(KEYINPUT0), .B(G543), .Z(n643) );
  NAND2_X1 U557 ( .A1(n650), .A2(G50), .ZN(n520) );
  XOR2_X1 U558 ( .A(G651), .B(KEYINPUT66), .Z(n521) );
  NOR2_X1 U559 ( .A1(G543), .A2(n521), .ZN(n518) );
  XOR2_X1 U560 ( .A(KEYINPUT1), .B(n518), .Z(n587) );
  BUF_X1 U561 ( .A(n587), .Z(n658) );
  NAND2_X1 U562 ( .A1(G62), .A2(n658), .ZN(n519) );
  NAND2_X1 U563 ( .A1(n520), .A2(n519), .ZN(n525) );
  NOR2_X1 U564 ( .A1(G651), .A2(G543), .ZN(n649) );
  NAND2_X1 U565 ( .A1(n649), .A2(G88), .ZN(n523) );
  NOR2_X1 U566 ( .A1(n643), .A2(n521), .ZN(n653) );
  NAND2_X1 U567 ( .A1(G75), .A2(n653), .ZN(n522) );
  NAND2_X1 U568 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U569 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U570 ( .A(n526), .B(KEYINPUT82), .ZN(G166) );
  INV_X1 U571 ( .A(G166), .ZN(G303) );
  INV_X1 U572 ( .A(G2105), .ZN(n532) );
  AND2_X1 U573 ( .A1(n532), .A2(G2104), .ZN(n876) );
  NAND2_X1 U574 ( .A1(G101), .A2(n876), .ZN(n528) );
  NOR2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n529) );
  XOR2_X1 U576 ( .A(KEYINPUT17), .B(n529), .Z(n562) );
  BUF_X1 U577 ( .A(n562), .Z(n875) );
  NAND2_X1 U578 ( .A1(G137), .A2(n875), .ZN(n530) );
  AND2_X1 U579 ( .A1(n531), .A2(n530), .ZN(n692) );
  NOR2_X1 U580 ( .A1(G2104), .A2(n532), .ZN(n879) );
  NAND2_X1 U581 ( .A1(G125), .A2(n879), .ZN(n534) );
  AND2_X1 U582 ( .A1(G2105), .A2(G2104), .ZN(n880) );
  NAND2_X1 U583 ( .A1(G113), .A2(n880), .ZN(n533) );
  AND2_X1 U584 ( .A1(n534), .A2(n533), .ZN(n691) );
  AND2_X1 U585 ( .A1(n692), .A2(n691), .ZN(G160) );
  NAND2_X1 U586 ( .A1(n649), .A2(G85), .ZN(n536) );
  NAND2_X1 U587 ( .A1(G72), .A2(n653), .ZN(n535) );
  NAND2_X1 U588 ( .A1(n536), .A2(n535), .ZN(n540) );
  NAND2_X1 U589 ( .A1(n650), .A2(G47), .ZN(n538) );
  NAND2_X1 U590 ( .A1(G60), .A2(n658), .ZN(n537) );
  NAND2_X1 U591 ( .A1(n538), .A2(n537), .ZN(n539) );
  OR2_X1 U592 ( .A1(n540), .A2(n539), .ZN(G290) );
  NAND2_X1 U593 ( .A1(n650), .A2(G52), .ZN(n542) );
  NAND2_X1 U594 ( .A1(G64), .A2(n658), .ZN(n541) );
  NAND2_X1 U595 ( .A1(n542), .A2(n541), .ZN(n549) );
  XNOR2_X1 U596 ( .A(KEYINPUT68), .B(KEYINPUT9), .ZN(n547) );
  NAND2_X1 U597 ( .A1(n649), .A2(G90), .ZN(n545) );
  NAND2_X1 U598 ( .A1(G77), .A2(n653), .ZN(n543) );
  XOR2_X1 U599 ( .A(KEYINPUT67), .B(n543), .Z(n544) );
  NAND2_X1 U600 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U601 ( .A(n547), .B(n546), .Z(n548) );
  NOR2_X1 U602 ( .A1(n549), .A2(n548), .ZN(G171) );
  XOR2_X1 U603 ( .A(G2443), .B(KEYINPUT104), .Z(n551) );
  XNOR2_X1 U604 ( .A(G2451), .B(G2427), .ZN(n550) );
  XNOR2_X1 U605 ( .A(n551), .B(n550), .ZN(n555) );
  XOR2_X1 U606 ( .A(G2435), .B(G2438), .Z(n553) );
  XNOR2_X1 U607 ( .A(G2454), .B(G2430), .ZN(n552) );
  XNOR2_X1 U608 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U609 ( .A(n555), .B(n554), .Z(n557) );
  XNOR2_X1 U610 ( .A(G2446), .B(KEYINPUT102), .ZN(n556) );
  XNOR2_X1 U611 ( .A(n557), .B(n556), .ZN(n560) );
  XOR2_X1 U612 ( .A(G1341), .B(G1348), .Z(n558) );
  XNOR2_X1 U613 ( .A(KEYINPUT103), .B(n558), .ZN(n559) );
  XOR2_X1 U614 ( .A(n560), .B(n559), .Z(n561) );
  AND2_X1 U615 ( .A1(G14), .A2(n561), .ZN(G401) );
  AND2_X1 U616 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U617 ( .A(G57), .ZN(G237) );
  NAND2_X1 U618 ( .A1(G138), .A2(n562), .ZN(n564) );
  NAND2_X1 U619 ( .A1(G102), .A2(n876), .ZN(n563) );
  NAND2_X1 U620 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U621 ( .A(n565), .B(KEYINPUT90), .ZN(n569) );
  NAND2_X1 U622 ( .A1(G126), .A2(n879), .ZN(n567) );
  NAND2_X1 U623 ( .A1(G114), .A2(n880), .ZN(n566) );
  NAND2_X1 U624 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U625 ( .A1(n569), .A2(n568), .ZN(G164) );
  NAND2_X1 U626 ( .A1(G7), .A2(G661), .ZN(n570) );
  XNOR2_X1 U627 ( .A(n570), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U628 ( .A(KEYINPUT11), .B(KEYINPUT70), .Z(n572) );
  INV_X1 U629 ( .A(G223), .ZN(n828) );
  NAND2_X1 U630 ( .A1(G567), .A2(n828), .ZN(n571) );
  XNOR2_X1 U631 ( .A(n572), .B(n571), .ZN(G234) );
  NAND2_X1 U632 ( .A1(G81), .A2(n649), .ZN(n573) );
  XNOR2_X1 U633 ( .A(n573), .B(KEYINPUT12), .ZN(n574) );
  XNOR2_X1 U634 ( .A(n574), .B(KEYINPUT72), .ZN(n576) );
  NAND2_X1 U635 ( .A1(G68), .A2(n653), .ZN(n575) );
  NAND2_X1 U636 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U637 ( .A(KEYINPUT13), .B(n577), .Z(n581) );
  NAND2_X1 U638 ( .A1(n587), .A2(G56), .ZN(n578) );
  XNOR2_X1 U639 ( .A(n578), .B(KEYINPUT14), .ZN(n579) );
  XNOR2_X1 U640 ( .A(n579), .B(KEYINPUT71), .ZN(n580) );
  NOR2_X1 U641 ( .A1(n581), .A2(n580), .ZN(n583) );
  NAND2_X1 U642 ( .A1(n650), .A2(G43), .ZN(n582) );
  NAND2_X1 U643 ( .A1(n583), .A2(n582), .ZN(n966) );
  INV_X1 U644 ( .A(G860), .ZN(n617) );
  OR2_X1 U645 ( .A1(n966), .A2(n617), .ZN(G153) );
  XNOR2_X1 U646 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U647 ( .A1(G868), .A2(G301), .ZN(n584) );
  XNOR2_X1 U648 ( .A(n584), .B(KEYINPUT74), .ZN(n594) );
  NAND2_X1 U649 ( .A1(n649), .A2(G92), .ZN(n586) );
  NAND2_X1 U650 ( .A1(G79), .A2(n653), .ZN(n585) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n591) );
  NAND2_X1 U652 ( .A1(n650), .A2(G54), .ZN(n589) );
  NAND2_X1 U653 ( .A1(G66), .A2(n587), .ZN(n588) );
  NAND2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U656 ( .A(KEYINPUT15), .B(n592), .Z(n976) );
  OR2_X1 U657 ( .A1(G868), .A2(n976), .ZN(n593) );
  NAND2_X1 U658 ( .A1(n594), .A2(n593), .ZN(G284) );
  NAND2_X1 U659 ( .A1(n653), .A2(G76), .ZN(n598) );
  XOR2_X1 U660 ( .A(KEYINPUT4), .B(KEYINPUT75), .Z(n596) );
  NAND2_X1 U661 ( .A1(G89), .A2(n649), .ZN(n595) );
  XNOR2_X1 U662 ( .A(n596), .B(n595), .ZN(n597) );
  NAND2_X1 U663 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U664 ( .A(n599), .B(KEYINPUT5), .ZN(n600) );
  XNOR2_X1 U665 ( .A(KEYINPUT76), .B(n600), .ZN(n606) );
  XNOR2_X1 U666 ( .A(KEYINPUT77), .B(KEYINPUT6), .ZN(n604) );
  NAND2_X1 U667 ( .A1(n650), .A2(G51), .ZN(n602) );
  NAND2_X1 U668 ( .A1(G63), .A2(n658), .ZN(n601) );
  NAND2_X1 U669 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U670 ( .A(n604), .B(n603), .ZN(n605) );
  NAND2_X1 U671 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U672 ( .A(n607), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U673 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U674 ( .A1(n650), .A2(G53), .ZN(n609) );
  NAND2_X1 U675 ( .A1(G65), .A2(n658), .ZN(n608) );
  NAND2_X1 U676 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U677 ( .A1(n649), .A2(G91), .ZN(n611) );
  NAND2_X1 U678 ( .A1(G78), .A2(n653), .ZN(n610) );
  NAND2_X1 U679 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U680 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U681 ( .A(n614), .B(KEYINPUT69), .ZN(G299) );
  NAND2_X1 U682 ( .A1(G286), .A2(G868), .ZN(n616) );
  INV_X1 U683 ( .A(G868), .ZN(n672) );
  NAND2_X1 U684 ( .A1(G299), .A2(n672), .ZN(n615) );
  NAND2_X1 U685 ( .A1(n616), .A2(n615), .ZN(G297) );
  NAND2_X1 U686 ( .A1(n617), .A2(G559), .ZN(n618) );
  NAND2_X1 U687 ( .A1(n618), .A2(n976), .ZN(n619) );
  XNOR2_X1 U688 ( .A(n619), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U689 ( .A1(G868), .A2(n966), .ZN(n622) );
  NAND2_X1 U690 ( .A1(G868), .A2(n976), .ZN(n620) );
  NOR2_X1 U691 ( .A1(G559), .A2(n620), .ZN(n621) );
  NOR2_X1 U692 ( .A1(n622), .A2(n621), .ZN(G282) );
  NAND2_X1 U693 ( .A1(G123), .A2(n879), .ZN(n623) );
  XNOR2_X1 U694 ( .A(n623), .B(KEYINPUT18), .ZN(n625) );
  NAND2_X1 U695 ( .A1(n876), .A2(G99), .ZN(n624) );
  NAND2_X1 U696 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U697 ( .A1(G135), .A2(n875), .ZN(n627) );
  NAND2_X1 U698 ( .A1(G111), .A2(n880), .ZN(n626) );
  NAND2_X1 U699 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U700 ( .A1(n629), .A2(n628), .ZN(n915) );
  XNOR2_X1 U701 ( .A(G2096), .B(n915), .ZN(n631) );
  INV_X1 U702 ( .A(G2100), .ZN(n630) );
  NAND2_X1 U703 ( .A1(n631), .A2(n630), .ZN(G156) );
  NAND2_X1 U704 ( .A1(G559), .A2(n976), .ZN(n632) );
  XNOR2_X1 U705 ( .A(n632), .B(n966), .ZN(n669) );
  NOR2_X1 U706 ( .A1(G860), .A2(n669), .ZN(n641) );
  NAND2_X1 U707 ( .A1(n649), .A2(G93), .ZN(n634) );
  NAND2_X1 U708 ( .A1(G80), .A2(n653), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n634), .A2(n633), .ZN(n639) );
  NAND2_X1 U710 ( .A1(n650), .A2(G55), .ZN(n636) );
  NAND2_X1 U711 ( .A1(G67), .A2(n658), .ZN(n635) );
  NAND2_X1 U712 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U713 ( .A(KEYINPUT79), .B(n637), .Z(n638) );
  NOR2_X1 U714 ( .A1(n639), .A2(n638), .ZN(n671) );
  XNOR2_X1 U715 ( .A(n671), .B(KEYINPUT78), .ZN(n640) );
  XNOR2_X1 U716 ( .A(n641), .B(n640), .ZN(G145) );
  NAND2_X1 U717 ( .A1(G74), .A2(G651), .ZN(n642) );
  XNOR2_X1 U718 ( .A(n642), .B(KEYINPUT80), .ZN(n648) );
  NAND2_X1 U719 ( .A1(G49), .A2(n650), .ZN(n645) );
  NAND2_X1 U720 ( .A1(G87), .A2(n643), .ZN(n644) );
  NAND2_X1 U721 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U722 ( .A1(n658), .A2(n646), .ZN(n647) );
  NAND2_X1 U723 ( .A1(n648), .A2(n647), .ZN(G288) );
  NAND2_X1 U724 ( .A1(G86), .A2(n649), .ZN(n652) );
  NAND2_X1 U725 ( .A1(G48), .A2(n650), .ZN(n651) );
  NAND2_X1 U726 ( .A1(n652), .A2(n651), .ZN(n657) );
  NAND2_X1 U727 ( .A1(n653), .A2(G73), .ZN(n654) );
  XNOR2_X1 U728 ( .A(n654), .B(KEYINPUT2), .ZN(n655) );
  XNOR2_X1 U729 ( .A(n655), .B(KEYINPUT81), .ZN(n656) );
  NOR2_X1 U730 ( .A1(n657), .A2(n656), .ZN(n660) );
  NAND2_X1 U731 ( .A1(G61), .A2(n658), .ZN(n659) );
  NAND2_X1 U732 ( .A1(n660), .A2(n659), .ZN(G305) );
  XOR2_X1 U733 ( .A(KEYINPUT85), .B(KEYINPUT83), .Z(n661) );
  XNOR2_X1 U734 ( .A(G288), .B(n661), .ZN(n662) );
  XNOR2_X1 U735 ( .A(KEYINPUT19), .B(n662), .ZN(n664) );
  XNOR2_X1 U736 ( .A(G290), .B(KEYINPUT84), .ZN(n663) );
  XNOR2_X1 U737 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U738 ( .A(n671), .B(n665), .ZN(n667) );
  XNOR2_X1 U739 ( .A(G305), .B(G303), .ZN(n666) );
  XNOR2_X1 U740 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U741 ( .A(n668), .B(G299), .ZN(n897) );
  XNOR2_X1 U742 ( .A(n669), .B(n897), .ZN(n670) );
  NAND2_X1 U743 ( .A1(n670), .A2(G868), .ZN(n674) );
  NAND2_X1 U744 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U745 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U746 ( .A(KEYINPUT86), .B(n675), .Z(G295) );
  XOR2_X1 U747 ( .A(KEYINPUT21), .B(KEYINPUT87), .Z(n679) );
  NAND2_X1 U748 ( .A1(G2084), .A2(G2078), .ZN(n676) );
  XOR2_X1 U749 ( .A(KEYINPUT20), .B(n676), .Z(n677) );
  NAND2_X1 U750 ( .A1(n677), .A2(G2090), .ZN(n678) );
  XNOR2_X1 U751 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U752 ( .A(KEYINPUT88), .B(n680), .ZN(n681) );
  NAND2_X1 U753 ( .A1(n681), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U755 ( .A(KEYINPUT22), .B(KEYINPUT89), .Z(n683) );
  NAND2_X1 U756 ( .A1(G132), .A2(G82), .ZN(n682) );
  XNOR2_X1 U757 ( .A(n683), .B(n682), .ZN(n684) );
  NOR2_X1 U758 ( .A1(n684), .A2(G218), .ZN(n685) );
  NAND2_X1 U759 ( .A1(G96), .A2(n685), .ZN(n832) );
  NAND2_X1 U760 ( .A1(n832), .A2(G2106), .ZN(n689) );
  NAND2_X1 U761 ( .A1(G69), .A2(G120), .ZN(n686) );
  NOR2_X1 U762 ( .A1(G237), .A2(n686), .ZN(n687) );
  NAND2_X1 U763 ( .A1(G108), .A2(n687), .ZN(n833) );
  NAND2_X1 U764 ( .A1(n833), .A2(G567), .ZN(n688) );
  NAND2_X1 U765 ( .A1(n689), .A2(n688), .ZN(n834) );
  NAND2_X1 U766 ( .A1(G483), .A2(G661), .ZN(n690) );
  NOR2_X1 U767 ( .A1(n834), .A2(n690), .ZN(n831) );
  NAND2_X1 U768 ( .A1(n831), .A2(G36), .ZN(G176) );
  NOR2_X1 U769 ( .A1(G164), .A2(G1384), .ZN(n793) );
  AND2_X1 U770 ( .A1(G40), .A2(n691), .ZN(n693) );
  NAND2_X1 U771 ( .A1(n693), .A2(n692), .ZN(n792) );
  INV_X1 U772 ( .A(n792), .ZN(n694) );
  NAND2_X1 U773 ( .A1(n793), .A2(n694), .ZN(n746) );
  INV_X1 U774 ( .A(G1996), .ZN(n695) );
  NOR2_X1 U775 ( .A1(n746), .A2(n695), .ZN(n697) );
  XOR2_X1 U776 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n696) );
  XNOR2_X1 U777 ( .A(n697), .B(n696), .ZN(n699) );
  NAND2_X1 U778 ( .A1(n746), .A2(G1341), .ZN(n698) );
  NAND2_X1 U779 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U780 ( .A1(n700), .A2(n966), .ZN(n706) );
  NAND2_X1 U781 ( .A1(n706), .A2(n976), .ZN(n704) );
  XNOR2_X1 U782 ( .A(n746), .B(KEYINPUT94), .ZN(n710) );
  INV_X1 U783 ( .A(n710), .ZN(n724) );
  NAND2_X1 U784 ( .A1(n724), .A2(G2067), .ZN(n702) );
  NAND2_X1 U785 ( .A1(G1348), .A2(n746), .ZN(n701) );
  NAND2_X1 U786 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U787 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U788 ( .A(KEYINPUT96), .B(n705), .Z(n708) );
  NOR2_X1 U789 ( .A1(n976), .A2(n706), .ZN(n707) );
  NOR2_X1 U790 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U791 ( .A(n709), .B(KEYINPUT97), .ZN(n716) );
  NAND2_X1 U792 ( .A1(n710), .A2(G1956), .ZN(n711) );
  XNOR2_X1 U793 ( .A(KEYINPUT95), .B(n711), .ZN(n714) );
  NAND2_X1 U794 ( .A1(G2072), .A2(n724), .ZN(n712) );
  XNOR2_X1 U795 ( .A(KEYINPUT27), .B(n712), .ZN(n713) );
  NOR2_X1 U796 ( .A1(n714), .A2(n713), .ZN(n718) );
  INV_X1 U797 ( .A(G299), .ZN(n717) );
  NAND2_X1 U798 ( .A1(n718), .A2(n717), .ZN(n715) );
  NAND2_X1 U799 ( .A1(n716), .A2(n715), .ZN(n721) );
  NOR2_X1 U800 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U801 ( .A(n719), .B(KEYINPUT28), .Z(n720) );
  NAND2_X1 U802 ( .A1(n721), .A2(n720), .ZN(n723) );
  XOR2_X1 U803 ( .A(KEYINPUT98), .B(KEYINPUT29), .Z(n722) );
  XNOR2_X1 U804 ( .A(n723), .B(n722), .ZN(n728) );
  XNOR2_X1 U805 ( .A(G2078), .B(KEYINPUT25), .ZN(n938) );
  NAND2_X1 U806 ( .A1(n724), .A2(n938), .ZN(n726) );
  INV_X1 U807 ( .A(G1961), .ZN(n1005) );
  NAND2_X1 U808 ( .A1(n1005), .A2(n746), .ZN(n725) );
  NAND2_X1 U809 ( .A1(n726), .A2(n725), .ZN(n732) );
  NAND2_X1 U810 ( .A1(n732), .A2(G171), .ZN(n727) );
  NAND2_X1 U811 ( .A1(n728), .A2(n727), .ZN(n737) );
  NOR2_X1 U812 ( .A1(G2084), .A2(n746), .ZN(n742) );
  NAND2_X1 U813 ( .A1(G8), .A2(n746), .ZN(n775) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n775), .ZN(n738) );
  NOR2_X1 U815 ( .A1(n742), .A2(n738), .ZN(n729) );
  NAND2_X1 U816 ( .A1(G8), .A2(n729), .ZN(n730) );
  XNOR2_X1 U817 ( .A(KEYINPUT30), .B(n730), .ZN(n731) );
  NOR2_X1 U818 ( .A1(G168), .A2(n731), .ZN(n734) );
  NOR2_X1 U819 ( .A1(G171), .A2(n732), .ZN(n733) );
  NOR2_X1 U820 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U821 ( .A(KEYINPUT31), .B(n735), .Z(n736) );
  NAND2_X1 U822 ( .A1(n737), .A2(n736), .ZN(n745) );
  INV_X1 U823 ( .A(n745), .ZN(n739) );
  NOR2_X1 U824 ( .A1(n739), .A2(n738), .ZN(n741) );
  XNOR2_X1 U825 ( .A(n741), .B(n740), .ZN(n744) );
  NAND2_X1 U826 ( .A1(G8), .A2(n742), .ZN(n743) );
  NAND2_X1 U827 ( .A1(n744), .A2(n743), .ZN(n755) );
  NAND2_X1 U828 ( .A1(G286), .A2(n745), .ZN(n751) );
  NOR2_X1 U829 ( .A1(G1971), .A2(n775), .ZN(n748) );
  NOR2_X1 U830 ( .A1(G2090), .A2(n746), .ZN(n747) );
  NOR2_X1 U831 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U832 ( .A1(G303), .A2(n749), .ZN(n750) );
  NAND2_X1 U833 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U834 ( .A1(G8), .A2(n752), .ZN(n753) );
  XNOR2_X1 U835 ( .A(n753), .B(KEYINPUT32), .ZN(n754) );
  NAND2_X1 U836 ( .A1(n755), .A2(n754), .ZN(n768) );
  NOR2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n761) );
  NOR2_X1 U838 ( .A1(G303), .A2(G1971), .ZN(n756) );
  NOR2_X1 U839 ( .A1(n761), .A2(n756), .ZN(n972) );
  NAND2_X1 U840 ( .A1(n768), .A2(n972), .ZN(n758) );
  NAND2_X1 U841 ( .A1(G288), .A2(G1976), .ZN(n757) );
  XNOR2_X1 U842 ( .A(n757), .B(KEYINPUT100), .ZN(n968) );
  NAND2_X1 U843 ( .A1(n758), .A2(n968), .ZN(n759) );
  NOR2_X1 U844 ( .A1(n759), .A2(n775), .ZN(n760) );
  NOR2_X1 U845 ( .A1(n760), .A2(KEYINPUT33), .ZN(n764) );
  NAND2_X1 U846 ( .A1(n761), .A2(KEYINPUT33), .ZN(n762) );
  NOR2_X1 U847 ( .A1(n775), .A2(n762), .ZN(n763) );
  NOR2_X1 U848 ( .A1(n764), .A2(n763), .ZN(n765) );
  XOR2_X1 U849 ( .A(G1981), .B(G305), .Z(n963) );
  NAND2_X1 U850 ( .A1(n765), .A2(n963), .ZN(n771) );
  NOR2_X1 U851 ( .A1(G303), .A2(G2090), .ZN(n766) );
  NAND2_X1 U852 ( .A1(G8), .A2(n766), .ZN(n767) );
  NAND2_X1 U853 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U854 ( .A1(n769), .A2(n775), .ZN(n770) );
  NAND2_X1 U855 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U856 ( .A(n772), .B(KEYINPUT101), .ZN(n814) );
  NOR2_X1 U857 ( .A1(G1981), .A2(G305), .ZN(n773) );
  XOR2_X1 U858 ( .A(n773), .B(KEYINPUT24), .Z(n774) );
  OR2_X1 U859 ( .A1(n775), .A2(n774), .ZN(n812) );
  NAND2_X1 U860 ( .A1(G141), .A2(n875), .ZN(n777) );
  NAND2_X1 U861 ( .A1(G129), .A2(n879), .ZN(n776) );
  NAND2_X1 U862 ( .A1(n777), .A2(n776), .ZN(n780) );
  NAND2_X1 U863 ( .A1(n876), .A2(G105), .ZN(n778) );
  XOR2_X1 U864 ( .A(KEYINPUT38), .B(n778), .Z(n779) );
  NOR2_X1 U865 ( .A1(n780), .A2(n779), .ZN(n782) );
  NAND2_X1 U866 ( .A1(n880), .A2(G117), .ZN(n781) );
  NAND2_X1 U867 ( .A1(n782), .A2(n781), .ZN(n890) );
  NOR2_X1 U868 ( .A1(G1996), .A2(n890), .ZN(n928) );
  NAND2_X1 U869 ( .A1(G119), .A2(n879), .ZN(n784) );
  NAND2_X1 U870 ( .A1(G107), .A2(n880), .ZN(n783) );
  NAND2_X1 U871 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U872 ( .A(KEYINPUT92), .B(n785), .Z(n789) );
  NAND2_X1 U873 ( .A1(G131), .A2(n875), .ZN(n787) );
  NAND2_X1 U874 ( .A1(G95), .A2(n876), .ZN(n786) );
  AND2_X1 U875 ( .A1(n787), .A2(n786), .ZN(n788) );
  NAND2_X1 U876 ( .A1(n789), .A2(n788), .ZN(n887) );
  XOR2_X1 U877 ( .A(KEYINPUT93), .B(G1991), .Z(n947) );
  AND2_X1 U878 ( .A1(n887), .A2(n947), .ZN(n791) );
  AND2_X1 U879 ( .A1(n890), .A2(G1996), .ZN(n790) );
  NOR2_X1 U880 ( .A1(n791), .A2(n790), .ZN(n914) );
  NOR2_X1 U881 ( .A1(n793), .A2(n792), .ZN(n820) );
  INV_X1 U882 ( .A(n820), .ZN(n794) );
  NOR2_X1 U883 ( .A1(n914), .A2(n794), .ZN(n816) );
  NOR2_X1 U884 ( .A1(n947), .A2(n887), .ZN(n916) );
  NOR2_X1 U885 ( .A1(G1986), .A2(G290), .ZN(n795) );
  NOR2_X1 U886 ( .A1(n916), .A2(n795), .ZN(n796) );
  NOR2_X1 U887 ( .A1(n816), .A2(n796), .ZN(n797) );
  NOR2_X1 U888 ( .A1(n928), .A2(n797), .ZN(n798) );
  XNOR2_X1 U889 ( .A(KEYINPUT39), .B(n798), .ZN(n808) );
  XNOR2_X1 U890 ( .A(G2067), .B(KEYINPUT37), .ZN(n809) );
  NAND2_X1 U891 ( .A1(G140), .A2(n875), .ZN(n800) );
  NAND2_X1 U892 ( .A1(G104), .A2(n876), .ZN(n799) );
  NAND2_X1 U893 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U894 ( .A(KEYINPUT34), .B(n801), .ZN(n806) );
  NAND2_X1 U895 ( .A1(G128), .A2(n879), .ZN(n803) );
  NAND2_X1 U896 ( .A1(G116), .A2(n880), .ZN(n802) );
  NAND2_X1 U897 ( .A1(n803), .A2(n802), .ZN(n804) );
  XOR2_X1 U898 ( .A(KEYINPUT35), .B(n804), .Z(n805) );
  NOR2_X1 U899 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U900 ( .A(KEYINPUT36), .B(n807), .ZN(n872) );
  NOR2_X1 U901 ( .A1(n809), .A2(n872), .ZN(n921) );
  NAND2_X1 U902 ( .A1(n820), .A2(n921), .ZN(n818) );
  NAND2_X1 U903 ( .A1(n808), .A2(n818), .ZN(n810) );
  NAND2_X1 U904 ( .A1(n809), .A2(n872), .ZN(n913) );
  NAND2_X1 U905 ( .A1(n810), .A2(n913), .ZN(n811) );
  NAND2_X1 U906 ( .A1(n811), .A2(n820), .ZN(n815) );
  AND2_X1 U907 ( .A1(n812), .A2(n815), .ZN(n813) );
  NAND2_X1 U908 ( .A1(n814), .A2(n813), .ZN(n826) );
  INV_X1 U909 ( .A(n815), .ZN(n824) );
  INV_X1 U910 ( .A(n816), .ZN(n817) );
  NAND2_X1 U911 ( .A1(n818), .A2(n817), .ZN(n822) );
  XOR2_X1 U912 ( .A(G1986), .B(KEYINPUT91), .Z(n819) );
  XNOR2_X1 U913 ( .A(G290), .B(n819), .ZN(n974) );
  AND2_X1 U914 ( .A1(n974), .A2(n820), .ZN(n821) );
  NOR2_X1 U915 ( .A1(n822), .A2(n821), .ZN(n823) );
  OR2_X1 U916 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U917 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U918 ( .A(n827), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n828), .ZN(G217) );
  AND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U921 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U923 ( .A1(n831), .A2(n830), .ZN(G188) );
  XNOR2_X1 U924 ( .A(G96), .B(KEYINPUT105), .ZN(G221) );
  INV_X1 U926 ( .A(G132), .ZN(G219) );
  INV_X1 U927 ( .A(G120), .ZN(G236) );
  INV_X1 U928 ( .A(G82), .ZN(G220) );
  INV_X1 U929 ( .A(G69), .ZN(G235) );
  NOR2_X1 U930 ( .A1(n833), .A2(n832), .ZN(G325) );
  INV_X1 U931 ( .A(G325), .ZN(G261) );
  INV_X1 U932 ( .A(n834), .ZN(G319) );
  XOR2_X1 U933 ( .A(KEYINPUT107), .B(G2678), .Z(n836) );
  XNOR2_X1 U934 ( .A(KEYINPUT43), .B(G2096), .ZN(n835) );
  XNOR2_X1 U935 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U936 ( .A(n837), .B(KEYINPUT42), .Z(n839) );
  XNOR2_X1 U937 ( .A(G2067), .B(G2084), .ZN(n838) );
  XNOR2_X1 U938 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U939 ( .A(G2100), .B(G2072), .Z(n841) );
  XNOR2_X1 U940 ( .A(G2090), .B(G2078), .ZN(n840) );
  XNOR2_X1 U941 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U942 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U943 ( .A(KEYINPUT106), .B(KEYINPUT108), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(G227) );
  XOR2_X1 U945 ( .A(G1956), .B(G1961), .Z(n847) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1981), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U948 ( .A(G1976), .B(G1971), .Z(n849) );
  XNOR2_X1 U949 ( .A(G1996), .B(G1991), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U951 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U952 ( .A(KEYINPUT109), .B(G2474), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(n855) );
  XOR2_X1 U954 ( .A(G1966), .B(KEYINPUT41), .Z(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(G229) );
  NAND2_X1 U956 ( .A1(n880), .A2(G112), .ZN(n862) );
  NAND2_X1 U957 ( .A1(G136), .A2(n875), .ZN(n857) );
  NAND2_X1 U958 ( .A1(G100), .A2(n876), .ZN(n856) );
  NAND2_X1 U959 ( .A1(n857), .A2(n856), .ZN(n860) );
  NAND2_X1 U960 ( .A1(n879), .A2(G124), .ZN(n858) );
  XOR2_X1 U961 ( .A(KEYINPUT44), .B(n858), .Z(n859) );
  NOR2_X1 U962 ( .A1(n860), .A2(n859), .ZN(n861) );
  NAND2_X1 U963 ( .A1(n862), .A2(n861), .ZN(n863) );
  XOR2_X1 U964 ( .A(KEYINPUT110), .B(n863), .Z(G162) );
  NAND2_X1 U965 ( .A1(G130), .A2(n879), .ZN(n865) );
  NAND2_X1 U966 ( .A1(G118), .A2(n880), .ZN(n864) );
  NAND2_X1 U967 ( .A1(n865), .A2(n864), .ZN(n871) );
  NAND2_X1 U968 ( .A1(G142), .A2(n875), .ZN(n867) );
  NAND2_X1 U969 ( .A1(G106), .A2(n876), .ZN(n866) );
  NAND2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U971 ( .A(KEYINPUT111), .B(n868), .ZN(n869) );
  XNOR2_X1 U972 ( .A(KEYINPUT45), .B(n869), .ZN(n870) );
  NOR2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U975 ( .A(n874), .B(G162), .ZN(n886) );
  NAND2_X1 U976 ( .A1(G139), .A2(n875), .ZN(n878) );
  NAND2_X1 U977 ( .A1(G103), .A2(n876), .ZN(n877) );
  NAND2_X1 U978 ( .A1(n878), .A2(n877), .ZN(n885) );
  NAND2_X1 U979 ( .A1(G127), .A2(n879), .ZN(n882) );
  NAND2_X1 U980 ( .A1(G115), .A2(n880), .ZN(n881) );
  NAND2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U982 ( .A(KEYINPUT47), .B(n883), .Z(n884) );
  NOR2_X1 U983 ( .A1(n885), .A2(n884), .ZN(n909) );
  XOR2_X1 U984 ( .A(n886), .B(n909), .Z(n889) );
  XOR2_X1 U985 ( .A(G164), .B(n887), .Z(n888) );
  XNOR2_X1 U986 ( .A(n889), .B(n888), .ZN(n895) );
  XOR2_X1 U987 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n892) );
  XOR2_X1 U988 ( .A(n890), .B(n915), .Z(n891) );
  XNOR2_X1 U989 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U990 ( .A(G160), .B(n893), .ZN(n894) );
  XNOR2_X1 U991 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U992 ( .A1(G37), .A2(n896), .ZN(G395) );
  XNOR2_X1 U993 ( .A(n966), .B(n897), .ZN(n899) );
  XNOR2_X1 U994 ( .A(G171), .B(n976), .ZN(n898) );
  XNOR2_X1 U995 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U996 ( .A(G286), .B(n900), .ZN(n901) );
  NOR2_X1 U997 ( .A1(G37), .A2(n901), .ZN(G397) );
  NOR2_X1 U998 ( .A1(G227), .A2(G229), .ZN(n902) );
  XOR2_X1 U999 ( .A(KEYINPUT49), .B(n902), .Z(n903) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n903), .ZN(n904) );
  NOR2_X1 U1001 ( .A1(G401), .A2(n904), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(KEYINPUT112), .B(n905), .ZN(n907) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n906) );
  NAND2_X1 U1004 ( .A1(n907), .A2(n906), .ZN(n908) );
  XOR2_X1 U1005 ( .A(KEYINPUT113), .B(n908), .Z(G225) );
  INV_X1 U1006 ( .A(G225), .ZN(G308) );
  INV_X1 U1007 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1008 ( .A(G2072), .B(n909), .Z(n911) );
  XOR2_X1 U1009 ( .A(G164), .B(G2078), .Z(n910) );
  NOR2_X1 U1010 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(KEYINPUT50), .B(n912), .ZN(n926) );
  NAND2_X1 U1012 ( .A1(n914), .A2(n913), .ZN(n924) );
  NOR2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(KEYINPUT114), .B(n917), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(G160), .B(G2084), .ZN(n918) );
  NAND2_X1 U1016 ( .A1(n919), .A2(n918), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(KEYINPUT115), .B(n922), .ZN(n923) );
  NOR2_X1 U1019 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1020 ( .A1(n926), .A2(n925), .ZN(n932) );
  XOR2_X1 U1021 ( .A(G2090), .B(G162), .Z(n927) );
  NOR2_X1 U1022 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1023 ( .A(KEYINPUT116), .B(n929), .ZN(n930) );
  XNOR2_X1 U1024 ( .A(KEYINPUT51), .B(n930), .ZN(n931) );
  NOR2_X1 U1025 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1026 ( .A(n933), .B(KEYINPUT52), .Z(n934) );
  XNOR2_X1 U1027 ( .A(KEYINPUT117), .B(n934), .ZN(n935) );
  INV_X1 U1028 ( .A(KEYINPUT55), .ZN(n957) );
  NAND2_X1 U1029 ( .A1(n935), .A2(n957), .ZN(n936) );
  NAND2_X1 U1030 ( .A1(n936), .A2(G29), .ZN(n1020) );
  XNOR2_X1 U1031 ( .A(G2090), .B(G35), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(n937), .B(KEYINPUT118), .ZN(n952) );
  XNOR2_X1 U1033 ( .A(G27), .B(n938), .ZN(n946) );
  XNOR2_X1 U1034 ( .A(G2067), .B(G26), .ZN(n940) );
  XNOR2_X1 U1035 ( .A(G33), .B(G2072), .ZN(n939) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1037 ( .A1(G28), .A2(n941), .ZN(n944) );
  XOR2_X1 U1038 ( .A(G32), .B(G1996), .Z(n942) );
  XNOR2_X1 U1039 ( .A(KEYINPUT119), .B(n942), .ZN(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(G25), .B(n947), .ZN(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(n950), .B(KEYINPUT53), .ZN(n951) );
  NOR2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n955) );
  XOR2_X1 U1046 ( .A(G2084), .B(G34), .Z(n953) );
  XNOR2_X1 U1047 ( .A(KEYINPUT54), .B(n953), .ZN(n954) );
  NAND2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(n957), .B(n956), .ZN(n959) );
  INV_X1 U1050 ( .A(G29), .ZN(n958) );
  NAND2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1052 ( .A1(G11), .A2(n960), .ZN(n1018) );
  XNOR2_X1 U1053 ( .A(G16), .B(KEYINPUT56), .ZN(n987) );
  XNOR2_X1 U1054 ( .A(G1966), .B(G168), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(n961), .B(KEYINPUT120), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n965) );
  XOR2_X1 U1057 ( .A(KEYINPUT121), .B(KEYINPUT57), .Z(n964) );
  XNOR2_X1 U1058 ( .A(n965), .B(n964), .ZN(n985) );
  XNOR2_X1 U1059 ( .A(n966), .B(G1341), .ZN(n983) );
  NAND2_X1 U1060 ( .A1(G303), .A2(G1971), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(G1956), .B(G299), .ZN(n969) );
  NOR2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1066 ( .A(KEYINPUT122), .B(n975), .ZN(n978) );
  XNOR2_X1 U1067 ( .A(n976), .B(G1348), .ZN(n977) );
  NAND2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n980) );
  XOR2_X1 U1069 ( .A(G171), .B(G1961), .Z(n979) );
  NOR2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1071 ( .A(KEYINPUT123), .B(n981), .ZN(n982) );
  NOR2_X1 U1072 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1073 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1074 ( .A1(n987), .A2(n986), .ZN(n1016) );
  INV_X1 U1075 ( .A(G16), .ZN(n1014) );
  XNOR2_X1 U1076 ( .A(KEYINPUT61), .B(KEYINPUT127), .ZN(n1012) );
  XNOR2_X1 U1077 ( .A(G1971), .B(G22), .ZN(n989) );
  XNOR2_X1 U1078 ( .A(G23), .B(G1976), .ZN(n988) );
  NOR2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n991) );
  XOR2_X1 U1080 ( .A(G1986), .B(G24), .Z(n990) );
  NAND2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n993) );
  XOR2_X1 U1082 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n992) );
  XNOR2_X1 U1083 ( .A(n993), .B(n992), .ZN(n1010) );
  XOR2_X1 U1084 ( .A(G1966), .B(G21), .Z(n1004) );
  XOR2_X1 U1085 ( .A(G1348), .B(KEYINPUT59), .Z(n994) );
  XNOR2_X1 U1086 ( .A(G4), .B(n994), .ZN(n1001) );
  XOR2_X1 U1087 ( .A(G1341), .B(G19), .Z(n998) );
  XNOR2_X1 U1088 ( .A(G1981), .B(G6), .ZN(n996) );
  XNOR2_X1 U1089 ( .A(G20), .B(G1956), .ZN(n995) );
  NOR2_X1 U1090 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1091 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1092 ( .A(KEYINPUT125), .B(n999), .Z(n1000) );
  NOR2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1094 ( .A(KEYINPUT60), .B(n1002), .ZN(n1003) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1008) );
  XOR2_X1 U1096 ( .A(KEYINPUT124), .B(n1005), .Z(n1006) );
  XNOR2_X1 U1097 ( .A(G5), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(n1012), .B(n1011), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1021), .Z(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
endmodule

