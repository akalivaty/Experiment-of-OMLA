//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 1 0 0 1 0 1 1 1 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1 1 0 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 1 0 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n231, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1263, new_n1264, new_n1265, new_n1267,
    new_n1268, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n205), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT1), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n202), .A2(G50), .ZN(new_n214));
  NAND3_X1  g0014(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT0), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n205), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n216), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n220), .B1(new_n217), .B2(new_n219), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n213), .A2(new_n221), .ZN(G361));
  XNOR2_X1  g0022(.A(G238), .B(G244), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(G232), .ZN(new_n224));
  XOR2_X1   g0024(.A(KEYINPUT2), .B(G226), .Z(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(G250), .B(G257), .Z(new_n227));
  XNOR2_X1  g0027(.A(G264), .B(G270), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n226), .B(new_n229), .Z(G358));
  XNOR2_X1  g0030(.A(G50), .B(G68), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G58), .B(G77), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n231), .B(new_n232), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT64), .ZN(new_n234));
  INV_X1    g0034(.A(G107), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n235), .A2(G97), .ZN(new_n236));
  INV_X1    g0036(.A(G97), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n237), .A2(G107), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G87), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n234), .B(new_n241), .ZN(G351));
  INV_X1    g0042(.A(KEYINPUT13), .ZN(new_n243));
  INV_X1    g0043(.A(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(KEYINPUT3), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT3), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  NAND4_X1  g0048(.A1(new_n245), .A2(new_n247), .A3(G226), .A4(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT72), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT3), .B(G33), .ZN(new_n252));
  NAND4_X1  g0052(.A1(new_n252), .A2(KEYINPUT72), .A3(G226), .A4(new_n248), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G97), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n252), .A2(G232), .A3(G1698), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n251), .A2(new_n253), .A3(new_n254), .A4(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G1), .A3(G13), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  INV_X1    g0061(.A(G45), .ZN(new_n262));
  AOI21_X1  g0062(.A(G1), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G274), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n258), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G238), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n264), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n243), .B1(new_n260), .B2(new_n270), .ZN(new_n271));
  AOI211_X1 g0071(.A(KEYINPUT13), .B(new_n269), .C1(new_n256), .C2(new_n259), .ZN(new_n272));
  OAI21_X1  g0072(.A(G169), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT14), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n260), .A2(new_n270), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT13), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n260), .A2(new_n243), .A3(new_n270), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(G179), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT14), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n279), .B(G169), .C1(new_n271), .C2(new_n272), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n274), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G1), .A2(G13), .ZN(new_n283));
  AND2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G20), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n244), .ZN(new_n287));
  INV_X1    g0087(.A(G50), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT74), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G77), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n286), .A2(G33), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n289), .B1(new_n286), .B2(G68), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  NOR3_X1   g0092(.A1(new_n287), .A2(KEYINPUT74), .A3(new_n288), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n285), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT11), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n265), .A2(G13), .A3(G20), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G68), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n297), .A2(KEYINPUT12), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT12), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(new_n296), .B2(G68), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n282), .B(new_n283), .C1(G1), .C2(new_n286), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n299), .B(new_n301), .C1(new_n302), .C2(new_n298), .ZN(new_n303));
  XOR2_X1   g0103(.A(new_n303), .B(KEYINPUT75), .Z(new_n304));
  AND2_X1   g0104(.A1(new_n295), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n281), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n276), .A2(new_n277), .ZN(new_n308));
  INV_X1    g0108(.A(G190), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT73), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT73), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n276), .A2(new_n311), .A3(G190), .A4(new_n277), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n308), .A2(G200), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n310), .A2(new_n305), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n307), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n316), .B(KEYINPUT76), .ZN(new_n317));
  OAI21_X1  g0117(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n318));
  INV_X1    g0118(.A(G150), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n318), .B1(new_n319), .B2(new_n287), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT66), .B(G58), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT8), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT67), .ZN(new_n323));
  INV_X1    g0123(.A(G58), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(KEYINPUT8), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT8), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(KEYINPUT67), .A3(G58), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n322), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n291), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n320), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(new_n284), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n297), .A2(new_n288), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n288), .B2(new_n302), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  OR3_X1    g0134(.A1(new_n334), .A2(KEYINPUT70), .A3(KEYINPUT9), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT70), .B1(new_n334), .B2(KEYINPUT9), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n252), .A2(G222), .A3(new_n248), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n252), .A2(G1698), .ZN(new_n339));
  INV_X1    g0139(.A(G223), .ZN(new_n340));
  OAI221_X1 g0140(.A(new_n338), .B1(new_n290), .B2(new_n252), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n259), .ZN(new_n342));
  INV_X1    g0142(.A(new_n264), .ZN(new_n343));
  INV_X1    g0143(.A(new_n267), .ZN(new_n344));
  XNOR2_X1  g0144(.A(KEYINPUT65), .B(G226), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n347), .A2(new_n309), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(G200), .B2(new_n347), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT9), .ZN(new_n350));
  NOR4_X1   g0150(.A1(new_n331), .A2(KEYINPUT71), .A3(new_n350), .A4(new_n333), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT71), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(new_n334), .B2(KEYINPUT9), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n349), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT10), .B1(new_n337), .B2(new_n354), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n353), .A2(new_n351), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n335), .A2(new_n336), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT10), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n356), .A2(new_n357), .A3(new_n358), .A4(new_n349), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT16), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT78), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(new_n244), .B2(KEYINPUT3), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n246), .A2(KEYINPUT78), .A3(G33), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n363), .A2(new_n245), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT7), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n366), .A2(G20), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n366), .B1(new_n252), .B2(G20), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n298), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G159), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT77), .B1(new_n287), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(G20), .A2(G33), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT77), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(new_n374), .A3(G159), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  AND2_X1   g0176(.A1(KEYINPUT66), .A2(G58), .ZN(new_n377));
  NOR2_X1   g0177(.A1(KEYINPUT66), .A2(G58), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n201), .B1(new_n379), .B2(G68), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n376), .B1(new_n380), .B2(new_n286), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n361), .B1(new_n370), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n245), .A2(new_n247), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT7), .B1(new_n383), .B2(new_n286), .ZN(new_n384));
  AOI211_X1 g0184(.A(new_n366), .B(G20), .C1(new_n245), .C2(new_n247), .ZN(new_n385));
  OAI21_X1  g0185(.A(G68), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n202), .B1(new_n321), .B2(new_n298), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n387), .A2(G20), .B1(new_n372), .B2(new_n375), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n388), .A3(KEYINPUT16), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n382), .A2(new_n285), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT79), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n322), .A2(new_n296), .A3(new_n325), .A4(new_n327), .ZN(new_n392));
  INV_X1    g0192(.A(new_n378), .ZN(new_n393));
  NAND2_X1  g0193(.A1(KEYINPUT66), .A2(G58), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n326), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n325), .A2(new_n327), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n302), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n391), .B1(new_n392), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n392), .A2(new_n397), .A3(new_n391), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n390), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n245), .A2(new_n247), .A3(G226), .A4(G1698), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n245), .A2(new_n247), .A3(G223), .A4(new_n248), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G87), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n259), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n258), .A2(G232), .A3(new_n266), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n264), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G169), .ZN(new_n412));
  OR2_X1    g0212(.A1(KEYINPUT68), .A2(G179), .ZN(new_n413));
  NAND2_X1  g0213(.A1(KEYINPUT68), .A2(G179), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n407), .A2(new_n410), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT80), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n412), .A2(KEYINPUT80), .A3(new_n416), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n402), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT18), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI211_X1 g0223(.A(new_n309), .B(new_n409), .C1(new_n259), .C2(new_n406), .ZN(new_n424));
  INV_X1    g0224(.A(G200), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n407), .B2(new_n410), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n390), .A2(new_n427), .A3(new_n401), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT17), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n390), .A2(new_n427), .A3(new_n401), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT17), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n402), .A2(new_n419), .A3(new_n420), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT18), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n423), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n347), .A2(new_n415), .ZN(new_n438));
  INV_X1    g0238(.A(G169), .ZN(new_n439));
  AOI211_X1 g0239(.A(new_n334), .B(new_n438), .C1(new_n439), .C2(new_n347), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  XNOR2_X1  g0241(.A(KEYINPUT8), .B(G58), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n443), .A2(new_n373), .B1(G20), .B2(G77), .ZN(new_n444));
  XOR2_X1   g0244(.A(KEYINPUT15), .B(G87), .Z(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n329), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n284), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n297), .A2(new_n290), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(new_n290), .B2(new_n302), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n252), .A2(G232), .A3(new_n248), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n383), .A2(G107), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n451), .B(new_n452), .C1(new_n339), .C2(new_n268), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n259), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT69), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n343), .B1(new_n344), .B2(G244), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n455), .B1(new_n454), .B2(new_n456), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n450), .B1(new_n459), .B2(new_n439), .ZN(new_n460));
  INV_X1    g0260(.A(new_n415), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(new_n457), .B2(new_n458), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n459), .A2(G200), .ZN(new_n465));
  OAI21_X1  g0265(.A(G190), .B1(new_n457), .B2(new_n458), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n465), .A2(new_n466), .A3(new_n450), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n360), .A2(new_n437), .A3(new_n441), .A4(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n317), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(G116), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n282), .A2(new_n283), .B1(G20), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G283), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n474), .B(new_n286), .C1(G33), .C2(new_n237), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n473), .A2(KEYINPUT20), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT86), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n473), .A2(new_n475), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT20), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT86), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n473), .A2(new_n481), .A3(new_n475), .A4(KEYINPUT20), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n477), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n296), .A2(G116), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n265), .A2(G33), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n284), .A2(new_n296), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n484), .B1(new_n486), .B2(G116), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT87), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n245), .A2(new_n247), .A3(G257), .A4(new_n248), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n245), .A2(new_n247), .A3(G264), .A4(G1698), .ZN(new_n491));
  INV_X1    g0291(.A(G303), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n490), .B(new_n491), .C1(new_n492), .C2(new_n252), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n259), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n262), .A2(G1), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n495), .B(KEYINPUT83), .C1(KEYINPUT5), .C2(new_n261), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n265), .B(G45), .C1(new_n261), .C2(KEYINPUT5), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT83), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(G274), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n500), .B1(KEYINPUT5), .B2(new_n261), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n496), .A2(new_n499), .A3(new_n258), .A4(new_n501), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n261), .A2(KEYINPUT5), .ZN(new_n503));
  OAI211_X1 g0303(.A(G270), .B(new_n258), .C1(new_n497), .C2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n494), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G200), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT87), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n483), .A2(new_n487), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n489), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT88), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n489), .A2(new_n506), .A3(KEYINPUT88), .A4(new_n508), .ZN(new_n512));
  OR2_X1    g0312(.A1(new_n505), .A2(new_n309), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n505), .A2(G169), .ZN(new_n515));
  INV_X1    g0315(.A(new_n508), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n507), .B1(new_n483), .B2(new_n487), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT21), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n489), .A2(new_n508), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n521), .A2(KEYINPUT21), .A3(new_n515), .ZN(new_n522));
  INV_X1    g0322(.A(G179), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n505), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n520), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n514), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(G87), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(KEYINPUT89), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n529), .A2(new_n245), .A3(new_n247), .A4(new_n286), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT22), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n252), .A2(KEYINPUT22), .A3(new_n286), .A4(new_n529), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G116), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n534), .A2(G20), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT23), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n286), .B2(G107), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n235), .A2(KEYINPUT23), .A3(G20), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n532), .A2(new_n533), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT24), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n284), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n532), .A2(new_n533), .A3(new_n539), .A4(KEYINPUT24), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n245), .A2(new_n247), .A3(G250), .A4(new_n248), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n245), .A2(new_n247), .A3(G257), .A4(G1698), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G294), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n548), .A2(new_n259), .ZN(new_n549));
  OAI211_X1 g0349(.A(G264), .B(new_n258), .C1(new_n497), .C2(new_n503), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n502), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(G200), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n297), .A2(KEYINPUT25), .A3(new_n235), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT25), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n296), .B2(G107), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n284), .A2(new_n296), .A3(new_n485), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n556), .B1(new_n235), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n548), .A2(new_n259), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n560), .A2(G190), .A3(new_n502), .A4(new_n550), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n544), .A2(new_n552), .A3(new_n559), .A4(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n558), .B1(new_n542), .B2(new_n543), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n560), .A2(new_n502), .A3(new_n550), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n439), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n560), .A2(new_n523), .A3(new_n502), .A4(new_n550), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n562), .B1(new_n563), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n252), .A2(G238), .A3(new_n248), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n245), .A2(new_n247), .A3(G244), .A4(G1698), .ZN(new_n570));
  AND3_X1   g0370(.A1(new_n569), .A2(new_n534), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(G250), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n265), .B2(G45), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n258), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n495), .A2(G274), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n574), .A2(KEYINPUT85), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT85), .B1(new_n574), .B2(new_n575), .ZN(new_n577));
  OAI22_X1  g0377(.A1(new_n571), .A2(new_n258), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G200), .ZN(new_n579));
  INV_X1    g0379(.A(new_n577), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n573), .A2(new_n258), .B1(new_n495), .B2(G274), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT85), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n569), .A2(new_n534), .A3(new_n570), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n580), .A2(new_n582), .B1(new_n583), .B2(new_n259), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(G190), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n445), .A2(new_n296), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n252), .A2(new_n286), .A3(G68), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT19), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n286), .B1(new_n254), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n528), .A2(new_n237), .A3(new_n235), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n588), .B1(new_n291), .B2(new_n237), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n587), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n586), .B1(new_n593), .B2(new_n285), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n486), .A2(G87), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n579), .A2(new_n585), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n580), .A2(new_n582), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n583), .A2(new_n259), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(new_n461), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n486), .A2(new_n445), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n594), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n600), .B(new_n602), .C1(G169), .C2(new_n584), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n568), .A2(new_n604), .ZN(new_n605));
  OAI211_X1 g0405(.A(G257), .B(new_n258), .C1(new_n497), .C2(new_n503), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n245), .A2(new_n247), .A3(G244), .A4(new_n248), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT82), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT4), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n609), .B1(new_n607), .B2(new_n608), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n245), .A2(new_n247), .A3(G250), .A4(G1698), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n474), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n502), .B(new_n606), .C1(new_n614), .C2(new_n258), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G200), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n297), .A2(KEYINPUT81), .A3(new_n237), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT81), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(new_n296), .B2(G97), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(new_n237), .B2(new_n557), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT6), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n236), .A2(new_n238), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n235), .A2(KEYINPUT6), .A3(G97), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n625), .A2(G20), .B1(G77), .B2(new_n373), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n383), .A2(new_n286), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n627), .A2(new_n366), .B1(new_n365), .B2(new_n367), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n626), .B1(new_n628), .B2(new_n235), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n621), .B1(new_n629), .B2(new_n285), .ZN(new_n630));
  INV_X1    g0430(.A(new_n606), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n607), .A2(new_n608), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT4), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n634));
  INV_X1    g0434(.A(new_n613), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n631), .B1(new_n636), .B2(new_n259), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n637), .A2(G190), .A3(new_n502), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n616), .A2(new_n630), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n636), .A2(new_n259), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n641), .A2(new_n461), .A3(new_n502), .A4(new_n606), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n629), .A2(new_n285), .ZN(new_n643));
  INV_X1    g0443(.A(new_n621), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n502), .ZN(new_n646));
  AOI211_X1 g0446(.A(new_n646), .B(new_n631), .C1(new_n636), .C2(new_n259), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n642), .B(new_n645), .C1(new_n647), .C2(G169), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT84), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n630), .B1(new_n439), .B2(new_n615), .ZN(new_n651));
  AOI21_X1  g0451(.A(KEYINPUT84), .B1(new_n651), .B2(new_n642), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n605), .B(new_n640), .C1(new_n650), .C2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n471), .A2(new_n527), .A3(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(G372));
  AOI22_X1  g0456(.A1(new_n390), .A2(new_n401), .B1(new_n412), .B2(new_n416), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n657), .B(KEYINPUT18), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n307), .A2(new_n464), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n314), .A2(new_n433), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n440), .B1(new_n661), .B2(new_n360), .ZN(new_n662));
  INV_X1    g0462(.A(new_n471), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n648), .A2(new_n649), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n651), .A2(KEYINPUT84), .A3(new_n642), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n664), .A2(new_n665), .A3(new_n603), .A4(new_n597), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(KEYINPUT26), .ZN(new_n667));
  INV_X1    g0467(.A(new_n603), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n594), .A2(new_n595), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT90), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n594), .A2(KEYINPUT90), .A3(new_n595), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n671), .A2(new_n579), .A3(new_n585), .A4(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n651), .A2(new_n673), .A3(new_n642), .A4(new_n603), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT26), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n668), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n639), .B1(new_n664), .B2(new_n665), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n673), .A2(new_n562), .A3(new_n603), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n567), .A2(new_n563), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT91), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n526), .ZN(new_n683));
  OAI211_X1 g0483(.A(new_n667), .B(new_n677), .C1(new_n680), .C2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n662), .B1(new_n663), .B2(new_n685), .ZN(G369));
  AND2_X1   g0486(.A1(new_n286), .A2(G13), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n265), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G213), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(G343), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n521), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n527), .A2(new_n694), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n520), .A2(new_n522), .A3(new_n525), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n695), .B1(new_n696), .B2(new_n694), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n567), .A2(new_n563), .ZN(new_n700));
  INV_X1    g0500(.A(new_n693), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n700), .B(new_n562), .C1(new_n563), .C2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n681), .A2(new_n693), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT92), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n702), .A2(KEYINPUT92), .A3(new_n703), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n699), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n526), .A2(new_n701), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n682), .A2(new_n701), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n709), .A2(new_n715), .ZN(G399));
  INV_X1    g0516(.A(new_n218), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(G41), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n590), .A2(G116), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(G1), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(new_n214), .B2(new_n719), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT28), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n520), .A2(new_n522), .A3(new_n525), .A4(new_n700), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n678), .A2(new_n679), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n668), .B1(new_n674), .B2(KEYINPUT26), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n666), .B2(KEYINPUT26), .ZN(new_n727));
  OAI211_X1 g0527(.A(KEYINPUT29), .B(new_n701), .C1(new_n725), .C2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n685), .A2(new_n693), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n728), .B1(new_n729), .B2(KEYINPUT29), .ZN(new_n730));
  INV_X1    g0530(.A(G330), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n578), .A2(new_n564), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(new_n524), .A3(new_n637), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT30), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n505), .A2(new_n461), .A3(new_n564), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n578), .A2(KEYINPUT93), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT93), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n584), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n736), .A2(new_n615), .A3(new_n737), .A4(new_n739), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n732), .A2(new_n524), .A3(KEYINPUT30), .A4(new_n637), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n735), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n693), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT31), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n742), .A2(KEYINPUT31), .A3(new_n693), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n527), .A2(new_n678), .A3(new_n605), .A4(new_n701), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n747), .B1(new_n748), .B2(KEYINPUT94), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT94), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n654), .A2(new_n750), .A3(new_n527), .A4(new_n701), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n731), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AND2_X1   g0553(.A1(new_n730), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n723), .B1(new_n754), .B2(G1), .ZN(G364));
  AOI21_X1  g0555(.A(new_n265), .B1(new_n687), .B2(G45), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n718), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G13), .A2(G33), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n697), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n283), .B1(G20), .B2(new_n439), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n233), .A2(new_n262), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n717), .A2(new_n252), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n214), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n770), .B1(new_n262), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n717), .A2(new_n383), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n773), .A2(G355), .B1(new_n472), .B2(new_n717), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n768), .A2(new_n772), .B1(KEYINPUT95), .B2(new_n775), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n775), .A2(KEYINPUT95), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n767), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n286), .A2(new_n309), .A3(G200), .ZN(new_n779));
  AND2_X1   g0579(.A1(new_n415), .A2(new_n779), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n309), .A2(G179), .A3(G200), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n286), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n780), .A2(new_n379), .B1(G97), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n286), .A2(G190), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n785), .A2(new_n523), .A3(G200), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n784), .B1(new_n235), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT32), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n785), .A2(new_n523), .A3(new_n425), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n788), .B1(new_n789), .B2(new_n371), .ZN(new_n790));
  INV_X1    g0590(.A(new_n789), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n791), .A2(KEYINPUT32), .A3(G159), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n787), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n286), .A2(new_n309), .A3(new_n425), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n523), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n415), .A2(new_n425), .A3(new_n785), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n252), .B1(new_n528), .B2(new_n795), .C1(new_n796), .C2(new_n290), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n415), .A2(G200), .A3(new_n785), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n797), .B1(G68), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT96), .ZN(new_n801));
  AND3_X1   g0601(.A1(new_n415), .A2(new_n801), .A3(new_n794), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n801), .B1(new_n415), .B2(new_n794), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n793), .B(new_n800), .C1(new_n288), .C2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT97), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G294), .ZN(new_n809));
  INV_X1    g0609(.A(G329), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n782), .A2(new_n809), .B1(new_n789), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G283), .ZN(new_n812));
  INV_X1    g0612(.A(G311), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n383), .B1(new_n812), .B2(new_n786), .C1(new_n796), .C2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n795), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n811), .B(new_n814), .C1(G303), .C2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n780), .A2(G322), .ZN(new_n817));
  XOR2_X1   g0617(.A(KEYINPUT33), .B(G317), .Z(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n798), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT98), .ZN(new_n820));
  INV_X1    g0620(.A(G326), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n816), .B(new_n820), .C1(new_n821), .C2(new_n805), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n806), .A2(new_n807), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n808), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n778), .B1(new_n824), .B2(new_n765), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n759), .B1(new_n764), .B2(new_n825), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n697), .A2(G330), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n758), .B1(new_n827), .B2(new_n698), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT99), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(G396));
  NOR2_X1   g0631(.A1(new_n765), .A2(new_n760), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n759), .B1(new_n290), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n765), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n252), .B1(new_n783), .B2(G97), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n835), .B1(new_n472), .B2(new_n796), .C1(new_n812), .C2(new_n798), .ZN(new_n836));
  INV_X1    g0636(.A(new_n786), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n815), .A2(G107), .B1(G87), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n780), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n838), .B1(new_n813), .B2(new_n789), .C1(new_n809), .C2(new_n839), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n836), .B(new_n840), .C1(G303), .C2(new_n804), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n383), .B1(new_n791), .B2(G132), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n843), .A2(KEYINPUT100), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n815), .A2(G50), .B1(G68), .B2(new_n837), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n845), .B1(new_n321), .B2(new_n782), .C1(new_n843), .C2(KEYINPUT100), .ZN(new_n846));
  INV_X1    g0646(.A(new_n796), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n847), .A2(G159), .B1(new_n780), .B2(G143), .ZN(new_n848));
  INV_X1    g0648(.A(G137), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n848), .B1(new_n319), .B2(new_n798), .C1(new_n805), .C2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT34), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n844), .B(new_n846), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  OR2_X1    g0652(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n841), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n450), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n693), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT101), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(new_n460), .B2(new_n462), .ZN(new_n858));
  INV_X1    g0658(.A(new_n458), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n859), .A2(new_n439), .A3(new_n860), .ZN(new_n861));
  AND4_X1   g0661(.A1(new_n857), .A2(new_n861), .A3(new_n462), .A4(new_n855), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n467), .B(new_n856), .C1(new_n858), .C2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n464), .A2(new_n693), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n833), .B1(new_n834), .B2(new_n854), .C1(new_n865), .C2(new_n761), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n858), .A2(new_n862), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n867), .A2(new_n468), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n684), .A2(new_n701), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n729), .B2(new_n865), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n758), .B1(new_n870), .B2(new_n753), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n870), .A2(new_n753), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n866), .B1(new_n872), .B2(new_n873), .ZN(G384));
  NAND3_X1  g0674(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n678), .A2(new_n696), .A3(new_n875), .A4(new_n605), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT94), .B1(new_n876), .B2(new_n693), .ZN(new_n877));
  INV_X1    g0677(.A(new_n747), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n877), .A2(new_n751), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n471), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n880), .B(KEYINPUT105), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n281), .A2(new_n306), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n306), .A2(new_n693), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n882), .A2(new_n314), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n281), .A2(new_n306), .A3(new_n693), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n865), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n749), .B2(new_n751), .ZN(new_n888));
  INV_X1    g0688(.A(new_n691), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n402), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(new_n658), .B2(new_n433), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT103), .B1(new_n428), .B2(new_n657), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT103), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n392), .A2(new_n397), .A3(new_n391), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n894), .A2(new_n398), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n383), .A2(KEYINPUT7), .A3(new_n286), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n298), .B1(new_n369), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n381), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n284), .B1(new_n898), .B2(KEYINPUT16), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n895), .B1(new_n899), .B2(new_n382), .ZN(new_n900));
  INV_X1    g0700(.A(new_n417), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n893), .B(new_n431), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n892), .A2(new_n890), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT37), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT37), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n434), .A2(new_n890), .A3(new_n905), .A4(new_n431), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n891), .B1(new_n907), .B2(KEYINPUT104), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n905), .B(new_n431), .C1(new_n900), .C2(new_n691), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n909), .A2(new_n421), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n903), .B2(KEYINPUT37), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT104), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT38), .B1(new_n908), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n361), .B1(new_n381), .B2(new_n897), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n915), .A2(new_n389), .A3(new_n285), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n401), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n889), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n436), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n917), .A2(new_n417), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n921), .A2(new_n918), .A3(new_n431), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT37), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n906), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n920), .A2(KEYINPUT38), .A3(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  OAI211_X1 g0726(.A(KEYINPUT40), .B(new_n888), .C1(new_n914), .C2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT38), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n430), .A2(new_n432), .B1(new_n434), .B2(KEYINPUT18), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n918), .B1(new_n929), .B2(new_n423), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n923), .A2(new_n906), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n925), .ZN(new_n933));
  INV_X1    g0733(.A(new_n887), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n879), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT40), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n927), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n731), .B1(new_n881), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n938), .B2(new_n881), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT106), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n867), .A2(new_n701), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n869), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n943), .A2(new_n933), .A3(new_n886), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n658), .B2(new_n889), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n882), .A2(new_n693), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n658), .A2(new_n433), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n900), .A2(new_n691), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n911), .B2(new_n912), .ZN(new_n950));
  AOI211_X1 g0750(.A(KEYINPUT104), .B(new_n910), .C1(KEYINPUT37), .C2(new_n903), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n928), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT39), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n952), .A2(new_n953), .A3(new_n925), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n933), .A2(KEYINPUT39), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n945), .B1(new_n946), .B2(new_n956), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n471), .B(new_n728), .C1(KEYINPUT29), .C2(new_n729), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n958), .A2(new_n662), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n957), .B(new_n959), .Z(new_n960));
  NOR2_X1   g0760(.A1(new_n941), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n941), .A2(new_n960), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n265), .B2(new_n687), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT107), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n964), .B2(new_n963), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n771), .B(G77), .C1(new_n298), .C2(new_n321), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n288), .A2(G68), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n265), .B(G13), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n215), .A2(new_n472), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n625), .B2(KEYINPUT35), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT102), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n971), .A2(new_n972), .B1(KEYINPUT35), .B2(new_n625), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n972), .B2(new_n971), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT36), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n969), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n966), .B(new_n976), .C1(new_n975), .C2(new_n974), .ZN(G367));
  NOR2_X1   g0777(.A1(new_n229), .A2(new_n770), .ZN(new_n978));
  INV_X1    g0778(.A(new_n445), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n766), .B1(new_n218), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n758), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n783), .A2(G68), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n849), .B2(new_n789), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n839), .A2(new_n319), .B1(new_n290), .B2(new_n786), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n983), .B(new_n984), .C1(new_n804), .C2(G143), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n252), .B1(new_n795), .B2(new_n321), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(G50), .B2(new_n847), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n985), .B(new_n987), .C1(new_n371), .C2(new_n798), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n815), .A2(KEYINPUT46), .A3(G116), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT46), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n795), .B2(new_n472), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n989), .B(new_n991), .C1(new_n812), .C2(new_n796), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n839), .A2(new_n492), .B1(new_n237), .B2(new_n786), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(G107), .B2(new_n783), .ZN(new_n994));
  INV_X1    g0794(.A(G317), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n383), .B1(new_n789), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(new_n799), .B2(G294), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n994), .B(new_n997), .C1(new_n813), .C2(new_n805), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n988), .B1(new_n992), .B2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT47), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n834), .B1(new_n999), .B2(new_n1000), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n981), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n671), .A2(new_n672), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n693), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1005), .A2(new_n603), .A3(new_n673), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n603), .B2(new_n1005), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1003), .B1(new_n763), .B2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT111), .Z(new_n1009));
  OAI21_X1  g0809(.A(new_n678), .B1(new_n630), .B2(new_n701), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n651), .A2(new_n642), .A3(new_n693), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n714), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT44), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n712), .A2(new_n713), .A3(new_n1012), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT45), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(KEYINPUT109), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n709), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n709), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1020), .A2(KEYINPUT109), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n708), .ZN(new_n1025));
  OR3_X1    g0825(.A1(new_n1025), .A2(KEYINPUT110), .A3(new_n710), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n698), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1025), .A2(new_n710), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1029), .A2(KEYINPUT110), .A3(new_n712), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n1028), .A2(new_n1030), .B1(new_n1023), .B2(KEYINPUT110), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n754), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1022), .A2(new_n1024), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n754), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n718), .B(KEYINPUT41), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n757), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OR3_X1    g0837(.A1(new_n712), .A2(KEYINPUT42), .A3(new_n1010), .ZN(new_n1038));
  OAI21_X1  g0838(.A(KEYINPUT42), .B1(new_n712), .B2(new_n1010), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n1012), .A2(new_n681), .B1(new_n664), .B2(new_n665), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1038), .B(new_n1039), .C1(new_n693), .C2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT108), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1007), .A2(KEYINPUT43), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1042), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n1045), .A2(new_n1046), .B1(KEYINPUT43), .B2(new_n1007), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1046), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1007), .A2(KEYINPUT43), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1048), .A2(new_n1049), .A3(new_n1044), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1047), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n709), .B2(new_n1013), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n709), .A2(new_n1013), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1047), .A2(new_n1050), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1009), .B1(new_n1037), .B2(new_n1055), .ZN(G387));
  NOR2_X1   g0856(.A1(new_n1033), .A2(new_n719), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n754), .B2(new_n1031), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1031), .A2(new_n757), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n770), .B1(new_n226), .B2(G45), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n720), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1060), .B1(new_n1061), .B2(new_n773), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  XOR2_X1   g0863(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n442), .B2(G50), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n443), .A2(new_n1064), .A3(new_n288), .ZN(new_n1067));
  AOI21_X1  g0867(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1066), .A2(new_n720), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1063), .A2(new_n1069), .B1(new_n235), .B2(new_n717), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n383), .B1(new_n837), .B2(G97), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n328), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1071), .B1(new_n796), .B2(new_n298), .C1(new_n1072), .C2(new_n798), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n979), .A2(new_n782), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(G150), .B2(new_n791), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n815), .A2(G77), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1075), .B(new_n1076), .C1(new_n288), .C2(new_n839), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1073), .B(new_n1077), .C1(G159), .C2(new_n804), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(KEYINPUT113), .B(G322), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n804), .A2(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n847), .A2(G303), .B1(new_n780), .B2(G317), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1080), .B(new_n1081), .C1(new_n813), .C2(new_n798), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT48), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n1083), .B1(new_n812), .B2(new_n782), .C1(new_n809), .C2(new_n795), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT49), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n383), .B1(new_n789), .B2(new_n821), .C1(new_n472), .C2(new_n786), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1078), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n758), .B1(new_n767), .B2(new_n1070), .C1(new_n1089), .C2(new_n834), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT114), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n708), .B2(new_n763), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1058), .B(new_n1059), .C1(new_n1092), .C2(new_n1094), .ZN(G393));
  OAI21_X1  g0895(.A(KEYINPUT115), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT115), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1016), .A2(new_n1019), .A3(new_n1098), .A4(new_n709), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n1096), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n718), .B(new_n1034), .C1(new_n1100), .C2(new_n1033), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1013), .A2(new_n762), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n805), .A2(new_n995), .B1(new_n813), .B2(new_n839), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT52), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n783), .A2(G116), .B1(new_n791), .B2(new_n1079), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n812), .B2(new_n795), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n252), .B1(new_n837), .B2(G107), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n1109), .B1(new_n798), .B2(new_n492), .C1(new_n809), .C2(new_n796), .ZN(new_n1110));
  NOR4_X1   g0910(.A1(new_n1105), .A2(new_n1106), .A3(new_n1108), .A4(new_n1110), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n804), .A2(G150), .B1(G159), .B2(new_n780), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT51), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n783), .A2(G77), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n791), .A2(G143), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1114), .B(new_n1115), .C1(new_n298), .C2(new_n795), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n383), .B1(new_n837), .B2(G87), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n1117), .B1(new_n798), .B2(new_n288), .C1(new_n442), .C2(new_n796), .ZN(new_n1118));
  NOR3_X1   g0918(.A1(new_n1113), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1111), .A2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1120), .A2(new_n834), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n241), .A2(new_n770), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n767), .B(new_n1122), .C1(G97), .C2(new_n717), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n1121), .A2(new_n759), .A3(new_n1123), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1100), .A2(new_n757), .B1(new_n1102), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1101), .A2(new_n1125), .ZN(G390));
  NAND2_X1  g0926(.A1(new_n952), .A2(new_n925), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n868), .B(new_n701), .C1(new_n725), .C2(new_n727), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n942), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT116), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n884), .A2(new_n1130), .A3(new_n885), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1130), .B1(new_n884), .B2(new_n885), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1129), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n946), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1127), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n946), .B1(new_n943), .B2(new_n886), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1136), .B1(new_n956), .B2(new_n1137), .ZN(new_n1138));
  AND4_X1   g0938(.A1(G330), .A2(new_n879), .A3(new_n865), .A4(new_n886), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n752), .A2(new_n865), .A3(new_n886), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1141), .B(new_n1136), .C1(new_n956), .C2(new_n1137), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n886), .B1(new_n752), .B2(new_n865), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n943), .B1(new_n1144), .B2(new_n1139), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1129), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n879), .A2(G330), .A3(new_n865), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1141), .B(new_n1146), .C1(new_n1147), .C2(new_n1133), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n471), .A2(G330), .A3(new_n879), .ZN(new_n1150));
  AND3_X1   g0950(.A1(new_n958), .A2(new_n662), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1143), .A2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1140), .A2(new_n1149), .A3(new_n1142), .A4(new_n1151), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1153), .A2(new_n718), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1140), .A2(new_n757), .A3(new_n1142), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n759), .B1(new_n1072), .B2(new_n832), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n780), .A2(G132), .B1(G50), .B2(new_n837), .ZN(new_n1158));
  INV_X1    g0958(.A(G125), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1158), .B1(new_n1159), .B2(new_n789), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n815), .A2(G150), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT53), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1160), .B(new_n1162), .C1(G128), .C2(new_n804), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n252), .B1(new_n371), .B2(new_n782), .C1(new_n798), .C2(new_n849), .ZN(new_n1164));
  XOR2_X1   g0964(.A(KEYINPUT54), .B(G143), .Z(new_n1165));
  AOI21_X1  g0965(.A(new_n1164), .B1(new_n847), .B2(new_n1165), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n780), .A2(G116), .B1(G294), .B2(new_n791), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1167), .B(new_n1114), .C1(new_n298), .C2(new_n786), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(G283), .B2(new_n804), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n383), .B1(new_n528), .B2(new_n795), .C1(new_n796), .C2(new_n237), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(G107), .B2(new_n799), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n1163), .A2(new_n1166), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1157), .B1(new_n834), .B2(new_n1172), .C1(new_n956), .C2(new_n761), .ZN(new_n1173));
  AND2_X1   g0973(.A1(new_n1156), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1155), .A2(new_n1174), .ZN(G378));
  NAND3_X1  g0975(.A1(new_n927), .A2(G330), .A3(new_n937), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(KEYINPUT119), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT119), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n927), .A2(new_n937), .A3(new_n1178), .A4(G330), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n360), .A2(new_n441), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n334), .A2(new_n691), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1180), .B(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1182), .B(new_n1183), .Z(new_n1184));
  NAND3_X1  g0984(.A1(new_n1177), .A2(new_n1179), .A3(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1182), .B(new_n1183), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n938), .A2(new_n1186), .A3(new_n1178), .A4(G330), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n957), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT120), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n957), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1185), .A2(new_n1191), .A3(new_n1187), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1189), .A2(new_n1190), .A3(new_n1192), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1185), .A2(new_n1191), .A3(KEYINPUT120), .A4(new_n1187), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1154), .A2(new_n1151), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT57), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1197), .B1(new_n1154), .B2(new_n1151), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1185), .A2(new_n1191), .A3(new_n1187), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1191), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1199), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n718), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1198), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1193), .A2(new_n757), .A3(new_n1194), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1186), .A2(new_n760), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n780), .A2(G107), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n791), .A2(G283), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n837), .A2(new_n379), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1208), .A2(new_n1076), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n252), .A2(G41), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n982), .A2(new_n1212), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(new_n237), .B2(new_n798), .C1(new_n979), .C2(new_n796), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1211), .B(new_n1214), .C1(G116), .C2(new_n804), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT117), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1216), .B(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(G33), .A2(G41), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(new_n1212), .A2(G50), .A3(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n815), .A2(new_n1165), .ZN(new_n1221));
  INV_X1    g1021(.A(G128), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1221), .B1(new_n839), .B2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(G150), .B2(new_n783), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G132), .A2(new_n799), .B1(new_n847), .B2(G137), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1224), .B(new_n1225), .C1(new_n1159), .C2(new_n805), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n1226), .A2(KEYINPUT59), .ZN(new_n1227));
  INV_X1    g1027(.A(G124), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1219), .B1(new_n789), .B2(new_n1228), .C1(new_n371), .C2(new_n786), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n1226), .B2(KEYINPUT59), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1220), .B1(new_n1227), .B2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n834), .B1(new_n1218), .B2(new_n1231), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n759), .B(new_n1232), .C1(new_n288), .C2(new_n832), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1207), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1206), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1205), .A2(new_n1236), .ZN(G375));
  INV_X1    g1037(.A(new_n1149), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1151), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1240), .A2(new_n1036), .A3(new_n1152), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n760), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1242), .A2(KEYINPUT121), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(KEYINPUT121), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n839), .A2(new_n812), .B1(new_n492), .B2(new_n789), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1074), .B(new_n1245), .C1(G97), .C2(new_n815), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n383), .B1(new_n290), .B2(new_n786), .C1(new_n798), .C2(new_n472), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G107), .B2(new_n847), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1246), .B(new_n1248), .C1(new_n809), .C2(new_n805), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(G150), .A2(new_n847), .B1(new_n799), .B2(new_n1165), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n780), .A2(G137), .B1(G50), .B2(new_n783), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1250), .A2(new_n252), .A3(new_n1210), .A4(new_n1251), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n795), .A2(new_n371), .B1(new_n1222), .B2(new_n789), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1253), .B(KEYINPUT122), .ZN(new_n1254));
  INV_X1    g1054(.A(G132), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1254), .B1(new_n805), .B2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1249), .B1(new_n1252), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n765), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n759), .B1(new_n298), .B2(new_n832), .ZN(new_n1259));
  AND4_X1   g1059(.A1(new_n1243), .A2(new_n1244), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n1149), .B2(new_n757), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1241), .A2(new_n1261), .ZN(G381));
  INV_X1    g1062(.A(G378), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1205), .A2(new_n1263), .A3(new_n1236), .ZN(new_n1264));
  OR4_X1    g1064(.A1(G396), .A2(G390), .A3(G393), .A4(G384), .ZN(new_n1265));
  OR4_X1    g1065(.A1(G387), .A2(new_n1264), .A3(new_n1265), .A4(G381), .ZN(G407));
  NAND2_X1  g1066(.A1(new_n692), .A2(G213), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(KEYINPUT123), .ZN(new_n1268));
  OAI211_X1 g1068(.A(G407), .B(G213), .C1(new_n1264), .C2(new_n1268), .ZN(G409));
  XNOR2_X1  g1069(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1268), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1205), .A2(G378), .A3(new_n1236), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n756), .B1(new_n1189), .B2(new_n1192), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(new_n1207), .B2(new_n1233), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1193), .A2(new_n1036), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1275));
  AOI21_X1  g1075(.A(G378), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1271), .B1(new_n1272), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT60), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1240), .A2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1238), .A2(new_n1239), .A3(KEYINPUT60), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1280), .A2(new_n718), .A3(new_n1152), .A4(new_n1281), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1282), .A2(G384), .A3(new_n1261), .ZN(new_n1283));
  AOI21_X1  g1083(.A(G384), .B1(new_n1282), .B2(new_n1261), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(G2897), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1285), .B1(new_n1286), .B2(new_n1267), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1271), .A2(G2897), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1287), .B1(new_n1285), .B2(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1270), .B1(new_n1278), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(KEYINPUT126), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT126), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1292), .B(new_n1270), .C1(new_n1278), .C2(new_n1289), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1203), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1294));
  NOR3_X1   g1094(.A1(new_n1294), .A2(new_n1263), .A3(new_n1235), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1267), .B(new_n1285), .C1(new_n1295), .C2(new_n1276), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT62), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1272), .A2(new_n1277), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1299), .A2(KEYINPUT62), .A3(new_n1268), .A4(new_n1285), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1291), .A2(new_n1293), .A3(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT124), .ZN(new_n1303));
  INV_X1    g1103(.A(G390), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1303), .B1(G387), .B2(new_n1304), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(G393), .B(new_n830), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1036), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1307), .B1(new_n1034), .B2(new_n754), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1054), .B(new_n1052), .C1(new_n1308), .C2(new_n757), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1309), .A2(G390), .A3(new_n1009), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(G390), .B1(new_n1309), .B2(new_n1009), .ZN(new_n1312));
  OAI22_X1  g1112(.A1(new_n1305), .A2(new_n1306), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1312), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(G393), .B(G396), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1314), .A2(new_n1303), .A3(new_n1310), .A4(new_n1315), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1313), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1302), .A2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1289), .B1(new_n1267), .B2(new_n1299), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT63), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1296), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1278), .A2(KEYINPUT63), .A3(new_n1285), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1317), .A2(KEYINPUT61), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1321), .A2(new_n1322), .A3(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1318), .A2(new_n1324), .ZN(G405));
  INV_X1    g1125(.A(KEYINPUT127), .ZN(new_n1326));
  OR2_X1    g1126(.A1(new_n1317), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1317), .A2(new_n1326), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(G375), .A2(new_n1263), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(new_n1272), .ZN(new_n1330));
  NOR3_X1   g1130(.A1(new_n1330), .A2(new_n1284), .A3(new_n1283), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1285), .B1(new_n1329), .B2(new_n1272), .ZN(new_n1332));
  OAI211_X1 g1132(.A(new_n1327), .B(new_n1328), .C1(new_n1331), .C2(new_n1332), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1334), .A2(new_n1326), .A3(new_n1317), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1333), .A2(new_n1335), .ZN(G402));
endmodule


