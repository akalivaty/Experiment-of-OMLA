//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 1 0 0 1 1 0 0 0 0 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n551, new_n552, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n565, new_n566, new_n567, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n608, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g025(.A1(G218), .A2(G221), .A3(G219), .A4(G220), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT67), .Z(new_n455));
  NAND2_X1  g030(.A1(new_n453), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  NAND2_X1  g032(.A1(new_n452), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n455), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(new_n462), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n462), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(G160));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  XOR2_X1   g052(.A(new_n477), .B(KEYINPUT69), .Z(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G112), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT70), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n475), .A2(new_n462), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(G124), .B2(new_n483), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n478), .A2(new_n484), .ZN(G162));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n487), .B(new_n488), .C1(new_n474), .C2(new_n473), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n488), .B1(new_n465), .B2(new_n487), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n465), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G126), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n462), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  OAI22_X1  g071(.A1(new_n493), .A2(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n492), .A2(new_n497), .ZN(G164));
  XNOR2_X1  g073(.A(KEYINPUT5), .B(G543), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n499), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  OR2_X1    g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  OAI211_X1 g080(.A(G50), .B(G543), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n507), .A2(new_n508), .B1(new_n504), .B2(new_n505), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT71), .B(G88), .ZN(new_n510));
  OAI211_X1 g085(.A(new_n503), .B(new_n506), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT71), .A2(G88), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT71), .A2(G88), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(new_n499), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n503), .B1(new_n517), .B2(new_n506), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n502), .B1(new_n512), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(G166));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  INV_X1    g097(.A(G89), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n522), .B1(new_n523), .B2(new_n509), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n525), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n516), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  AND2_X1   g104(.A1(G63), .A2(G651), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n529), .A2(G51), .B1(new_n499), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n526), .A2(new_n527), .A3(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT74), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n533), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(G168));
  AOI22_X1  g111(.A1(new_n499), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n501), .ZN(new_n538));
  INV_X1    g113(.A(G52), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n528), .A2(new_n539), .B1(new_n509), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  AOI22_X1  g117(.A1(new_n499), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n501), .ZN(new_n544));
  INV_X1    g119(.A(G43), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n528), .A2(new_n545), .B1(new_n509), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  NAND3_X1  g128(.A1(new_n516), .A2(G53), .A3(G543), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT9), .ZN(new_n555));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n508), .A2(new_n507), .ZN(new_n557));
  INV_X1    g132(.A(G65), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n509), .ZN(new_n560));
  AOI22_X1  g135(.A1(G651), .A2(new_n559), .B1(new_n560), .B2(G91), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n555), .A2(new_n561), .ZN(G299));
  INV_X1    g137(.A(G171), .ZN(G301));
  INV_X1    g138(.A(G168), .ZN(G286));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n519), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g141(.A(new_n502), .B(KEYINPUT75), .C1(new_n512), .C2(new_n518), .ZN(new_n567));
  AND2_X1   g142(.A1(new_n566), .A2(new_n567), .ZN(G303));
  NAND2_X1  g143(.A1(new_n560), .A2(G87), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n499), .B2(G74), .ZN(new_n571));
  INV_X1    g146(.A(G49), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n572), .B2(new_n528), .ZN(new_n573));
  OR3_X1    g148(.A1(new_n570), .A2(new_n573), .A3(KEYINPUT76), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT76), .B1(new_n570), .B2(new_n573), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G288));
  INV_X1    g152(.A(G48), .ZN(new_n578));
  INV_X1    g153(.A(G86), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n528), .A2(new_n578), .B1(new_n509), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n499), .A2(G61), .ZN(new_n581));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n501), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G305));
  AOI22_X1  g160(.A1(new_n499), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(new_n501), .ZN(new_n587));
  XOR2_X1   g162(.A(KEYINPUT77), .B(G47), .Z(new_n588));
  INV_X1    g163(.A(G85), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n528), .A2(new_n588), .B1(new_n509), .B2(new_n589), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n587), .A2(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n560), .A2(G92), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n593), .B(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n499), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n501), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(new_n597), .B2(new_n596), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n529), .A2(G54), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n595), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n592), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n592), .B1(new_n602), .B2(G868), .ZN(G321));
  NOR2_X1   g179(.A1(G299), .A2(G868), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g181(.A(new_n605), .B1(G168), .B2(G868), .ZN(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n602), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND2_X1  g184(.A1(new_n602), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n465), .A2(new_n463), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT12), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT13), .ZN(new_n616));
  INV_X1    g191(.A(G2100), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  AOI22_X1  g194(.A1(G123), .A2(new_n483), .B1(new_n476), .B2(G135), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  INV_X1    g196(.A(G111), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n621), .A2(KEYINPUT79), .B1(new_n622), .B2(G2105), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(KEYINPUT79), .B2(new_n621), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(G2096), .Z(new_n626));
  NAND3_X1  g201(.A1(new_n618), .A2(new_n619), .A3(new_n626), .ZN(G156));
  XNOR2_X1  g202(.A(KEYINPUT15), .B(G2435), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT81), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G2427), .B(G2430), .Z(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n632), .A2(KEYINPUT14), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G1341), .B(G1348), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n634), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G2451), .B(G2454), .Z(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(G14), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n638), .A2(new_n641), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(G401));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT82), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT17), .ZN(new_n649));
  XOR2_X1   g224(.A(G2067), .B(G2678), .Z(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2084), .B(G2090), .ZN(new_n652));
  NOR3_X1   g227(.A1(new_n649), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n652), .B1(new_n648), .B2(new_n651), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n654), .B1(new_n649), .B2(new_n651), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n650), .A2(new_n652), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n648), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT18), .ZN(new_n658));
  OR3_X1    g233(.A1(new_n653), .A2(new_n655), .A3(new_n658), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n659), .A2(KEYINPUT83), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(KEYINPUT83), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2096), .B(G2100), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n660), .A2(new_n661), .A3(new_n663), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1956), .B(G2474), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1961), .B(G1966), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n671), .B(new_n672), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n671), .A2(new_n672), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n670), .A2(new_n675), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n676), .A2(KEYINPUT20), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(KEYINPUT20), .ZN(new_n678));
  OAI221_X1 g253(.A(new_n673), .B1(new_n670), .B2(new_n674), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1991), .B(G1996), .Z(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1981), .B(G1986), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n681), .A2(new_n683), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n685), .B1(new_n684), .B2(new_n686), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(G229));
  XNOR2_X1  g265(.A(KEYINPUT87), .B(G16), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G20), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT23), .Z(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(G299), .B2(G16), .ZN(new_n694));
  INV_X1    g269(.A(G1956), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(G29), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G35), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G162), .B2(new_n697), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT29), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n696), .B1(new_n700), .B2(G2090), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT96), .Z(new_n702));
  NAND2_X1  g277(.A1(new_n602), .A2(G16), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G4), .B2(G16), .ZN(new_n704));
  INV_X1    g279(.A(G1348), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  INV_X1    g282(.A(G2084), .ZN(new_n708));
  INV_X1    g283(.A(G34), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n709), .A2(KEYINPUT24), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(KEYINPUT24), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n697), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G160), .B2(new_n697), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT94), .Z(new_n714));
  OAI211_X1 g289(.A(new_n706), .B(new_n707), .C1(new_n708), .C2(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT93), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT92), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT25), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n717), .A2(KEYINPUT92), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n717), .A2(KEYINPUT92), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n721), .A2(KEYINPUT25), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(G115), .A2(G2104), .ZN(new_n724));
  INV_X1    g299(.A(G127), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n475), .B2(new_n725), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n726), .A2(G2105), .B1(new_n476), .B2(G139), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n720), .A2(new_n723), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G29), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n697), .A2(G33), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI22_X1  g306(.A1(new_n700), .A2(G2090), .B1(G2072), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n714), .A2(new_n708), .ZN(new_n733));
  INV_X1    g308(.A(G16), .ZN(new_n734));
  NOR2_X1   g309(.A1(G171), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G5), .B2(new_n734), .ZN(new_n736));
  INV_X1    g311(.A(G1961), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n697), .A2(G32), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n476), .A2(G141), .B1(G105), .B2(new_n463), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n483), .A2(G129), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT26), .Z(new_n742));
  AND3_X1   g317(.A1(new_n739), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n738), .B1(new_n743), .B2(new_n697), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT27), .B(G1996), .Z(new_n745));
  AOI22_X1  g320(.A1(new_n736), .A2(new_n737), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n733), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT95), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n697), .A2(G27), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G164), .B2(new_n697), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n752), .A2(G2078), .ZN(new_n753));
  OAI221_X1 g328(.A(new_n753), .B1(new_n744), .B2(new_n745), .C1(new_n736), .C2(new_n737), .ZN(new_n754));
  INV_X1    g329(.A(new_n691), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n755), .A2(G19), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n548), .B2(new_n755), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G1341), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n752), .A2(G2078), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n620), .A2(G29), .A3(new_n624), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT30), .B(G28), .ZN(new_n761));
  OR2_X1    g336(.A1(KEYINPUT31), .A2(G11), .ZN(new_n762));
  NAND2_X1  g337(.A1(KEYINPUT31), .A2(G11), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n761), .A2(new_n697), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n759), .A2(new_n760), .A3(new_n764), .ZN(new_n765));
  NOR3_X1   g340(.A1(new_n754), .A2(new_n758), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n731), .A2(G2072), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR4_X1   g343(.A1(new_n715), .A2(new_n732), .A3(new_n750), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n476), .A2(G140), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n483), .A2(G128), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n462), .A2(G116), .ZN(new_n772));
  OAI21_X1  g347(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n770), .B(new_n771), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(G29), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT90), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n697), .A2(G26), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT28), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT91), .ZN(new_n780));
  INV_X1    g355(.A(G2067), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n734), .A2(G21), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G168), .B2(new_n734), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G1966), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n749), .B2(new_n748), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n702), .A2(new_n769), .A3(new_n782), .A4(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(G6), .A2(G16), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n584), .B2(G16), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT32), .ZN(new_n790));
  INV_X1    g365(.A(G1981), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n691), .A2(G22), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G166), .B2(new_n691), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n794), .A2(G1971), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(G1971), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n734), .A2(G23), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n570), .A2(new_n573), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(new_n734), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT33), .B(G1976), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n792), .A2(new_n795), .A3(new_n796), .A4(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT89), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT88), .B(KEYINPUT34), .Z(new_n804));
  OR2_X1    g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n697), .A2(G25), .ZN(new_n807));
  OR2_X1    g382(.A1(G95), .A2(G2105), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n808), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT85), .Z(new_n810));
  AOI22_X1  g385(.A1(G119), .A2(new_n483), .B1(new_n476), .B2(G131), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT86), .Z(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n807), .B1(new_n814), .B2(new_n697), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT35), .B(G1991), .Z(new_n816));
  XOR2_X1   g391(.A(new_n815), .B(new_n816), .Z(new_n817));
  MUX2_X1   g392(.A(G24), .B(G290), .S(new_n755), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(G1986), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n805), .A2(new_n806), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(KEYINPUT36), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n806), .A2(new_n820), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT36), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n823), .A2(new_n824), .A3(new_n805), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n787), .B1(new_n822), .B2(new_n825), .ZN(G311));
  INV_X1    g401(.A(new_n787), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n821), .A2(KEYINPUT36), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n824), .B1(new_n823), .B2(new_n805), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(G150));
  NAND2_X1  g405(.A1(new_n602), .A2(G559), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT38), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n499), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n833), .A2(new_n501), .ZN(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT97), .B(G55), .ZN(new_n835));
  INV_X1    g410(.A(G93), .ZN(new_n836));
  OAI22_X1  g411(.A1(new_n528), .A2(new_n835), .B1(new_n509), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n548), .B(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n832), .B(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n841), .A2(KEYINPUT39), .ZN(new_n842));
  INV_X1    g417(.A(G860), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(KEYINPUT39), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n838), .A2(new_n843), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT37), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(G145));
  INV_X1    g423(.A(KEYINPUT101), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n495), .A2(new_n496), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(new_n483), .B2(G126), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n487), .B1(new_n473), .B2(new_n474), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(KEYINPUT4), .ZN(new_n853));
  AND3_X1   g428(.A1(new_n853), .A2(KEYINPUT99), .A3(new_n489), .ZN(new_n854));
  AOI21_X1  g429(.A(KEYINPUT99), .B1(new_n853), .B2(new_n489), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n851), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n774), .ZN(new_n857));
  AOI22_X1  g432(.A1(G130), .A2(new_n483), .B1(new_n476), .B2(G142), .ZN(new_n858));
  OAI21_X1  g433(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n859));
  INV_X1    g434(.A(G118), .ZN(new_n860));
  AOI22_X1  g435(.A1(new_n859), .A2(KEYINPUT100), .B1(new_n860), .B2(G2105), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(KEYINPUT100), .B2(new_n859), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n857), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n728), .B(new_n743), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n812), .B(new_n615), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n866), .A2(new_n868), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n865), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(G162), .B(new_n625), .ZN(new_n873));
  XOR2_X1   g448(.A(G160), .B(KEYINPUT98), .Z(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n866), .A2(new_n868), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n876), .A2(new_n864), .A3(new_n869), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n872), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(G37), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n875), .B1(new_n872), .B2(new_n877), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n849), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n872), .A2(new_n877), .ZN(new_n883));
  INV_X1    g458(.A(new_n875), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n885), .A2(KEYINPUT101), .A3(new_n879), .A4(new_n878), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g463(.A(new_n519), .B(G290), .Z(new_n889));
  XNOR2_X1  g464(.A(G305), .B(new_n798), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n889), .B(new_n890), .Z(new_n891));
  XNOR2_X1  g466(.A(new_n610), .B(new_n839), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n601), .A2(G299), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n601), .A2(G299), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n894), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n601), .A2(G299), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT41), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n892), .B1(new_n897), .B2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n610), .B(new_n840), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n904), .A2(new_n895), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n891), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n902), .A2(new_n897), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n904), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n892), .A2(new_n900), .ZN(new_n909));
  INV_X1    g484(.A(new_n891), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  XOR2_X1   g486(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n912));
  AND3_X1   g487(.A1(new_n906), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n912), .B1(new_n906), .B2(new_n911), .ZN(new_n914));
  OAI21_X1  g489(.A(G868), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n838), .A2(G868), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(G295));
  INV_X1    g492(.A(KEYINPUT104), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n915), .A2(new_n918), .A3(new_n916), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n918), .B1(new_n915), .B2(new_n916), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(G331));
  NAND3_X1  g496(.A1(new_n534), .A2(new_n535), .A3(G301), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(G301), .B1(new_n534), .B2(new_n535), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n839), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(G168), .A2(G171), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(new_n840), .A3(new_n922), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n925), .A2(new_n927), .A3(new_n900), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n893), .A2(new_n894), .A3(new_n896), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(new_n900), .B2(KEYINPUT41), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n930), .B1(new_n927), .B2(new_n925), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n928), .B1(new_n931), .B2(KEYINPUT105), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n925), .A2(new_n927), .ZN(new_n933));
  INV_X1    g508(.A(new_n930), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n933), .A2(KEYINPUT105), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n891), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n925), .A2(new_n927), .A3(new_n900), .ZN(new_n937));
  AOI22_X1  g512(.A1(new_n925), .A2(new_n927), .B1(new_n902), .B2(new_n897), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(G37), .B1(new_n939), .B2(new_n910), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n936), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n933), .A2(new_n907), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n944), .A2(new_n910), .A3(new_n928), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n879), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n910), .B1(new_n944), .B2(new_n928), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT43), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n942), .A2(new_n943), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n891), .B1(new_n937), .B2(new_n938), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n940), .A2(KEYINPUT106), .A3(new_n941), .A4(new_n950), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n950), .A2(new_n945), .A3(new_n941), .A4(new_n879), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n933), .A2(new_n934), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT105), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n931), .A2(KEYINPUT105), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(new_n958), .A3(new_n928), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n946), .B1(new_n891), .B2(new_n959), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n951), .B(new_n954), .C1(new_n960), .C2(new_n941), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n949), .B1(KEYINPUT44), .B2(new_n961), .ZN(G397));
  INV_X1    g537(.A(G1966), .ZN(new_n963));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n964), .B1(new_n492), .B2(new_n497), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT117), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G40), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n468), .A2(new_n471), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n853), .A2(new_n489), .ZN(new_n970));
  AOI21_X1  g545(.A(G1384), .B1(new_n851), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT117), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(new_n972), .A3(KEYINPUT45), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n967), .A2(new_n969), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT45), .B1(new_n856), .B2(new_n964), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n963), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n856), .A2(new_n977), .A3(new_n964), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT109), .B1(new_n971), .B2(new_n977), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n856), .A2(KEYINPUT109), .A3(new_n977), .A4(new_n964), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n980), .A2(new_n708), .A3(new_n981), .A4(new_n969), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n976), .A2(new_n982), .A3(G168), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n983), .A2(new_n984), .A3(G8), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n976), .A2(new_n982), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(G286), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n987), .A2(G8), .A3(new_n983), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n985), .B1(new_n988), .B2(KEYINPUT51), .ZN(new_n989));
  XNOR2_X1  g564(.A(KEYINPUT112), .B(G1981), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT113), .B1(new_n584), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n993));
  NOR4_X1   g568(.A1(new_n580), .A2(new_n583), .A3(new_n993), .A4(new_n990), .ZN(new_n994));
  OAI22_X1  g569(.A1(new_n992), .A2(new_n994), .B1(new_n791), .B2(new_n584), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT49), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI221_X1 g572(.A(KEYINPUT49), .B1(new_n791), .B2(new_n584), .C1(new_n992), .C2(new_n994), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n856), .A2(new_n964), .A3(new_n969), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n999), .A2(G8), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n997), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n798), .A2(G1976), .ZN(new_n1003));
  INV_X1    g578(.A(G1976), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n574), .A2(new_n575), .A3(new_n1004), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1000), .A2(new_n1002), .A3(new_n1003), .A4(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n999), .A2(G8), .A3(new_n1003), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n1007), .A2(new_n1008), .A3(KEYINPUT52), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1008), .B1(new_n1007), .B2(KEYINPUT52), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1001), .B(new_n1006), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n566), .A2(G8), .A3(new_n567), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n566), .A2(KEYINPUT55), .A3(G8), .A4(new_n567), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n856), .A2(KEYINPUT45), .A3(new_n964), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n965), .A2(new_n966), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1017), .A2(new_n969), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1971), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n476), .A2(G137), .B1(G101), .B2(new_n463), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n469), .A2(new_n470), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1022), .B(G40), .C1(new_n462), .C2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1024), .B1(new_n977), .B2(new_n971), .ZN(new_n1025));
  INV_X1    g600(.A(G2090), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT99), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1027), .B1(new_n490), .B2(new_n491), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n853), .A2(KEYINPUT99), .A3(new_n489), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n497), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1030), .A2(G1384), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1025), .B(new_n1026), .C1(new_n977), .C2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1021), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1016), .B1(new_n1033), .B2(G8), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1011), .A2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n980), .A2(new_n1026), .A3(new_n981), .A4(new_n969), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT110), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1024), .B1(new_n978), .B2(new_n979), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT110), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1038), .A2(new_n1039), .A3(new_n1026), .A4(new_n981), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1037), .A2(new_n1040), .A3(new_n1021), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1041), .A2(G8), .A3(new_n1016), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1035), .A2(new_n1042), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1030), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT109), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1045), .B1(new_n965), .B2(KEYINPUT50), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n981), .B(new_n969), .C1(new_n1044), .C2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n737), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT123), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT123), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1047), .A2(new_n1050), .A3(new_n737), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n975), .A2(new_n1052), .A3(G2078), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1024), .B1(new_n1031), .B2(KEYINPUT45), .ZN(new_n1054));
  INV_X1    g629(.A(G2078), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1017), .A2(new_n1055), .A3(new_n969), .A4(new_n1018), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1053), .A2(new_n1054), .B1(new_n1056), .B2(new_n1052), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1049), .A2(G301), .A3(new_n1051), .A4(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1052), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n973), .A2(new_n969), .ZN(new_n1060));
  INV_X1    g635(.A(new_n975), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1052), .A2(G2078), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1060), .A2(new_n1061), .A3(new_n967), .A4(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1048), .A2(new_n1059), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(G171), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT54), .B1(new_n1058), .B2(new_n1065), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n989), .A2(new_n1043), .A3(new_n1066), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n1064), .A2(G171), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1049), .A2(new_n1051), .A3(new_n1057), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT124), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(G171), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1073));
  OAI211_X1 g648(.A(KEYINPUT54), .B(new_n1068), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1996), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1017), .A2(new_n1075), .A3(new_n969), .A4(new_n1018), .ZN(new_n1076));
  XOR2_X1   g651(.A(KEYINPUT58), .B(G1341), .Z(new_n1077));
  NAND2_X1  g652(.A1(new_n999), .A2(new_n1077), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT121), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT59), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n548), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  OAI22_X1  g657(.A1(new_n1079), .A2(new_n1082), .B1(KEYINPUT121), .B2(KEYINPUT59), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1084), .A2(new_n1080), .A3(new_n1081), .A4(new_n548), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT57), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1087), .A2(KEYINPUT57), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(G299), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n555), .A2(new_n561), .A3(KEYINPUT119), .A4(new_n1092), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n977), .B1(new_n856), .B2(new_n964), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n969), .B1(new_n965), .B2(KEYINPUT50), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n695), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT56), .B(G2072), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1017), .A2(new_n969), .A3(new_n1018), .A4(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1094), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1097), .A2(new_n1094), .A3(new_n1099), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1101), .A2(KEYINPUT61), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(KEYINPUT120), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1097), .A2(new_n1094), .A3(new_n1099), .A4(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1100), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1086), .B(new_n1103), .C1(new_n1107), .C2(KEYINPUT61), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n999), .A2(G2067), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1110), .B1(new_n1047), .B2(new_n705), .ZN(new_n1111));
  AOI211_X1 g686(.A(new_n1109), .B(new_n602), .C1(new_n1111), .C2(KEYINPUT60), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1047), .A2(new_n705), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1110), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(KEYINPUT60), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n601), .B1(new_n1115), .B2(KEYINPUT122), .ZN(new_n1116));
  OAI22_X1  g691(.A1(new_n1112), .A2(new_n1116), .B1(KEYINPUT122), .B2(new_n1115), .ZN(new_n1117));
  OR2_X1    g692(.A1(new_n1111), .A2(KEYINPUT60), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1108), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1111), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1100), .B1(new_n1120), .B2(new_n602), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1121), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1067), .B(new_n1074), .C1(new_n1119), .C2(new_n1122), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n986), .A2(G8), .A3(G168), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1035), .A2(new_n1042), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT63), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT118), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1125), .A2(new_n1129), .A3(new_n1126), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1011), .B(KEYINPUT114), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1041), .A2(G8), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1132), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1124), .A2(KEYINPUT63), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1131), .A2(new_n1042), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1128), .A2(new_n1130), .A3(new_n1135), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1064), .A2(G171), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1035), .A2(new_n1042), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT62), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1138), .B1(new_n1139), .B2(new_n989), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n983), .A2(G8), .ZN(new_n1141));
  AOI21_X1  g716(.A(G168), .B1(new_n976), .B2(new_n982), .ZN(new_n1142));
  OAI21_X1  g717(.A(KEYINPUT51), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n983), .A2(new_n984), .A3(G8), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT125), .B1(new_n1145), .B2(KEYINPUT62), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT125), .ZN(new_n1147));
  AOI211_X1 g722(.A(new_n1147), .B(new_n1139), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1140), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n576), .A2(new_n1004), .ZN(new_n1150));
  XOR2_X1   g725(.A(new_n1150), .B(KEYINPUT115), .Z(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n1001), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1152), .B1(new_n992), .B2(new_n994), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT116), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1000), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1156), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1042), .ZN(new_n1158));
  AOI22_X1  g733(.A1(new_n1155), .A2(new_n1157), .B1(new_n1131), .B2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1123), .A2(new_n1136), .A3(new_n1149), .A4(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n975), .A2(new_n969), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n774), .B(new_n781), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1163), .B1(new_n1075), .B2(new_n743), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1161), .A2(G1996), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1166), .A2(KEYINPUT107), .A3(new_n743), .ZN(new_n1167));
  AOI21_X1  g742(.A(KEYINPUT107), .B1(new_n1166), .B2(new_n743), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1165), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1169), .B(KEYINPUT108), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n812), .B(new_n816), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1170), .B1(new_n1161), .B2(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g747(.A(G290), .B(G1986), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1172), .B1(new_n1162), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1160), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1161), .B1(new_n743), .B2(new_n1163), .ZN(new_n1176));
  XOR2_X1   g751(.A(new_n1176), .B(KEYINPUT126), .Z(new_n1177));
  XOR2_X1   g752(.A(new_n1166), .B(KEYINPUT46), .Z(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1179), .B(KEYINPUT47), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n1161), .A2(G1986), .A3(G290), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(KEYINPUT48), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1180), .B1(new_n1172), .B2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1170), .A2(new_n814), .A3(new_n816), .ZN(new_n1184));
  OR2_X1    g759(.A1(new_n774), .A2(G2067), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1161), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1175), .A2(new_n1187), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g763(.A1(new_n665), .A2(G319), .A3(new_n645), .A4(new_n666), .ZN(new_n1190));
  INV_X1    g764(.A(new_n1190), .ZN(new_n1191));
  OAI211_X1 g765(.A(new_n1191), .B(KEYINPUT127), .C1(new_n688), .C2(new_n689), .ZN(new_n1192));
  INV_X1    g766(.A(KEYINPUT127), .ZN(new_n1193));
  OAI21_X1  g767(.A(new_n1193), .B1(G229), .B2(new_n1190), .ZN(new_n1194));
  NAND2_X1  g768(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g769(.A1(new_n942), .A2(new_n948), .ZN(new_n1196));
  NAND3_X1  g770(.A1(new_n1195), .A2(new_n887), .A3(new_n1196), .ZN(G225));
  INV_X1    g771(.A(G225), .ZN(G308));
endmodule


