//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 1 1 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G119), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G128), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT24), .B(G110), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT79), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n193), .B(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n187), .A2(KEYINPUT23), .A3(G119), .ZN(new_n196));
  INV_X1    g010(.A(new_n188), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n190), .B(new_n196), .C1(new_n197), .C2(KEYINPUT23), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT78), .ZN(new_n199));
  OR3_X1    g013(.A1(new_n198), .A2(new_n199), .A3(G110), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n199), .B1(new_n198), .B2(G110), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n195), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  OAI21_X1  g017(.A(G140), .B1(new_n203), .B2(KEYINPUT77), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT77), .ZN(new_n205));
  INV_X1    g019(.A(G140), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G125), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n207), .A3(KEYINPUT16), .ZN(new_n208));
  OR3_X1    g022(.A1(new_n203), .A2(KEYINPUT16), .A3(G140), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(G146), .A3(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(G125), .B(G140), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n202), .A2(new_n210), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n208), .A2(new_n209), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n215), .B(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n198), .A2(G110), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n217), .B1(new_n191), .B2(new_n192), .ZN(new_n218));
  OR2_X1    g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT80), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT80), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n214), .A2(new_n219), .A3(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT22), .B(G137), .ZN(new_n224));
  INV_X1    g038(.A(G953), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(G221), .A3(G234), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n224), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n227), .B(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n221), .A2(new_n223), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G902), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n214), .A2(new_n219), .A3(new_n229), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  OR2_X1    g048(.A1(new_n234), .A2(KEYINPUT25), .ZN(new_n235));
  INV_X1    g049(.A(G234), .ZN(new_n236));
  OAI21_X1  g050(.A(G217), .B1(new_n236), .B2(G902), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n237), .B1(new_n234), .B2(KEYINPUT25), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n231), .A2(new_n233), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT83), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n237), .A2(new_n232), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n239), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(G214), .B1(G237), .B2(G902), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(G116), .B(G119), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT5), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n189), .A2(G116), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n249), .B(G113), .C1(KEYINPUT5), .C2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT2), .ZN(new_n252));
  INV_X1    g066(.A(G113), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(KEYINPUT68), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n255), .B1(KEYINPUT2), .B2(G113), .ZN(new_n256));
  AOI22_X1  g070(.A1(new_n254), .A2(new_n256), .B1(KEYINPUT2), .B2(G113), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n248), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n251), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G107), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G104), .ZN(new_n261));
  INV_X1    g075(.A(G104), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G107), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G101), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT85), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT3), .B1(new_n262), .B2(G107), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT3), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(new_n260), .A3(G104), .ZN(new_n270));
  INV_X1    g084(.A(G101), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n268), .A2(new_n270), .A3(new_n271), .A4(new_n263), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n264), .A2(KEYINPUT85), .A3(G101), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n267), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  OR2_X1    g088(.A1(new_n259), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n272), .A2(KEYINPUT4), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n268), .A2(new_n270), .A3(new_n263), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G101), .ZN(new_n278));
  XOR2_X1   g092(.A(new_n276), .B(new_n278), .Z(new_n279));
  XOR2_X1   g093(.A(new_n257), .B(new_n248), .Z(new_n280));
  OAI21_X1  g094(.A(new_n275), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(G110), .B(G122), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n275), .B(new_n282), .C1(new_n279), .C2(new_n280), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(KEYINPUT6), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(G143), .B(G146), .ZN(new_n287));
  NAND2_X1  g101(.A1(KEYINPUT0), .A2(G128), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XOR2_X1   g103(.A(KEYINPUT0), .B(G128), .Z(new_n290));
  OAI211_X1 g104(.A(new_n289), .B(G125), .C1(new_n287), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n212), .A2(G143), .ZN(new_n292));
  INV_X1    g106(.A(G143), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G146), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n212), .A2(G143), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n295), .A2(new_n187), .B1(KEYINPUT1), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT1), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n287), .A2(new_n298), .A3(G128), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n291), .B1(new_n300), .B2(G125), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n225), .A2(G224), .ZN(new_n302));
  XOR2_X1   g116(.A(new_n302), .B(KEYINPUT88), .Z(new_n303));
  XNOR2_X1  g117(.A(new_n301), .B(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT6), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n281), .A2(new_n305), .A3(new_n283), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n286), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT90), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n291), .A2(new_n308), .B1(KEYINPUT7), .B2(new_n302), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n309), .B(new_n301), .ZN(new_n310));
  OR3_X1    g124(.A1(new_n259), .A2(new_n274), .A3(KEYINPUT89), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n259), .A2(new_n274), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT89), .B1(new_n259), .B2(new_n274), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n282), .B(KEYINPUT8), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n310), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(G902), .B1(new_n316), .B2(new_n285), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n307), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(G210), .B1(G237), .B2(G902), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n307), .A2(new_n317), .A3(new_n319), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n247), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G237), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(new_n225), .A3(G214), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n293), .ZN(new_n326));
  NOR2_X1   g140(.A1(G237), .A2(G953), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(G143), .A3(G214), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT66), .B(G131), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT17), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n329), .A2(new_n331), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n329), .A2(KEYINPUT17), .A3(new_n331), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n216), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(KEYINPUT91), .A2(KEYINPUT18), .A3(G131), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n204), .A2(new_n207), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G146), .ZN(new_n341));
  AOI22_X1  g155(.A1(new_n330), .A2(new_n339), .B1(new_n341), .B2(new_n213), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n342), .B1(new_n330), .B2(new_n339), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT95), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT95), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n338), .A2(new_n346), .A3(new_n343), .ZN(new_n347));
  XNOR2_X1  g161(.A(G113), .B(G122), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n348), .B(KEYINPUT92), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n349), .B(new_n262), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n345), .A2(KEYINPUT96), .A3(new_n347), .A4(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n338), .A2(new_n343), .A3(new_n350), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n350), .B1(new_n344), .B2(KEYINPUT95), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT96), .B1(new_n355), .B2(new_n347), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n232), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n333), .A2(new_n335), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n204), .A2(new_n207), .A3(KEYINPUT19), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n359), .B1(KEYINPUT19), .B2(new_n211), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n212), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n358), .A2(new_n361), .A3(new_n210), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n343), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n351), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n353), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT93), .ZN(new_n366));
  NOR2_X1   g180(.A1(G475), .A2(G902), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT93), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n364), .A2(new_n368), .A3(new_n353), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n366), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(KEYINPUT20), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT20), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n373), .B1(new_n364), .B2(new_n353), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT94), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n374), .B(new_n375), .ZN(new_n376));
  AOI22_X1  g190(.A1(new_n357), .A2(G475), .B1(new_n371), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G952), .ZN(new_n378));
  AOI211_X1 g192(.A(G953), .B(new_n378), .C1(G234), .C2(G237), .ZN(new_n379));
  XOR2_X1   g193(.A(KEYINPUT21), .B(G898), .Z(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(KEYINPUT100), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  AOI211_X1 g196(.A(new_n232), .B(new_n225), .C1(G234), .C2(G237), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n379), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n187), .A2(G143), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT97), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n386), .B(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G134), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n293), .A2(G128), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT98), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT98), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n388), .A2(new_n393), .A3(new_n389), .A4(new_n390), .ZN(new_n394));
  XNOR2_X1  g208(.A(G116), .B(G122), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(new_n260), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n386), .B(KEYINPUT97), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT13), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n390), .B(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(G134), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n392), .A2(new_n394), .A3(new_n396), .A4(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT14), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n395), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G122), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(G116), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n260), .B1(new_n405), .B2(KEYINPUT14), .ZN(new_n406));
  AOI22_X1  g220(.A1(new_n403), .A2(new_n406), .B1(new_n260), .B2(new_n395), .ZN(new_n407));
  INV_X1    g221(.A(new_n391), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n389), .B1(new_n388), .B2(new_n390), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(KEYINPUT9), .B(G234), .ZN(new_n411));
  INV_X1    g225(.A(G217), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n411), .A2(new_n412), .A3(G953), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n401), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n413), .B1(new_n401), .B2(new_n410), .ZN(new_n415));
  OR2_X1    g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n232), .ZN(new_n417));
  OR2_X1    g231(.A1(KEYINPUT99), .A2(KEYINPUT15), .ZN(new_n418));
  NAND2_X1  g232(.A1(KEYINPUT99), .A2(KEYINPUT15), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(G478), .A3(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n417), .B(new_n420), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n323), .A2(new_n377), .A3(new_n385), .A4(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G469), .ZN(new_n423));
  INV_X1    g237(.A(new_n300), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n424), .A2(new_n274), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n276), .B(new_n278), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n289), .B1(new_n287), .B2(new_n290), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT69), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT69), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n289), .B(new_n429), .C1(new_n287), .C2(new_n290), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  AOI22_X1  g245(.A1(KEYINPUT10), .A2(new_n425), .B1(new_n426), .B2(new_n431), .ZN(new_n432));
  AND2_X1   g246(.A1(KEYINPUT11), .A2(G134), .ZN(new_n433));
  OR2_X1    g247(.A1(KEYINPUT11), .A2(G134), .ZN(new_n434));
  INV_X1    g248(.A(G137), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  AND2_X1   g251(.A1(KEYINPUT64), .A2(G137), .ZN(new_n438));
  NOR2_X1   g252(.A1(KEYINPUT64), .A2(G137), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(KEYINPUT65), .B1(new_n440), .B2(new_n433), .ZN(new_n441));
  NAND2_X1  g255(.A1(KEYINPUT11), .A2(G134), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT65), .ZN(new_n443));
  NOR4_X1   g257(.A1(new_n438), .A2(new_n439), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n437), .B(new_n332), .C1(new_n441), .C2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G131), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT64), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n435), .ZN(new_n448));
  NAND2_X1  g262(.A1(KEYINPUT64), .A2(G137), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n449), .A3(new_n433), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n443), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n448), .A2(new_n433), .A3(KEYINPUT65), .A4(new_n449), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n436), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n445), .B1(new_n446), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n300), .A2(new_n272), .A3(new_n273), .A4(new_n267), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT86), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT10), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n457), .B1(new_n456), .B2(new_n458), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n432), .B(new_n455), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(G110), .B(G140), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(KEYINPUT84), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n225), .A2(G227), .ZN(new_n464));
  XOR2_X1   g278(.A(new_n463), .B(new_n464), .Z(new_n465));
  NAND2_X1  g279(.A1(new_n424), .A2(new_n274), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT87), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(new_n456), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT12), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n424), .A2(new_n274), .A3(KEYINPUT87), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n468), .A2(new_n469), .A3(new_n454), .A4(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n468), .A2(new_n454), .A3(new_n470), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT12), .ZN(new_n473));
  AND4_X1   g287(.A1(new_n461), .A2(new_n465), .A3(new_n471), .A4(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n459), .A2(new_n460), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n426), .A2(new_n431), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(new_n458), .B2(new_n456), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n454), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n465), .B1(new_n478), .B2(new_n461), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n423), .B(new_n232), .C1(new_n474), .C2(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n423), .A2(new_n232), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n461), .A2(new_n471), .A3(new_n473), .ZN(new_n483));
  INV_X1    g297(.A(new_n465), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n478), .A2(new_n461), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n485), .B1(new_n486), .B2(new_n484), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n480), .B(new_n482), .C1(new_n487), .C2(new_n423), .ZN(new_n488));
  OAI21_X1  g302(.A(G221), .B1(new_n411), .B2(G902), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n422), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT73), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT30), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n440), .A2(new_n389), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n446), .B1(G134), .B2(G137), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n297), .A2(new_n299), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n445), .ZN(new_n498));
  INV_X1    g312(.A(new_n427), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n437), .B1(new_n441), .B2(new_n444), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G131), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n499), .B1(new_n501), .B2(new_n445), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n498), .B1(new_n502), .B2(KEYINPUT67), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n454), .A2(KEYINPUT67), .A3(new_n427), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n494), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n280), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n497), .A2(new_n445), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n508), .B1(new_n454), .B2(new_n431), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT30), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n506), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n327), .A2(G210), .ZN(new_n512));
  XOR2_X1   g326(.A(new_n512), .B(KEYINPUT27), .Z(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(KEYINPUT26), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(new_n271), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n454), .A2(new_n431), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n516), .A2(new_n280), .A3(new_n498), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n511), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT31), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT31), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n511), .A2(new_n521), .A3(new_n515), .A4(new_n518), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n515), .B(KEYINPUT70), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n516), .A2(new_n498), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT72), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n507), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n509), .A2(KEYINPUT72), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT28), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n451), .A2(new_n452), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n446), .B1(new_n530), .B2(new_n437), .ZN(new_n531));
  AOI211_X1 g345(.A(new_n436), .B(new_n331), .C1(new_n451), .C2(new_n452), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n427), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT67), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n508), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n280), .B1(new_n535), .B2(new_n504), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT28), .B1(new_n536), .B2(new_n517), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT71), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n529), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI211_X1 g353(.A(KEYINPUT71), .B(KEYINPUT28), .C1(new_n536), .C2(new_n517), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n524), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n493), .B1(new_n523), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n533), .A2(new_n534), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(new_n504), .A3(new_n498), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n517), .B1(new_n544), .B2(new_n507), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT28), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n538), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n527), .A2(new_n528), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n546), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n547), .A2(new_n540), .A3(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n524), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n552), .A2(KEYINPUT73), .A3(new_n520), .A4(new_n522), .ZN(new_n553));
  NOR2_X1   g367(.A1(G472), .A2(G902), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n542), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT74), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT32), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n542), .A2(new_n553), .A3(KEYINPUT74), .A4(new_n554), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(G472), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n509), .A2(new_n280), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT28), .B1(new_n562), .B2(new_n517), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n549), .A2(KEYINPUT29), .A3(new_n515), .A4(new_n563), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n564), .A2(KEYINPUT76), .A3(new_n232), .ZN(new_n565));
  AOI21_X1  g379(.A(KEYINPUT76), .B1(new_n564), .B2(new_n232), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n547), .A2(new_n524), .A3(new_n540), .A4(new_n549), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT75), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n539), .A2(KEYINPUT75), .A3(new_n524), .A4(new_n540), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n511), .A2(new_n518), .ZN(new_n572));
  INV_X1    g386(.A(new_n515), .ZN(new_n573));
  AOI21_X1  g387(.A(KEYINPUT29), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n570), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n561), .B1(new_n567), .B2(new_n575), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n542), .A2(new_n553), .A3(new_n554), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n576), .B1(new_n577), .B2(KEYINPUT32), .ZN(new_n578));
  AOI211_X1 g392(.A(new_n245), .B(new_n492), .C1(new_n560), .C2(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(new_n271), .ZN(G3));
  NAND3_X1  g394(.A1(new_n542), .A2(new_n553), .A3(new_n232), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(G472), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n245), .A2(new_n490), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n557), .A2(new_n582), .A3(new_n559), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n323), .A2(new_n385), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT101), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n401), .A2(new_n410), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT33), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT33), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n416), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n587), .B1(new_n414), .B2(new_n415), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(new_n590), .A3(new_n589), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n232), .A2(G478), .ZN(new_n596));
  INV_X1    g410(.A(G478), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n595), .A2(new_n596), .B1(new_n597), .B2(new_n417), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n377), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n586), .A2(new_n599), .ZN(new_n600));
  OR2_X1    g414(.A1(new_n584), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT34), .B(G104), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G6));
  AND2_X1   g417(.A1(new_n366), .A2(new_n369), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n604), .A2(new_n372), .A3(new_n367), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n605), .A2(KEYINPUT102), .A3(new_n371), .ZN(new_n606));
  INV_X1    g420(.A(new_n421), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n357), .A2(G475), .ZN(new_n608));
  OR3_X1    g422(.A1(new_n370), .A2(KEYINPUT102), .A3(KEYINPUT20), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n606), .A2(new_n607), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n584), .A2(new_n585), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT35), .B(G107), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G9));
  NOR2_X1   g427(.A1(new_n230), .A2(KEYINPUT36), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT103), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n221), .A2(new_n223), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n244), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n618), .A2(new_n619), .B1(new_n235), .B2(new_n238), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n422), .A2(new_n490), .A3(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n621), .A2(new_n557), .A3(new_n582), .A4(new_n559), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT104), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT37), .B(G110), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G12));
  INV_X1    g439(.A(G900), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n383), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n379), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n610), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n323), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n620), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n490), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n631), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n560), .B2(new_n578), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(new_n187), .ZN(G30));
  XNOR2_X1  g451(.A(new_n629), .B(KEYINPUT39), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT40), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n321), .A2(new_n322), .ZN(new_n641));
  XOR2_X1   g455(.A(new_n641), .B(KEYINPUT38), .Z(new_n642));
  NAND2_X1  g456(.A1(new_n371), .A2(new_n376), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n608), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n607), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n620), .A2(new_n246), .ZN(new_n646));
  NOR4_X1   g460(.A1(new_n640), .A2(new_n642), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n562), .A2(new_n517), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n519), .B1(new_n524), .B2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n561), .B1(new_n649), .B2(new_n232), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n577), .B2(KEYINPUT32), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n560), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(new_n293), .ZN(G45));
  NAND2_X1  g468(.A1(new_n560), .A2(new_n578), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n377), .A2(new_n598), .A3(new_n630), .ZN(new_n656));
  AND3_X1   g470(.A1(new_n633), .A2(new_n634), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G146), .ZN(G48));
  INV_X1    g473(.A(new_n245), .ZN(new_n660));
  INV_X1    g474(.A(new_n489), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n232), .B1(new_n474), .B2(new_n479), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(G469), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n663), .A2(KEYINPUT105), .A3(new_n480), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n662), .A2(new_n665), .A3(G469), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n661), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n600), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n655), .A2(new_n660), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT41), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G113), .ZN(G15));
  NOR3_X1   g486(.A1(new_n668), .A2(new_n585), .A3(new_n610), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n655), .A2(new_n660), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G116), .ZN(G18));
  NAND2_X1  g489(.A1(new_n667), .A2(new_n323), .ZN(new_n676));
  INV_X1    g490(.A(new_n620), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n677), .A2(new_n421), .A3(new_n377), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n676), .A2(new_n678), .A3(new_n384), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n655), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G119), .ZN(G21));
  XNOR2_X1  g495(.A(KEYINPUT106), .B(G472), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n581), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n524), .B1(new_n549), .B2(new_n563), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n554), .B1(new_n523), .B2(new_n684), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n683), .A2(new_n660), .A3(new_n685), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n676), .A2(new_n384), .A3(new_n645), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT107), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G122), .ZN(G24));
  AND2_X1   g504(.A1(new_n683), .A2(new_n685), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n667), .A2(new_n323), .A3(new_n656), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n691), .A2(new_n677), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G125), .ZN(G27));
  NAND2_X1  g508(.A1(new_n487), .A2(KEYINPUT108), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n696), .B1(new_n486), .B2(new_n484), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n695), .A2(G469), .A3(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n480), .A3(new_n482), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n641), .A2(new_n661), .A3(new_n247), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n656), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n655), .A2(new_n660), .A3(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT42), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n555), .A2(new_n558), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n245), .B1(new_n578), .B2(new_n706), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n701), .A2(new_n702), .A3(new_n705), .ZN(new_n708));
  AOI22_X1  g522(.A1(new_n704), .A2(new_n705), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n446), .ZN(G33));
  NOR3_X1   g524(.A1(new_n701), .A2(new_n610), .A3(new_n630), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n655), .A2(new_n660), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G134), .ZN(G36));
  INV_X1    g527(.A(new_n480), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n695), .A2(KEYINPUT45), .A3(new_n697), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT45), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n423), .B1(new_n487), .B2(new_n716), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  OR2_X1    g532(.A1(new_n718), .A2(new_n481), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT46), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n714), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n721), .B1(new_n720), .B2(new_n719), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(new_n489), .A3(new_n638), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n557), .A2(new_n559), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n582), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n644), .A2(new_n598), .ZN(new_n726));
  XOR2_X1   g540(.A(new_n726), .B(KEYINPUT43), .Z(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n620), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n725), .A2(new_n728), .A3(KEYINPUT44), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT44), .B1(new_n725), .B2(new_n728), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n641), .A2(new_n247), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NOR4_X1   g547(.A1(new_n723), .A2(new_n730), .A3(new_n731), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n435), .ZN(G39));
  NAND2_X1  g549(.A1(new_n722), .A2(new_n489), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(KEYINPUT47), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n245), .A2(new_n656), .A3(new_n732), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n737), .A2(new_n655), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n206), .ZN(G42));
  NOR2_X1   g554(.A1(new_n727), .A2(new_n628), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n741), .A2(new_n686), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n742), .A2(new_n732), .ZN(new_n743));
  INV_X1    g557(.A(new_n737), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n744), .A2(KEYINPUT116), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n664), .A2(new_n666), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT117), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n661), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n748), .B1(new_n744), .B2(KEYINPUT116), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n743), .B1(new_n745), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(KEYINPUT118), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n742), .A2(new_n247), .A3(new_n642), .A4(new_n667), .ZN(new_n752));
  XOR2_X1   g566(.A(new_n752), .B(KEYINPUT50), .Z(new_n753));
  INV_X1    g567(.A(KEYINPUT118), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n754), .B(new_n743), .C1(new_n745), .C2(new_n749), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n667), .A2(new_n379), .A3(new_n732), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n727), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(KEYINPUT119), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n677), .A3(new_n691), .ZN(new_n759));
  OR3_X1    g573(.A1(new_n652), .A2(new_n245), .A3(new_n756), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n377), .A2(new_n598), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(KEYINPUT51), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n751), .A2(new_n753), .A3(new_n755), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n737), .A2(new_n748), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n743), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n766), .B(new_n753), .C1(KEYINPUT120), .C2(new_n762), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n762), .A2(KEYINPUT120), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT51), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n764), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT112), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n622), .B1(new_n584), .B2(new_n600), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n377), .A2(new_n607), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT110), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n586), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT110), .B1(new_n585), .B2(new_n774), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n584), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n773), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n579), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n772), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR4_X1   g597(.A1(new_n579), .A2(new_n773), .A3(new_n780), .A4(KEYINPUT111), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n655), .A2(new_n660), .A3(new_n711), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n606), .A2(new_n609), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n608), .A2(new_n421), .A3(new_n629), .ZN(new_n788));
  NOR4_X1   g602(.A1(new_n733), .A2(new_n490), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n655), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n691), .A2(new_n703), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n786), .B1(new_n792), .B2(new_n677), .ZN(new_n793));
  AOI22_X1  g607(.A1(new_n655), .A2(new_n679), .B1(new_n686), .B2(new_n687), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n794), .A2(new_n670), .A3(new_n674), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n704), .A2(new_n705), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n707), .A2(new_n708), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n793), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n771), .B1(new_n785), .B2(new_n799), .ZN(new_n800));
  AOI22_X1  g614(.A1(new_n655), .A2(new_n789), .B1(new_n691), .B2(new_n703), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n712), .B1(new_n801), .B2(new_n620), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n794), .A2(new_n670), .A3(new_n674), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n802), .A2(new_n709), .A3(new_n803), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n777), .A2(new_n778), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n724), .A2(new_n805), .A3(new_n582), .A4(new_n583), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n601), .A2(new_n806), .A3(new_n622), .ZN(new_n807));
  OAI21_X1  g621(.A(KEYINPUT111), .B1(new_n807), .B2(new_n579), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n781), .A2(new_n782), .A3(new_n772), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n804), .A2(new_n810), .A3(KEYINPUT112), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n645), .A2(new_n632), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n629), .B(KEYINPUT114), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n677), .A2(new_n661), .A3(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n652), .A2(new_n699), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n815), .A2(KEYINPUT52), .ZN(new_n816));
  AND4_X1   g630(.A1(new_n677), .A2(new_n692), .A3(new_n685), .A4(new_n683), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(new_n636), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n658), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(new_n658), .A3(new_n815), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n800), .A2(new_n811), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(KEYINPUT53), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n800), .A2(new_n811), .ZN(new_n826));
  INV_X1    g640(.A(new_n658), .ZN(new_n827));
  INV_X1    g641(.A(new_n635), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n655), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n693), .A3(KEYINPUT113), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT113), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n831), .B1(new_n817), .B2(new_n636), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n827), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n833), .A2(new_n816), .B1(new_n821), .B2(new_n820), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n834), .A2(KEYINPUT53), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n825), .B(KEYINPUT54), .C1(new_n826), .C2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n709), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n803), .A2(KEYINPUT115), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n794), .A2(new_n840), .A3(new_n670), .A4(new_n674), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n838), .A2(new_n839), .A3(new_n793), .A4(new_n841), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n842), .A2(new_n834), .A3(new_n785), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n843), .B1(new_n824), .B2(new_n837), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n758), .A2(new_n707), .ZN(new_n847));
  NOR2_X1   g661(.A1(KEYINPUT121), .A2(KEYINPUT48), .ZN(new_n848));
  AND2_X1   g662(.A1(KEYINPUT121), .A2(KEYINPUT48), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n676), .ZN(new_n851));
  AOI211_X1 g665(.A(new_n378), .B(G953), .C1(new_n742), .C2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n599), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n852), .B1(new_n853), .B2(new_n760), .ZN(new_n854));
  AOI211_X1 g668(.A(new_n850), .B(new_n854), .C1(new_n848), .C2(new_n847), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n770), .A2(new_n836), .A3(new_n846), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n378), .A2(new_n225), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n245), .A2(new_n661), .A3(new_n247), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT109), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n642), .A3(new_n726), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n859), .A2(new_n860), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n746), .B(KEYINPUT49), .Z(new_n864));
  OR4_X1    g678(.A1(new_n652), .A2(new_n862), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n858), .A2(new_n865), .ZN(G75));
  NOR2_X1   g680(.A1(new_n844), .A2(new_n232), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(G210), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT56), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n286), .A2(new_n306), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(new_n304), .Z(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT55), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n225), .A2(G952), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n870), .A2(new_n873), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n877), .A2(new_n878), .ZN(G51));
  XNOR2_X1  g693(.A(new_n481), .B(KEYINPUT57), .ZN(new_n880));
  AOI211_X1 g694(.A(KEYINPUT54), .B(new_n843), .C1(new_n837), .C2(new_n824), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n824), .A2(new_n837), .ZN(new_n882));
  INV_X1    g696(.A(new_n843), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n845), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n880), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n474), .A2(new_n479), .ZN(new_n888));
  OAI211_X1 g702(.A(KEYINPUT122), .B(new_n880), .C1(new_n881), .C2(new_n884), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n867), .A2(new_n718), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n875), .B1(new_n890), .B2(new_n891), .ZN(G54));
  AND2_X1   g706(.A1(KEYINPUT58), .A2(G475), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n867), .A2(new_n604), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n604), .B1(new_n867), .B2(new_n893), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n894), .A2(new_n895), .A3(new_n875), .ZN(G60));
  NAND2_X1  g710(.A1(G478), .A2(G902), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT59), .Z(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(new_n592), .B2(new_n594), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n899), .B1(new_n881), .B2(new_n884), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n900), .A2(KEYINPUT123), .A3(new_n876), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT123), .B1(new_n900), .B2(new_n876), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n898), .B1(new_n836), .B2(new_n846), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n903), .A2(new_n595), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(G63));
  NAND2_X1  g719(.A1(G217), .A2(G902), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT60), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n243), .B1(new_n844), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n876), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n844), .A2(new_n617), .A3(new_n907), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT61), .ZN(G66));
  INV_X1    g726(.A(G224), .ZN(new_n913));
  OAI21_X1  g727(.A(G953), .B1(new_n382), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n785), .A2(new_n803), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n914), .B1(new_n915), .B2(G953), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n871), .B1(G898), .B2(new_n225), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n916), .B(new_n917), .ZN(G69));
  NAND2_X1  g732(.A1(new_n506), .A2(new_n510), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n360), .B(KEYINPUT124), .Z(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n921), .B1(new_n626), .B2(new_n225), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n723), .A2(new_n632), .A3(new_n645), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n923), .A2(new_n707), .ZN(new_n924));
  OR4_X1    g738(.A1(new_n709), .A2(new_n739), .A3(new_n786), .A4(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n833), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n734), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT125), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n922), .B1(new_n929), .B2(new_n225), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n225), .B1(G227), .B2(G900), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n926), .A2(new_n653), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n932), .A2(KEYINPUT62), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n655), .A2(new_n660), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n732), .B1(new_n775), .B2(new_n599), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n934), .A2(new_n639), .A3(new_n935), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n739), .A2(new_n734), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n932), .A2(KEYINPUT62), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n933), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n921), .B1(new_n939), .B2(new_n225), .ZN(new_n940));
  OR3_X1    g754(.A1(new_n930), .A2(new_n931), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n931), .B1(new_n930), .B2(new_n940), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(G72));
  NAND2_X1  g757(.A1(G472), .A2(G902), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT63), .Z(new_n945));
  INV_X1    g759(.A(new_n915), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n945), .B1(new_n939), .B2(new_n946), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n572), .B(KEYINPUT126), .Z(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n949), .A2(new_n573), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n875), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n945), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(new_n929), .B2(new_n915), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n949), .A2(new_n573), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n825), .B1(new_n826), .B2(new_n835), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n572), .A2(new_n573), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n519), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n945), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n956), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  OR3_X1    g775(.A1(new_n957), .A2(new_n956), .A3(new_n960), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n955), .B1(new_n961), .B2(new_n962), .ZN(G57));
endmodule


