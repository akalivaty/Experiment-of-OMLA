//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 0 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 0 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n569, new_n570, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n604,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT66), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT67), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT68), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  AND2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n461), .A2(new_n463), .A3(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND4_X1  g041(.A1(new_n461), .A2(new_n463), .A3(G137), .A4(new_n459), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n459), .A2(G101), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n466), .A2(new_n469), .ZN(G160));
  NAND2_X1  g045(.A1(new_n461), .A2(new_n463), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(new_n459), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G124), .ZN(new_n473));
  XOR2_X1   g048(.A(new_n473), .B(KEYINPUT69), .Z(new_n474));
  OR2_X1    g049(.A1(G100), .A2(G2105), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n475), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n471), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  AND3_X1   g053(.A1(new_n474), .A2(new_n476), .A3(new_n478), .ZN(G162));
  OAI21_X1  g054(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(G114), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT70), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G114), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(KEYINPUT71), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT71), .ZN(new_n488));
  AOI211_X1 g063(.A(new_n488), .B(new_n459), .C1(new_n483), .C2(new_n485), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n481), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n461), .A2(new_n463), .A3(G138), .A4(new_n459), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT72), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g068(.A(KEYINPUT3), .B(G2104), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n494), .A2(KEYINPUT72), .A3(G138), .A4(new_n459), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n493), .A2(new_n495), .A3(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n491), .A2(new_n492), .A3(new_n497), .ZN(new_n498));
  AND3_X1   g073(.A1(new_n494), .A2(G126), .A3(G2105), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n490), .A2(new_n496), .A3(new_n498), .A4(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  OR2_X1    g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G50), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n504), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n508), .A2(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n506), .A2(new_n507), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT73), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI221_X1 g092(.A(KEYINPUT73), .B1(new_n513), .B2(new_n514), .C1(new_n506), .C2(new_n507), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(new_n508), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(new_n509), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G62), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n517), .A2(new_n518), .B1(G651), .B2(new_n524), .ZN(G166));
  NAND2_X1  g100(.A1(new_n505), .A2(G89), .ZN(new_n526));
  NAND2_X1  g101(.A1(G63), .A2(G651), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n522), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  INV_X1    g105(.A(G51), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n506), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n528), .A2(new_n532), .ZN(G168));
  AOI22_X1  g108(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G651), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(G52), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n506), .A2(new_n537), .B1(new_n513), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G171));
  AOI22_X1  g115(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n535), .ZN(new_n542));
  XNOR2_X1  g117(.A(KEYINPUT74), .B(G43), .ZN(new_n543));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n506), .A2(new_n543), .B1(new_n513), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(G188));
  NAND2_X1  g127(.A1(G78), .A2(G543), .ZN(new_n553));
  XNOR2_X1  g128(.A(KEYINPUT76), .B(G65), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n522), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n520), .A2(new_n509), .B1(new_n503), .B2(new_n504), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n555), .A2(G651), .B1(new_n556), .B2(G91), .ZN(new_n557));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  OAI21_X1  g133(.A(KEYINPUT9), .B1(new_n506), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(G543), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n560), .B1(new_n503), .B2(new_n504), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n561), .A2(new_n562), .A3(G53), .ZN(new_n563));
  AND3_X1   g138(.A1(new_n559), .A2(KEYINPUT75), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g139(.A(KEYINPUT75), .B1(new_n559), .B2(new_n563), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n557), .B1(new_n564), .B2(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  INV_X1    g142(.A(G168), .ZN(G286));
  NAND2_X1  g143(.A1(new_n517), .A2(new_n518), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n524), .A2(G651), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(G303));
  NAND2_X1  g146(.A1(new_n556), .A2(G87), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n561), .A2(G49), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  NAND3_X1  g150(.A1(new_n521), .A2(new_n505), .A3(G86), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n561), .A2(G48), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(new_n520), .B2(new_n509), .ZN(new_n580));
  AND2_X1   g155(.A1(G73), .A2(G543), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n578), .A2(new_n582), .ZN(G305));
  NAND2_X1  g158(.A1(new_n556), .A2(G85), .ZN(new_n584));
  XNOR2_X1  g159(.A(KEYINPUT77), .B(G47), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OAI221_X1 g161(.A(new_n584), .B1(new_n506), .B2(new_n585), .C1(new_n535), .C2(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n556), .A2(G92), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G66), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n522), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n594), .A2(G651), .B1(G54), .B2(new_n561), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n588), .B1(new_n597), .B2(G868), .ZN(G284));
  OAI21_X1  g173(.A(new_n588), .B1(new_n597), .B2(G868), .ZN(G321));
  NAND2_X1  g174(.A1(G286), .A2(G868), .ZN(new_n600));
  INV_X1    g175(.A(G299), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(G868), .ZN(G297));
  OAI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(G868), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n597), .B1(new_n604), .B2(G860), .ZN(G148));
  NAND2_X1  g180(.A1(new_n597), .A2(new_n604), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G868), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g184(.A(KEYINPUT12), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n477), .A2(new_n610), .A3(G2104), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n494), .A2(new_n459), .ZN(new_n612));
  OAI21_X1  g187(.A(KEYINPUT12), .B1(new_n612), .B2(new_n460), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  INV_X1    g190(.A(G2100), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n615), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n477), .A2(G135), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n472), .A2(G123), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n459), .A2(G111), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n619), .B(new_n620), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(G2096), .Z(new_n624));
  NAND3_X1  g199(.A1(new_n617), .A2(new_n618), .A3(new_n624), .ZN(G156));
  INV_X1    g200(.A(KEYINPUT14), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2427), .B(G2438), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2430), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT15), .B(G2435), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n626), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(new_n629), .B2(new_n628), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(G1341), .B(G1348), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n631), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  AND3_X1   g214(.A1(new_n638), .A2(G14), .A3(new_n639), .ZN(G401));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n643), .A2(KEYINPUT17), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n641), .A2(new_n642), .ZN(new_n645));
  AOI21_X1  g220(.A(KEYINPUT18), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  AOI21_X1  g222(.A(new_n647), .B1(new_n643), .B2(KEYINPUT18), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n646), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2096), .B(G2100), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(G227));
  XNOR2_X1  g226(.A(G1961), .B(G1966), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT78), .ZN(new_n653));
  XOR2_X1   g228(.A(G1956), .B(G2474), .Z(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1971), .B(G1976), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n653), .A2(new_n654), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n655), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(new_n657), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT20), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n658), .A2(KEYINPUT20), .A3(new_n657), .ZN(new_n663));
  OAI221_X1 g238(.A(new_n659), .B1(new_n657), .B2(new_n655), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G1991), .B(G1996), .Z(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1981), .B(G1986), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n666), .A2(new_n668), .ZN(new_n671));
  AND3_X1   g246(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n670), .B1(new_n669), .B2(new_n671), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(G229));
  NAND3_X1  g249(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT25), .Z(new_n676));
  INV_X1    g251(.A(G139), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n676), .B1(new_n677), .B2(new_n612), .ZN(new_n678));
  NAND2_X1  g253(.A1(G115), .A2(G2104), .ZN(new_n679));
  INV_X1    g254(.A(G127), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n679), .B1(new_n471), .B2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT88), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n459), .B1(new_n681), .B2(new_n682), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n678), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(G29), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(new_n686), .B2(G33), .ZN(new_n688));
  INV_X1    g263(.A(G2072), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT89), .Z(new_n691));
  XOR2_X1   g266(.A(KEYINPUT82), .B(G16), .Z(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G20), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT96), .B(KEYINPUT23), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n601), .B2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G1956), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(G171), .A2(new_n696), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G5), .B2(new_n696), .ZN(new_n701));
  INV_X1    g276(.A(G1961), .ZN(new_n702));
  INV_X1    g277(.A(G2084), .ZN(new_n703));
  NAND2_X1  g278(.A1(G160), .A2(G29), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT90), .B(KEYINPUT24), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(G34), .Z(new_n706));
  OAI21_X1  g281(.A(new_n704), .B1(G29), .B2(new_n706), .ZN(new_n707));
  AOI22_X1  g282(.A1(new_n701), .A2(new_n702), .B1(new_n703), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(new_n702), .B2(new_n701), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n686), .A2(G26), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT28), .Z(new_n711));
  NAND2_X1  g286(.A1(new_n477), .A2(G140), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT87), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n459), .A2(G116), .ZN(new_n715));
  OAI21_X1  g290(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  AOI22_X1  g292(.A1(new_n472), .A2(G128), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n711), .B1(new_n719), .B2(G29), .ZN(new_n720));
  INV_X1    g295(.A(G2067), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n688), .A2(new_n689), .ZN(new_n723));
  NOR3_X1   g298(.A1(new_n709), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n686), .A2(G27), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT93), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n501), .B2(G29), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT94), .B(G2078), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n691), .A2(new_n699), .A3(new_n724), .A4(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n686), .A2(G35), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT95), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G162), .B2(new_n686), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT29), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G2090), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n472), .A2(G129), .ZN(new_n736));
  NAND3_X1  g311(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT91), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT26), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n477), .A2(G141), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n459), .A2(G105), .A3(G2104), .ZN(new_n741));
  AND4_X1   g316(.A1(new_n736), .A2(new_n739), .A3(new_n740), .A4(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n742), .A2(new_n686), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n686), .B2(G32), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT27), .B(G1996), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT92), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n692), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(G19), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n546), .B2(new_n748), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT86), .B(G1341), .Z(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT30), .B(G28), .ZN(new_n753));
  OR2_X1    g328(.A1(KEYINPUT31), .A2(G11), .ZN(new_n754));
  NAND2_X1  g329(.A1(KEYINPUT31), .A2(G11), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n753), .A2(new_n686), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI221_X1 g331(.A(new_n756), .B1(new_n686), .B2(new_n623), .C1(new_n707), .C2(new_n703), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n752), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n696), .A2(G21), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G168), .B2(new_n696), .ZN(new_n760));
  INV_X1    g335(.A(G1966), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n747), .A2(new_n758), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G4), .A2(G16), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n597), .B2(G16), .ZN(new_n765));
  INV_X1    g340(.A(G1348), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n744), .B2(new_n746), .ZN(new_n768));
  NOR4_X1   g343(.A1(new_n730), .A2(new_n735), .A3(new_n763), .A4(new_n768), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT97), .Z(new_n770));
  NAND2_X1  g345(.A1(G166), .A2(new_n748), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G22), .B2(new_n748), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT84), .B(G1971), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  MUX2_X1   g350(.A(G6), .B(G305), .S(G16), .Z(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT32), .B(G1981), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT83), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n776), .B(new_n778), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n774), .A2(new_n775), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n696), .A2(G23), .ZN(new_n781));
  INV_X1    g356(.A(G288), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(new_n696), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT33), .ZN(new_n784));
  INV_X1    g359(.A(G1976), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n780), .A2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT34), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT85), .ZN(new_n790));
  MUX2_X1   g365(.A(G24), .B(G290), .S(new_n748), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1986), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n477), .A2(G131), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n472), .A2(G119), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n459), .A2(G107), .ZN(new_n795));
  OAI21_X1  g370(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n793), .B(new_n794), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT79), .ZN(new_n798));
  MUX2_X1   g373(.A(G25), .B(new_n798), .S(G29), .Z(new_n799));
  XOR2_X1   g374(.A(KEYINPUT35), .B(G1991), .Z(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT80), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT81), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n799), .B(new_n802), .ZN(new_n803));
  AOI211_X1 g378(.A(new_n792), .B(new_n803), .C1(new_n787), .C2(new_n788), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n790), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT36), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n770), .A2(new_n806), .ZN(G150));
  INV_X1    g382(.A(G150), .ZN(G311));
  NAND2_X1  g383(.A1(new_n597), .A2(G559), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT38), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(new_n535), .ZN(new_n812));
  INV_X1    g387(.A(G55), .ZN(new_n813));
  INV_X1    g388(.A(G93), .ZN(new_n814));
  OAI22_X1  g389(.A1(new_n506), .A2(new_n813), .B1(new_n513), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n546), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n546), .A2(new_n816), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n810), .B(new_n820), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n821), .A2(KEYINPUT39), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n821), .A2(KEYINPUT39), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n822), .A2(new_n823), .A3(G860), .ZN(new_n824));
  OAI21_X1  g399(.A(G860), .B1(new_n812), .B2(new_n815), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT98), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT37), .Z(new_n827));
  OR2_X1    g402(.A1(new_n824), .A2(new_n827), .ZN(G145));
  NAND2_X1  g403(.A1(new_n477), .A2(G142), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n472), .A2(G130), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n459), .A2(G118), .ZN(new_n831));
  OAI21_X1  g406(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n829), .B(new_n830), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(new_n614), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n797), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT101), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n719), .B(new_n501), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(new_n742), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n837), .A2(new_n742), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT100), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n685), .A2(new_n841), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n839), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n685), .B(new_n841), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n837), .A2(new_n742), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n844), .B1(new_n845), .B2(new_n838), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n836), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n845), .A2(new_n841), .A3(new_n685), .A4(new_n838), .ZN(new_n848));
  INV_X1    g423(.A(new_n835), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n839), .A2(new_n840), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n848), .B(new_n849), .C1(new_n850), .C2(new_n844), .ZN(new_n851));
  XOR2_X1   g426(.A(G160), .B(KEYINPUT99), .Z(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n623), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(G162), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n847), .A2(new_n851), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(KEYINPUT102), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT102), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n847), .A2(new_n851), .A3(new_n857), .A4(new_n854), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT101), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n835), .B(new_n860), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n861), .B(new_n848), .C1(new_n850), .C2(new_n844), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n854), .B1(new_n862), .B2(new_n847), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n863), .A2(G37), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g441(.A(G303), .B(G290), .ZN(new_n867));
  XNOR2_X1  g442(.A(G305), .B(G288), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n867), .B(new_n868), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT42), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n601), .A2(new_n596), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n597), .A2(G299), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n872), .A3(KEYINPUT103), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT41), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n874), .B(new_n875), .C1(KEYINPUT103), .C2(new_n871), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n871), .A2(new_n872), .A3(KEYINPUT41), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n606), .B(new_n819), .Z(new_n879));
  MUX2_X1   g454(.A(new_n873), .B(new_n878), .S(new_n879), .Z(new_n880));
  AND2_X1   g455(.A1(new_n870), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n870), .A2(new_n880), .ZN(new_n882));
  OAI21_X1  g457(.A(G868), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(G868), .B2(new_n816), .ZN(G295));
  OAI21_X1  g459(.A(new_n883), .B1(G868), .B2(new_n816), .ZN(G331));
  NAND2_X1  g460(.A1(G301), .A2(KEYINPUT105), .ZN(new_n886));
  OR3_X1    g461(.A1(new_n536), .A2(new_n539), .A3(KEYINPUT105), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n886), .A2(G168), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(G168), .B1(new_n886), .B2(new_n887), .ZN(new_n889));
  OR3_X1    g464(.A1(new_n888), .A2(new_n889), .A3(new_n819), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n819), .B1(new_n888), .B2(new_n889), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n878), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n869), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  OAI211_X1 g471(.A(KEYINPUT106), .B(new_n819), .C1(new_n888), .C2(new_n889), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n896), .A2(new_n890), .A3(new_n873), .A4(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n893), .A2(new_n894), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT107), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n893), .A2(new_n898), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n869), .ZN(new_n902));
  INV_X1    g477(.A(G37), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n893), .A2(new_n894), .A3(new_n904), .A4(new_n898), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n900), .A2(new_n902), .A3(new_n903), .A4(new_n905), .ZN(new_n906));
  XOR2_X1   g481(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n896), .A2(new_n890), .A3(new_n897), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n874), .B(KEYINPUT41), .C1(KEYINPUT103), .C2(new_n871), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n910), .B(new_n911), .C1(KEYINPUT41), .C2(new_n873), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n890), .A2(new_n873), .A3(new_n891), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n869), .ZN(new_n915));
  AOI21_X1  g490(.A(G37), .B1(new_n899), .B2(KEYINPUT107), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n915), .A2(new_n916), .A3(new_n905), .A4(new_n907), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n909), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n918), .A2(KEYINPUT44), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n915), .A2(new_n916), .A3(new_n905), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT43), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n921), .B1(new_n906), .B2(new_n908), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n919), .B1(KEYINPUT44), .B2(new_n922), .ZN(G397));
  INV_X1    g498(.A(KEYINPUT126), .ZN(new_n924));
  INV_X1    g499(.A(G1384), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n501), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT45), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n464), .A2(new_n465), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(G2105), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n467), .A2(new_n468), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n931), .A3(G40), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(G160), .A2(KEYINPUT108), .A3(G40), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n928), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n719), .A2(G2067), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n714), .A2(new_n721), .A3(new_n718), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n941), .A2(KEYINPUT109), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(KEYINPUT109), .ZN(new_n943));
  INV_X1    g518(.A(G1996), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n742), .B(new_n944), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n942), .A2(new_n943), .B1(new_n937), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n797), .B(new_n801), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n937), .A2(new_n947), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(G290), .A2(G1986), .ZN(new_n950));
  AND2_X1   g525(.A1(G290), .A2(G1986), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n937), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT110), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n949), .A2(KEYINPUT110), .A3(new_n952), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT112), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT55), .ZN(new_n959));
  NAND4_X1  g534(.A1(G303), .A2(new_n958), .A3(new_n959), .A4(G8), .ZN(new_n960));
  NAND2_X1  g535(.A1(KEYINPUT112), .A2(KEYINPUT55), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n958), .A2(new_n959), .ZN(new_n962));
  INV_X1    g537(.A(G8), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n961), .B(new_n962), .C1(G166), .C2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n960), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G2090), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n926), .A2(KEYINPUT50), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT108), .B1(G160), .B2(G40), .ZN(new_n969));
  INV_X1    g544(.A(G40), .ZN(new_n970));
  NOR4_X1   g545(.A1(new_n466), .A2(new_n469), .A3(new_n933), .A4(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g547(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n973));
  NAND3_X1  g548(.A1(new_n501), .A2(new_n925), .A3(new_n973), .ZN(new_n974));
  AND4_X1   g549(.A1(new_n967), .A2(new_n968), .A3(new_n972), .A4(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n936), .B1(new_n926), .B2(new_n927), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n925), .ZN(new_n977));
  AOI21_X1  g552(.A(G1971), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n966), .B(G8), .C1(new_n975), .C2(new_n978), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n501), .A2(new_n934), .A3(new_n925), .A4(new_n935), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n782), .A2(G1976), .ZN(new_n981));
  XNOR2_X1  g556(.A(KEYINPUT113), .B(G1976), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT52), .B1(G288), .B2(new_n982), .ZN(new_n983));
  AND4_X1   g558(.A1(G8), .A2(new_n980), .A3(new_n981), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT114), .ZN(new_n985));
  INV_X1    g560(.A(G1981), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n582), .A2(new_n576), .A3(new_n986), .A4(new_n577), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT115), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT115), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n578), .A2(new_n989), .A3(new_n986), .A4(new_n582), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(G305), .A2(G1981), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT49), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(KEYINPUT70), .B(G114), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n488), .B1(new_n995), .B2(new_n459), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n486), .A2(KEYINPUT71), .A3(G2105), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n480), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n498), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n998), .A2(new_n999), .A3(new_n499), .ZN(new_n1000));
  AOI21_X1  g575(.A(G1384), .B1(new_n1000), .B2(new_n496), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n963), .B1(new_n1001), .B2(new_n972), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n991), .A2(KEYINPUT49), .A3(new_n992), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n994), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n985), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n980), .A2(G8), .A3(new_n981), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT52), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n984), .B1(new_n1007), .B2(KEYINPUT114), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n979), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1002), .B(KEYINPUT116), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1004), .A2(new_n785), .A3(new_n782), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1010), .B1(new_n1011), .B2(new_n991), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n984), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1006), .A2(KEYINPUT52), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n991), .A2(KEYINPUT49), .A3(new_n992), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1018), .A2(new_n993), .ZN(new_n1019));
  AOI22_X1  g594(.A1(new_n1019), .A2(new_n1002), .B1(new_n984), .B2(KEYINPUT114), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n979), .A2(new_n1017), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n501), .A2(new_n1022), .A3(new_n925), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT117), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT117), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n501), .A2(new_n1025), .A3(new_n1022), .A4(new_n925), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n973), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n936), .B1(new_n926), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n967), .A3(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n928), .A2(new_n972), .A3(new_n977), .ZN(new_n1031));
  INV_X1    g606(.A(G1971), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n966), .B1(new_n1034), .B2(G8), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1021), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1031), .A2(new_n761), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n968), .A2(new_n703), .A3(new_n972), .A4(new_n974), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(G168), .A2(G8), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT63), .B1(new_n1036), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n936), .B1(new_n926), .B2(KEYINPUT50), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1043), .A2(new_n967), .A3(new_n974), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n963), .B1(new_n1033), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n965), .B1(new_n1045), .B2(KEYINPUT118), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n1047));
  AOI211_X1 g622(.A(new_n1047), .B(new_n963), .C1(new_n1033), .C2(new_n1044), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT63), .ZN(new_n1051));
  AOI211_X1 g626(.A(new_n1051), .B(new_n1040), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1050), .A2(new_n979), .A3(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1013), .B1(new_n1042), .B2(new_n1054), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n925), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT45), .B1(new_n501), .B2(new_n925), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1056), .A2(new_n1057), .A3(new_n936), .ZN(new_n1058));
  OAI211_X1 g633(.A(G168), .B(new_n1038), .C1(new_n1058), .C2(G1966), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(G8), .ZN(new_n1060));
  AOI21_X1  g635(.A(G168), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT51), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT62), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT51), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1059), .A2(new_n1064), .A3(G8), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1062), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1063), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1035), .ZN(new_n1069));
  INV_X1    g644(.A(G2078), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n928), .A2(new_n1070), .A3(new_n972), .A4(new_n977), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n968), .A2(new_n972), .A3(new_n974), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n702), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n976), .A2(KEYINPUT53), .A3(new_n1070), .A4(new_n977), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1073), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(G171), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1069), .A2(new_n1079), .A3(new_n979), .A4(new_n1050), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n1067), .A2(new_n1068), .A3(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1055), .A2(new_n1081), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n932), .A2(new_n1072), .A3(G2078), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n928), .A2(new_n977), .A3(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1073), .A2(new_n1075), .A3(G301), .A4(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT123), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1072), .A2(new_n1071), .B1(new_n1074), .B2(new_n702), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1088), .A2(KEYINPUT123), .A3(G301), .A4(new_n1084), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1087), .A2(new_n1089), .A3(new_n1078), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1088), .A2(new_n1084), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(G171), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1094), .B(KEYINPUT54), .C1(G171), .C2(new_n1077), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1096));
  AND4_X1   g671(.A1(new_n1092), .A2(new_n1095), .A3(new_n1096), .A4(new_n1036), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n698), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n1100));
  XNOR2_X1  g675(.A(KEYINPUT56), .B(G2072), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n976), .A2(new_n1100), .A3(new_n977), .A4(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n928), .A2(new_n972), .A3(new_n977), .A4(new_n1101), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT119), .ZN(new_n1104));
  NAND2_X1  g679(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT57), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n559), .A2(new_n563), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n557), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1099), .A2(new_n1102), .A3(new_n1104), .A4(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(KEYINPUT61), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1109), .A2(KEYINPUT121), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT121), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1114), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1104), .A2(new_n1102), .ZN(new_n1117));
  AOI21_X1  g692(.A(G1956), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1116), .B(KEYINPUT122), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1112), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1001), .A2(KEYINPUT120), .A3(new_n972), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n980), .A2(new_n1125), .ZN(new_n1126));
  XOR2_X1   g701(.A(KEYINPUT58), .B(G1341), .Z(new_n1127));
  NAND3_X1  g702(.A1(new_n1124), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n928), .A2(new_n944), .A3(new_n972), .A4(new_n977), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n546), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(KEYINPUT59), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1130), .A2(new_n1133), .A3(new_n546), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(G2067), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1136));
  AOI21_X1  g711(.A(G1348), .B1(new_n1043), .B2(new_n974), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1136), .A2(new_n1137), .A3(new_n597), .ZN(new_n1138));
  AOI21_X1  g713(.A(KEYINPUT120), .B1(new_n1001), .B2(new_n972), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n980), .A2(new_n1125), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n721), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1074), .A2(new_n766), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n596), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(KEYINPUT60), .B1(new_n1138), .B2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n596), .A2(KEYINPUT60), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1141), .A2(new_n1142), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1135), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1109), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT61), .B1(new_n1148), .B2(new_n1111), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n1123), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1111), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1143), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1097), .B1(new_n1150), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n957), .B1(new_n1082), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n937), .A2(new_n950), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT125), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1158), .B(KEYINPUT48), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(new_n949), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT46), .ZN(new_n1161));
  INV_X1    g736(.A(new_n937), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1161), .B1(new_n1162), .B2(G1996), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n937), .A2(KEYINPUT46), .A3(new_n944), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n938), .A2(new_n742), .A3(new_n939), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1163), .B(new_n1164), .C1(new_n1162), .C2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1166), .B(KEYINPUT47), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1160), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n798), .A2(new_n801), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n946), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n939), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1162), .B1(new_n1172), .B2(KEYINPUT124), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT124), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1168), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n924), .B1(new_n1156), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(new_n957), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1092), .A2(new_n1095), .A3(new_n1096), .A4(new_n1036), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1123), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1154), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1180), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NOR4_X1   g760(.A1(new_n1021), .A2(new_n1035), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1186));
  OAI22_X1  g761(.A1(new_n1186), .A2(KEYINPUT63), .B1(new_n1049), .B2(new_n1053), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1096), .A2(KEYINPUT62), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1188), .A2(new_n1079), .A3(new_n1036), .A4(new_n1066), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1187), .A2(new_n1189), .A3(new_n1013), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1179), .B1(new_n1185), .B2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1191), .A2(KEYINPUT126), .A3(new_n1176), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1178), .A2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g768(.A(G319), .ZN(new_n1195));
  NOR3_X1   g769(.A1(G401), .A2(new_n1195), .A3(G227), .ZN(new_n1196));
  OAI21_X1  g770(.A(new_n1196), .B1(new_n672), .B2(new_n673), .ZN(new_n1197));
  AOI21_X1  g771(.A(new_n1197), .B1(new_n859), .B2(new_n864), .ZN(new_n1198));
  AND3_X1   g772(.A1(new_n1198), .A2(new_n918), .A3(KEYINPUT127), .ZN(new_n1199));
  AOI21_X1  g773(.A(KEYINPUT127), .B1(new_n1198), .B2(new_n918), .ZN(new_n1200));
  NOR2_X1   g774(.A1(new_n1199), .A2(new_n1200), .ZN(G308));
  NAND2_X1  g775(.A1(new_n1198), .A2(new_n918), .ZN(G225));
endmodule


