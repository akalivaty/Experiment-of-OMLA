//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 0 1 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050;
  INV_X1    g000(.A(KEYINPUT16), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(G125), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n189), .B1(new_n193), .B2(new_n187), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  OAI211_X1 g010(.A(G146), .B(new_n189), .C1(new_n193), .C2(new_n187), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n199));
  INV_X1    g013(.A(G119), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(G128), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT23), .A3(G119), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n201), .B(new_n203), .C1(G119), .C2(new_n202), .ZN(new_n204));
  XNOR2_X1  g018(.A(G119), .B(G128), .ZN(new_n205));
  XOR2_X1   g019(.A(KEYINPUT24), .B(G110), .Z(new_n206));
  AOI22_X1  g020(.A1(new_n204), .A2(G110), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n198), .A2(new_n207), .ZN(new_n208));
  OAI22_X1  g022(.A1(new_n204), .A2(G110), .B1(new_n205), .B2(new_n206), .ZN(new_n209));
  AND2_X1   g023(.A1(new_n190), .A2(new_n192), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(new_n195), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n209), .A2(new_n197), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT22), .B(G137), .ZN(new_n214));
  INV_X1    g028(.A(G953), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(G221), .A3(G234), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n214), .B(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G902), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n208), .A2(new_n212), .A3(new_n217), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  OR2_X1    g036(.A1(new_n222), .A2(KEYINPUT25), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(KEYINPUT25), .ZN(new_n224));
  NAND2_X1  g038(.A1(G217), .A2(G902), .ZN(new_n225));
  INV_X1    g039(.A(G217), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(G234), .ZN(new_n227));
  XNOR2_X1  g041(.A(new_n227), .B(KEYINPUT74), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n223), .A2(new_n224), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT75), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n223), .A2(KEYINPUT75), .A3(new_n224), .A4(new_n228), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n219), .A2(new_n221), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n228), .A2(G902), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n231), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT73), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n195), .A2(G143), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n202), .B1(new_n239), .B2(KEYINPUT1), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G143), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT64), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT64), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G143), .ZN(new_n245));
  AOI21_X1  g059(.A(G146), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n195), .A2(G143), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n241), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT66), .ZN(new_n249));
  INV_X1    g063(.A(new_n239), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT64), .B(G143), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n250), .B1(new_n251), .B2(G146), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n249), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n243), .A2(new_n245), .A3(G146), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n255), .A2(new_n249), .A3(new_n239), .A4(new_n253), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n248), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT11), .ZN(new_n259));
  INV_X1    g073(.A(G134), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n259), .B1(new_n260), .B2(G137), .ZN(new_n261));
  INV_X1    g075(.A(G137), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(KEYINPUT11), .A3(G134), .ZN(new_n263));
  INV_X1    g077(.A(G131), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n260), .A2(G137), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n261), .A2(new_n263), .A3(new_n264), .A4(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n260), .A2(G137), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n262), .A2(G134), .ZN(new_n268));
  OAI21_X1  g082(.A(G131), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n258), .A2(new_n271), .ZN(new_n272));
  OR2_X1    g086(.A1(KEYINPUT69), .A2(G116), .ZN(new_n273));
  NAND2_X1  g087(.A1(KEYINPUT69), .A2(G116), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n273), .A2(G119), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT68), .ZN(new_n276));
  INV_X1    g090(.A(G116), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n276), .B1(new_n277), .B2(G119), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n200), .A2(KEYINPUT68), .A3(G116), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n275), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT2), .ZN(new_n281));
  INV_X1    g095(.A(G113), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n282), .A3(KEYINPUT67), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT67), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n284), .B1(KEYINPUT2), .B2(G113), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(KEYINPUT2), .A2(G113), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n280), .A2(new_n288), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n278), .A2(new_n279), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n290), .A2(new_n286), .A3(new_n287), .A4(new_n275), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  AND2_X1   g107(.A1(KEYINPUT0), .A2(G128), .ZN(new_n294));
  NOR2_X1   g108(.A1(KEYINPUT0), .A2(G128), .ZN(new_n295));
  OR2_X1    g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n244), .A2(G143), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n242), .A2(KEYINPUT64), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n195), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n247), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n296), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n255), .A2(new_n239), .A3(new_n294), .ZN(new_n302));
  OAI21_X1  g116(.A(KEYINPUT70), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n261), .A2(new_n263), .A3(new_n265), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G131), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n266), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n294), .A2(new_n295), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n307), .B1(new_n246), .B2(new_n247), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT70), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n255), .A2(new_n239), .A3(new_n294), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n303), .A2(new_n306), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n272), .A2(new_n293), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT28), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(KEYINPUT71), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT71), .B1(new_n313), .B2(new_n314), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G237), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(new_n215), .A3(G210), .ZN(new_n320));
  XOR2_X1   g134(.A(new_n320), .B(KEYINPUT27), .Z(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT26), .B(G101), .ZN(new_n322));
  XOR2_X1   g136(.A(new_n321), .B(new_n322), .Z(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT29), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AND3_X1   g140(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n309), .B1(new_n308), .B2(new_n310), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n305), .A2(new_n266), .ZN(new_n329));
  NOR3_X1   g143(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n255), .A2(new_n239), .A3(new_n253), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT66), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n256), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n270), .B1(new_n333), .B2(new_n248), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n292), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n313), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT72), .B1(new_n336), .B2(KEYINPUT28), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT72), .ZN(new_n338));
  AOI211_X1 g152(.A(new_n338), .B(new_n314), .C1(new_n335), .C2(new_n313), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n318), .B(new_n326), .C1(new_n337), .C2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n238), .B1(new_n340), .B2(new_n220), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n238), .A3(new_n220), .ZN(new_n343));
  INV_X1    g157(.A(new_n313), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT65), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n270), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n266), .A2(new_n269), .A3(KEYINPUT65), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n258), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n306), .A2(new_n310), .A3(new_n308), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n293), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT28), .B1(new_n344), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n318), .A2(new_n351), .A3(new_n323), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT30), .B1(new_n330), .B2(new_n334), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT30), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n240), .B1(new_n299), .B2(new_n300), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n355), .B1(new_n332), .B2(new_n256), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n346), .A2(new_n347), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n354), .B(new_n349), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n293), .B1(new_n353), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n324), .B1(new_n359), .B2(new_n344), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n352), .A2(new_n325), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n342), .A2(new_n343), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G472), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n354), .B1(new_n272), .B2(new_n312), .ZN(new_n364));
  INV_X1    g178(.A(new_n358), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n292), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(new_n313), .A3(new_n323), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT31), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n366), .A2(KEYINPUT31), .A3(new_n313), .A4(new_n323), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n313), .A2(new_n314), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT71), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n351), .A2(new_n373), .A3(new_n315), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n369), .A2(new_n370), .B1(new_n374), .B2(new_n324), .ZN(new_n375));
  NOR2_X1   g189(.A1(G472), .A2(G902), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT32), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n374), .A2(new_n324), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n353), .A2(new_n358), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n344), .B1(new_n380), .B2(new_n292), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT31), .B1(new_n381), .B2(new_n323), .ZN(new_n382));
  INV_X1    g196(.A(new_n370), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n379), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT32), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(new_n376), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n378), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n237), .B1(new_n363), .B2(new_n387), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n319), .A2(new_n215), .A3(G143), .A4(G214), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n243), .A2(new_n245), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n319), .A2(new_n215), .A3(G214), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G131), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT17), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n319), .A2(new_n215), .A3(G214), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n251), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(new_n264), .A3(new_n389), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n393), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n264), .B1(new_n396), .B2(new_n389), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT17), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n398), .A2(new_n196), .A3(new_n400), .A4(new_n197), .ZN(new_n401));
  XNOR2_X1  g215(.A(G113), .B(G122), .ZN(new_n402));
  INV_X1    g216(.A(G104), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n402), .B(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT18), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n396), .B(new_n389), .C1(new_n405), .C2(new_n264), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n193), .A2(G146), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n211), .A2(new_n407), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n406), .B(new_n408), .C1(new_n393), .C2(new_n405), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n401), .A2(new_n404), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n398), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n196), .B(new_n197), .C1(new_n393), .C2(new_n394), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT86), .ZN(new_n414));
  INV_X1    g228(.A(new_n404), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n414), .B1(new_n413), .B2(new_n415), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n410), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n220), .ZN(new_n420));
  INV_X1    g234(.A(new_n397), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(new_n399), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n193), .B(KEYINPUT19), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n197), .B1(new_n423), .B2(G146), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n409), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n415), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n410), .ZN(new_n427));
  INV_X1    g241(.A(G475), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n428), .A3(new_n220), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT20), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT20), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n427), .A2(new_n431), .A3(new_n428), .A4(new_n220), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n420), .A2(G475), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(G234), .A2(G237), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(G952), .A3(new_n215), .ZN(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(G898), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(G902), .A3(G953), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n435), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(KEYINPUT90), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n433), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT87), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n242), .A2(G128), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n443), .B1(new_n251), .B2(G128), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n260), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n273), .A2(G122), .A3(new_n274), .ZN(new_n446));
  INV_X1    g260(.A(G107), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n277), .A2(G122), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n446), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n447), .B1(new_n446), .B2(new_n449), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n445), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT13), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n243), .A2(new_n245), .A3(new_n454), .A4(G128), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G134), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n456), .B1(KEYINPUT13), .B2(new_n444), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n442), .B1(new_n453), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n443), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n459), .B1(new_n390), .B2(new_n202), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G134), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n451), .B1(new_n461), .B2(new_n445), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT14), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n446), .A2(new_n463), .A3(new_n449), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n464), .B(G107), .C1(new_n463), .C2(new_n446), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g280(.A(G134), .B(new_n455), .C1(new_n460), .C2(new_n454), .ZN(new_n467));
  INV_X1    g281(.A(new_n274), .ZN(new_n468));
  NOR2_X1   g282(.A1(KEYINPUT69), .A2(G116), .ZN(new_n469));
  INV_X1    g283(.A(G122), .ZN(new_n470));
  NOR3_X1   g284(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(G107), .B1(new_n471), .B2(new_n448), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n450), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n467), .A2(new_n473), .A3(KEYINPUT87), .A4(new_n445), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT9), .B(G234), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n475), .A2(new_n226), .A3(G953), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n458), .A2(new_n466), .A3(new_n474), .A4(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT88), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n467), .A2(new_n473), .A3(new_n445), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n480), .A2(new_n442), .B1(new_n462), .B2(new_n465), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n481), .A2(KEYINPUT88), .A3(new_n474), .A4(new_n476), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n458), .A2(new_n466), .A3(new_n474), .ZN(new_n483));
  INV_X1    g297(.A(new_n476), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n479), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n220), .ZN(new_n487));
  INV_X1    g301(.A(G478), .ZN(new_n488));
  NOR2_X1   g302(.A1(KEYINPUT89), .A2(KEYINPUT15), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(KEYINPUT89), .A2(KEYINPUT15), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n487), .B(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n441), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(G221), .B1(new_n475), .B2(G902), .ZN(new_n495));
  XOR2_X1   g309(.A(new_n495), .B(KEYINPUT76), .Z(new_n496));
  XNOR2_X1  g310(.A(G110), .B(G140), .ZN(new_n497));
  INV_X1    g311(.A(G227), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n498), .A2(G953), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n497), .B(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n202), .B1(new_n299), .B2(KEYINPUT1), .ZN(new_n502));
  OAI22_X1  g316(.A1(new_n254), .A2(new_n257), .B1(new_n252), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n447), .A2(G104), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n403), .A2(G107), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT77), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT3), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n504), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n447), .A2(G104), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT3), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n510), .A2(KEYINPUT77), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n506), .A2(KEYINPUT3), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G101), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n508), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(G101), .B1(new_n505), .B2(new_n504), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n503), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n356), .A2(new_n517), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(KEYINPUT12), .B1(new_n521), .B2(new_n306), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT12), .ZN(new_n523));
  AOI211_X1 g337(.A(new_n523), .B(new_n329), .C1(new_n519), .C2(new_n520), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT10), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n503), .A2(new_n526), .A3(new_n518), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT10), .B1(new_n356), .B2(new_n517), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n510), .A2(KEYINPUT77), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n505), .B1(new_n507), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n403), .A2(G107), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n532), .B1(new_n511), .B2(new_n509), .ZN(new_n533));
  OAI21_X1  g347(.A(G101), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(new_n515), .A3(KEYINPUT4), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT4), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n536), .B(G101), .C1(new_n531), .C2(new_n533), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n327), .A2(new_n328), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT78), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n303), .A2(new_n535), .A3(new_n311), .A4(new_n537), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT78), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n329), .B(new_n529), .C1(new_n540), .C2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n501), .B1(new_n525), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n529), .B1(new_n540), .B2(new_n543), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n546), .A2(new_n306), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n544), .A2(new_n501), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(G469), .B1(new_n550), .B2(G902), .ZN(new_n551));
  INV_X1    g365(.A(G469), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT79), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n544), .A2(new_n553), .A3(new_n501), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n553), .B1(new_n544), .B2(new_n501), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n522), .A2(new_n524), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n546), .A2(new_n306), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n501), .B1(new_n558), .B2(new_n544), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n552), .B(new_n220), .C1(new_n557), .C2(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n496), .B1(new_n551), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(G214), .B1(G237), .B2(G902), .ZN(new_n562));
  XOR2_X1   g376(.A(new_n562), .B(KEYINPUT80), .Z(new_n563));
  OAI21_X1  g377(.A(G210), .B1(G237), .B2(G902), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(KEYINPUT85), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n535), .A2(new_n292), .A3(new_n537), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n277), .A2(G119), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT5), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n282), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(new_n280), .B2(new_n568), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n570), .A2(new_n291), .A3(new_n515), .A4(new_n516), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(G110), .B(G122), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n566), .A2(new_n573), .A3(new_n571), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(KEYINPUT6), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT6), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n572), .A2(new_n578), .A3(new_n574), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n191), .B(new_n248), .C1(new_n254), .C2(new_n257), .ZN(new_n580));
  OAI21_X1  g394(.A(G125), .B1(new_n301), .B2(new_n302), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(G224), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(G953), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n584), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n580), .A2(new_n581), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n577), .A2(new_n579), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n220), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n586), .A2(KEYINPUT7), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n580), .A2(new_n581), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT84), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n582), .A2(new_n591), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT84), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n580), .A2(new_n596), .A3(new_n581), .A4(new_n592), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n594), .A2(new_n595), .A3(new_n597), .A4(new_n576), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT82), .B1(new_n517), .B2(KEYINPUT81), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n570), .A2(new_n291), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT82), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n515), .A2(new_n601), .A3(new_n516), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n573), .B(KEYINPUT8), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n604), .B1(new_n599), .B2(new_n600), .ZN(new_n605));
  OAI21_X1  g419(.A(KEYINPUT83), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  OR2_X1    g420(.A1(new_n599), .A2(new_n600), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT83), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n607), .A2(new_n608), .A3(new_n609), .A4(new_n604), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n598), .B1(new_n606), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n565), .B1(new_n590), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n606), .A2(new_n610), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n594), .A2(new_n576), .A3(new_n595), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n613), .A2(new_n597), .A3(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n565), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n615), .A2(new_n220), .A3(new_n616), .A4(new_n589), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n563), .B1(new_n612), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n388), .A2(new_n494), .A3(new_n561), .A4(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G101), .ZN(G3));
  NAND2_X1  g434(.A1(new_n384), .A2(new_n220), .ZN(new_n621));
  AOI22_X1  g435(.A1(new_n621), .A2(G472), .B1(new_n384), .B2(new_n376), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n561), .A2(new_n236), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n562), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(new_n612), .B2(new_n617), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n626), .B1(new_n483), .B2(new_n484), .ZN(new_n627));
  AOI22_X1  g441(.A1(new_n486), .A2(new_n626), .B1(new_n477), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n488), .A2(G902), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(G478), .B1(new_n486), .B2(new_n220), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n410), .ZN(new_n633));
  INV_X1    g447(.A(new_n418), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n633), .B1(new_n634), .B2(new_n416), .ZN(new_n635));
  OAI21_X1  g449(.A(G475), .B1(new_n635), .B2(G902), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n430), .A2(new_n432), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n630), .A2(new_n632), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT91), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n625), .A2(new_n638), .A3(new_n639), .A4(new_n440), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n625), .A2(new_n638), .A3(new_n440), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(KEYINPUT91), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n623), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(new_n403), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT92), .B(KEYINPUT34), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  NAND2_X1  g460(.A1(new_n612), .A2(new_n617), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n562), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n493), .A2(new_n433), .ZN(new_n649));
  INV_X1    g463(.A(new_n440), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n623), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT35), .B(G107), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  NOR2_X1   g469(.A1(new_n218), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n213), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n234), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT93), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n231), .A2(new_n659), .A3(new_n232), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n494), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n662), .A2(new_n561), .A3(new_n618), .A4(new_n622), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT37), .B(G110), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G12));
  AND3_X1   g479(.A1(new_n231), .A2(new_n659), .A3(new_n232), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n648), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n551), .A2(new_n560), .ZN(new_n668));
  INV_X1    g482(.A(new_n496), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n343), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n352), .A2(new_n325), .A3(new_n360), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n671), .A2(new_n341), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(G472), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n387), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n435), .B(KEYINPUT94), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n676), .B1(G900), .B2(new_n438), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n677), .B(KEYINPUT95), .Z(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n493), .A2(new_n433), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n670), .A2(new_n675), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  XOR2_X1   g497(.A(new_n678), .B(KEYINPUT39), .Z(new_n684));
  NAND2_X1  g498(.A1(new_n561), .A2(new_n684), .ZN(new_n685));
  OR2_X1    g499(.A1(new_n685), .A2(KEYINPUT40), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(KEYINPUT40), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n688), .B(KEYINPUT96), .Z(new_n689));
  AND3_X1   g503(.A1(new_n612), .A2(new_n617), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n689), .B1(new_n612), .B2(new_n617), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n636), .A2(new_n637), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n493), .A2(new_n693), .ZN(new_n694));
  NOR4_X1   g508(.A1(new_n692), .A2(new_n624), .A3(new_n660), .A4(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n686), .A2(new_n687), .A3(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT100), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT99), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n336), .A2(new_n324), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n367), .A2(KEYINPUT98), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n220), .ZN(new_n701));
  AOI21_X1  g515(.A(KEYINPUT98), .B1(new_n367), .B2(new_n699), .ZN(new_n702));
  OAI21_X1  g516(.A(G472), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n387), .A2(new_n698), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n698), .B1(new_n387), .B2(new_n703), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n697), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n375), .A2(KEYINPUT32), .A3(new_n377), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n385), .B1(new_n384), .B2(new_n376), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n703), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT99), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n387), .A2(new_n698), .A3(new_n703), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(KEYINPUT100), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n706), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n696), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(new_n251), .ZN(G45));
  AOI21_X1  g529(.A(new_n631), .B1(new_n628), .B2(new_n629), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n716), .A2(new_n433), .A3(new_n678), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n670), .A2(new_n675), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G146), .ZN(G48));
  NAND2_X1  g533(.A1(new_n642), .A2(new_n640), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n556), .B1(new_n548), .B2(KEYINPUT79), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n544), .A2(new_n553), .A3(new_n501), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n559), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(G469), .B1(new_n723), .B2(G902), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n724), .A2(new_n669), .A3(new_n560), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n720), .A2(new_n675), .A3(new_n236), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT41), .B(G113), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G15));
  NAND4_X1  g542(.A1(new_n675), .A2(new_n236), .A3(new_n651), .A4(new_n725), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G116), .ZN(G18));
  NAND4_X1  g544(.A1(new_n724), .A2(new_n560), .A3(new_n669), .A4(new_n625), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n675), .A2(new_n662), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G119), .ZN(G21));
  NAND3_X1  g548(.A1(new_n724), .A2(new_n560), .A3(new_n669), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n625), .A2(new_n493), .A3(new_n693), .A4(new_n440), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n369), .A2(new_n370), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n373), .A2(new_n315), .ZN(new_n739));
  INV_X1    g553(.A(new_n337), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n336), .A2(KEYINPUT72), .A3(KEYINPUT28), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n738), .B1(new_n742), .B2(new_n323), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n376), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT101), .B(G472), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n745), .B1(new_n375), .B2(G902), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n744), .A2(new_n236), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n737), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(KEYINPUT102), .B(G122), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G24));
  AOI22_X1  g565(.A1(new_n621), .A2(new_n745), .B1(new_n743), .B2(new_n376), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n660), .A3(new_n717), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n731), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n191), .ZN(G27));
  NAND3_X1  g569(.A1(new_n551), .A2(new_n560), .A3(KEYINPUT103), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT103), .B1(new_n551), .B2(new_n560), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n647), .A2(new_n624), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n669), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n388), .A3(new_n717), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT42), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n761), .A2(new_n388), .A3(KEYINPUT42), .A4(new_n717), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XOR2_X1   g580(.A(KEYINPUT104), .B(G131), .Z(new_n767));
  XNOR2_X1  g581(.A(new_n766), .B(new_n767), .ZN(G33));
  NAND3_X1  g582(.A1(new_n761), .A2(new_n388), .A3(new_n681), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G134), .ZN(G36));
  INV_X1    g584(.A(new_n759), .ZN(new_n771));
  OAI21_X1  g585(.A(KEYINPUT43), .B1(new_n716), .B2(new_n693), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n630), .A2(new_n632), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT43), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n774), .A3(new_n433), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n622), .A2(new_n776), .A3(new_n666), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n771), .B1(new_n777), .B2(KEYINPUT44), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n778), .B1(KEYINPUT44), .B2(new_n777), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n780), .B1(new_n545), .B2(new_n549), .ZN(new_n781));
  INV_X1    g595(.A(new_n544), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n500), .B1(new_n782), .B2(new_n556), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n783), .B(KEYINPUT45), .C1(new_n547), .C2(new_n548), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n781), .A2(new_n784), .A3(G469), .ZN(new_n785));
  NAND2_X1  g599(.A1(G469), .A2(G902), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT46), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n785), .A2(KEYINPUT46), .A3(new_n786), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n560), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n669), .A3(new_n684), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n779), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(new_n262), .ZN(G39));
  XNOR2_X1  g608(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n560), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n797), .B1(new_n787), .B2(new_n788), .ZN(new_n798));
  AOI211_X1 g612(.A(new_n496), .B(new_n796), .C1(new_n798), .C2(new_n790), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n795), .B1(new_n791), .B2(new_n669), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n341), .A2(new_n672), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n674), .B1(new_n802), .B2(new_n343), .ZN(new_n803));
  INV_X1    g617(.A(new_n387), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n805), .A2(new_n237), .A3(new_n717), .A4(new_n759), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n801), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(new_n188), .ZN(G42));
  INV_X1    g622(.A(KEYINPUT51), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n724), .A2(new_n560), .ZN(new_n810));
  XOR2_X1   g624(.A(new_n810), .B(KEYINPUT106), .Z(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n496), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT117), .B1(new_n801), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n676), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n772), .A2(new_n775), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n747), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n759), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT112), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT112), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n816), .A2(new_n819), .A3(new_n759), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n813), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n801), .A2(KEYINPUT117), .A3(new_n812), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n809), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n690), .A2(new_n691), .A3(new_n562), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n725), .A2(KEYINPUT113), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT113), .ZN(new_n827));
  INV_X1    g641(.A(new_n689), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n647), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n612), .A2(new_n617), .A3(new_n689), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(new_n624), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n827), .B1(new_n735), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n826), .A2(new_n832), .A3(new_n816), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT50), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n826), .A2(new_n832), .A3(new_n816), .A4(KEYINPUT50), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n835), .A2(KEYINPUT114), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT114), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n833), .A2(new_n838), .A3(new_n834), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n725), .A2(new_n759), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n815), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n752), .A2(new_n660), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n237), .A2(new_n435), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n725), .A2(new_n759), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n773), .A2(new_n693), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n704), .A2(new_n705), .A3(new_n697), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT100), .B1(new_n710), .B2(new_n711), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n846), .B(new_n847), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n837), .A2(new_n839), .A3(new_n843), .A4(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n841), .A2(new_n388), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n853), .A2(KEYINPUT48), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(KEYINPUT48), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n845), .B1(new_n706), .B2(new_n712), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n638), .ZN(new_n858));
  INV_X1    g672(.A(G952), .ZN(new_n859));
  AOI211_X1 g673(.A(new_n859), .B(G953), .C1(new_n816), .C2(new_n732), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n856), .A2(KEYINPUT118), .A3(new_n858), .A4(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n860), .B1(new_n854), .B2(new_n855), .ZN(new_n863));
  INV_X1    g677(.A(new_n858), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n824), .A2(new_n852), .B1(new_n861), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT116), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n821), .B1(new_n801), .B2(new_n812), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n868), .B1(new_n851), .B2(KEYINPUT115), .ZN(new_n869));
  AOI22_X1  g683(.A1(new_n857), .A2(new_n847), .B1(new_n842), .B2(new_n841), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT115), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n870), .A2(new_n871), .A3(new_n837), .A4(new_n839), .ZN(new_n872));
  AOI211_X1 g686(.A(new_n867), .B(KEYINPUT51), .C1(new_n869), .C2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n850), .A2(new_n839), .A3(new_n843), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n835), .A2(KEYINPUT114), .A3(new_n836), .ZN(new_n875));
  OAI21_X1  g689(.A(KEYINPUT115), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n868), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n876), .A2(new_n872), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT116), .B1(new_n878), .B2(new_n809), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n866), .B1(new_n873), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT119), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT119), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n866), .B(new_n882), .C1(new_n873), .C2(new_n879), .ZN(new_n883));
  INV_X1    g697(.A(new_n492), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n487), .B(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT109), .B1(new_n885), .B2(new_n693), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT109), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n493), .A2(new_n887), .A3(new_n433), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n886), .A2(new_n888), .A3(new_n440), .A4(new_n618), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n618), .A2(new_n440), .ZN(new_n890));
  AOI22_X1  g704(.A1(new_n889), .A2(KEYINPUT110), .B1(new_n890), .B2(new_n638), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT110), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n890), .A2(new_n892), .A3(new_n886), .A4(new_n888), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n619), .B(new_n663), .C1(new_n894), .C2(new_n623), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n726), .A2(new_n729), .A3(new_n733), .A4(new_n749), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(KEYINPUT108), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n661), .B1(new_n363), .B2(new_n387), .ZN(new_n898));
  AOI22_X1  g712(.A1(new_n898), .A2(new_n732), .B1(new_n748), .B2(new_n737), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT108), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n899), .A2(new_n900), .A3(new_n726), .A4(new_n729), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n895), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  NOR4_X1   g716(.A1(new_n666), .A2(new_n493), .A3(new_n693), .A4(new_n678), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n675), .A2(new_n561), .A3(new_n759), .A4(new_n903), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n752), .A2(new_n660), .A3(new_n717), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n761), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n769), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n764), .B2(new_n765), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT52), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n905), .A2(new_n732), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n682), .A2(new_n718), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n679), .A2(new_n669), .ZN(new_n912));
  NOR4_X1   g726(.A1(new_n648), .A2(new_n694), .A3(new_n660), .A4(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n758), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n914), .A3(new_n756), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n915), .B1(new_n711), .B2(new_n710), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n909), .B1(new_n911), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n680), .B1(new_n363), .B2(new_n387), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n754), .B1(new_n670), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n757), .A2(new_n758), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n920), .B(new_n913), .C1(new_n704), .C2(new_n705), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n919), .A2(new_n921), .A3(KEYINPUT52), .A4(new_n718), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n917), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n902), .A2(new_n908), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(KEYINPUT53), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n919), .A2(new_n921), .A3(new_n718), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT111), .ZN(new_n927));
  AOI22_X1  g741(.A1(new_n917), .A2(new_n922), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n926), .A2(new_n927), .A3(KEYINPUT52), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT53), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n902), .A2(new_n932), .A3(new_n908), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n925), .B(KEYINPUT54), .C1(new_n931), .C2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n924), .A2(new_n932), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n236), .B1(new_n803), .B2(new_n804), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n561), .A2(new_n494), .A3(new_n618), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n663), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n623), .B1(new_n891), .B2(new_n893), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n938), .A2(new_n939), .A3(new_n932), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n769), .A2(new_n904), .A3(new_n906), .ZN(new_n941));
  INV_X1    g755(.A(new_n896), .ZN(new_n942));
  AND4_X1   g756(.A1(new_n766), .A2(new_n940), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n943), .B1(new_n928), .B2(new_n930), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT54), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n935), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n934), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n881), .A2(new_n883), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n859), .A2(new_n215), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n773), .A2(new_n433), .ZN(new_n951));
  NOR4_X1   g765(.A1(new_n237), .A2(new_n951), .A3(new_n496), .A4(new_n563), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT49), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n952), .B1(new_n811), .B2(new_n953), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT107), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n811), .A2(new_n953), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n955), .A2(new_n713), .A3(new_n692), .A4(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n950), .A2(new_n957), .ZN(G75));
  NOR2_X1   g772(.A1(new_n215), .A2(G952), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n220), .B1(new_n935), .B2(new_n944), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT56), .B1(new_n961), .B2(new_n565), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n577), .A2(new_n579), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(new_n588), .ZN(new_n964));
  XNOR2_X1  g778(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n964), .B(new_n965), .Z(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n960), .B1(new_n962), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n962), .B2(new_n967), .ZN(G51));
  INV_X1    g783(.A(KEYINPUT121), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n946), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n935), .A2(new_n944), .A3(KEYINPUT121), .A4(new_n945), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n935), .A2(new_n944), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(KEYINPUT54), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n971), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n786), .B(KEYINPUT57), .Z(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n723), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n785), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n961), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n959), .B1(new_n979), .B2(new_n981), .ZN(G54));
  AND2_X1   g796(.A1(KEYINPUT58), .A2(G475), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n961), .A2(new_n427), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n427), .B1(new_n961), .B2(new_n983), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n984), .A2(new_n985), .A3(new_n959), .ZN(G60));
  NAND2_X1  g800(.A1(G478), .A2(G902), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT59), .Z(new_n988));
  AOI21_X1  g802(.A(new_n988), .B1(new_n934), .B2(new_n946), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n960), .B1(new_n989), .B2(new_n628), .ZN(new_n990));
  INV_X1    g804(.A(new_n988), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n628), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n990), .B1(new_n975), .B2(new_n992), .ZN(G63));
  XNOR2_X1  g807(.A(new_n225), .B(KEYINPUT60), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n994), .B1(new_n935), .B2(new_n944), .ZN(new_n995));
  OR2_X1    g809(.A1(new_n995), .A2(new_n233), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n657), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n996), .A2(new_n960), .A3(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT61), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n996), .A2(KEYINPUT61), .A3(new_n960), .A4(new_n997), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(G66));
  NOR2_X1   g816(.A1(new_n902), .A2(G953), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT122), .Z(new_n1004));
  OAI21_X1  g818(.A(G953), .B1(new_n436), .B2(new_n583), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT123), .Z(new_n1006));
  NAND2_X1  g820(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n963), .B1(G898), .B2(new_n215), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1007), .B(new_n1008), .ZN(G69));
  XOR2_X1   g823(.A(new_n380), .B(new_n423), .Z(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n638), .B1(new_n886), .B2(new_n888), .ZN(new_n1012));
  NOR4_X1   g826(.A1(new_n936), .A2(new_n685), .A3(new_n771), .A4(new_n1012), .ZN(new_n1013));
  NOR3_X1   g827(.A1(new_n807), .A2(new_n793), .A3(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(KEYINPUT62), .B1(new_n714), .B2(new_n911), .ZN(new_n1015));
  OR3_X1    g829(.A1(new_n714), .A2(KEYINPUT62), .A3(new_n911), .ZN(new_n1016));
  AND3_X1   g830(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1011), .B1(new_n1017), .B2(G953), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n215), .A2(G900), .ZN(new_n1019));
  INV_X1    g833(.A(new_n807), .ZN(new_n1020));
  NOR3_X1   g834(.A1(new_n936), .A2(new_n648), .A3(new_n694), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n1021), .A2(new_n669), .A3(new_n684), .A4(new_n791), .ZN(new_n1022));
  AND4_X1   g836(.A1(new_n766), .A2(new_n1020), .A3(new_n769), .A4(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n911), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1024), .B1(new_n792), .B2(new_n779), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1025), .B(KEYINPUT125), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1019), .B1(new_n1027), .B2(new_n215), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1018), .B1(new_n1028), .B2(new_n1011), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n215), .B1(G227), .B2(G900), .ZN(new_n1030));
  XOR2_X1   g844(.A(new_n1030), .B(KEYINPUT124), .Z(new_n1031));
  XNOR2_X1  g845(.A(new_n1029), .B(new_n1031), .ZN(G72));
  NOR2_X1   g846(.A1(new_n381), .A2(new_n324), .ZN(new_n1033));
  INV_X1    g847(.A(new_n1033), .ZN(new_n1034));
  NAND4_X1  g848(.A1(new_n1014), .A2(new_n1016), .A3(new_n902), .A4(new_n1015), .ZN(new_n1035));
  NAND2_X1  g849(.A1(G472), .A2(G902), .ZN(new_n1036));
  XOR2_X1   g850(.A(new_n1036), .B(KEYINPUT63), .Z(new_n1037));
  AOI21_X1  g851(.A(new_n1034), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  XOR2_X1   g852(.A(new_n1038), .B(KEYINPUT126), .Z(new_n1039));
  NAND2_X1  g853(.A1(new_n381), .A2(new_n324), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n1023), .A2(new_n1026), .A3(new_n902), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1041), .A2(new_n1037), .ZN(new_n1042));
  INV_X1    g856(.A(KEYINPUT127), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n1041), .A2(KEYINPUT127), .A3(new_n1037), .ZN(new_n1045));
  AOI21_X1  g859(.A(new_n1040), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g860(.A(new_n1037), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n1047), .B1(new_n360), .B2(new_n367), .ZN(new_n1048));
  OAI211_X1 g862(.A(new_n925), .B(new_n1048), .C1(new_n931), .C2(new_n933), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n1049), .A2(new_n960), .ZN(new_n1050));
  NOR3_X1   g864(.A1(new_n1039), .A2(new_n1046), .A3(new_n1050), .ZN(G57));
endmodule


