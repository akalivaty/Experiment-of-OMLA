

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U549 ( .A1(n532), .A2(G2104), .ZN(n995) );
  OR2_X2 U550 ( .A1(n523), .A2(n602), .ZN(n519) );
  NAND2_X2 U551 ( .A1(n703), .A2(n702), .ZN(n742) );
  NOR2_X1 U552 ( .A1(n778), .A2(n777), .ZN(n790) );
  XOR2_X1 U553 ( .A(G543), .B(KEYINPUT0), .Z(n602) );
  XNOR2_X1 U554 ( .A(KEYINPUT72), .B(n564), .ZN(n516) );
  AND2_X1 U555 ( .A1(n565), .A2(n516), .ZN(n517) );
  INV_X1 U556 ( .A(G168), .ZN(n719) );
  XNOR2_X1 U557 ( .A(n752), .B(KEYINPUT29), .ZN(n753) );
  INV_X1 U558 ( .A(KEYINPUT90), .ZN(n715) );
  AND2_X1 U559 ( .A1(n781), .A2(n776), .ZN(n777) );
  NOR2_X1 U560 ( .A1(G2104), .A2(G2105), .ZN(n536) );
  NOR2_X1 U561 ( .A1(n792), .A2(n791), .ZN(n794) );
  XOR2_X1 U562 ( .A(n569), .B(KEYINPUT15), .Z(n1009) );
  NOR2_X1 U563 ( .A1(G651), .A2(G543), .ZN(n629) );
  AND2_X1 U564 ( .A1(n563), .A2(n562), .ZN(n954) );
  NAND2_X1 U565 ( .A1(n629), .A2(G89), .ZN(n518) );
  XNOR2_X1 U566 ( .A(n518), .B(KEYINPUT4), .ZN(n521) );
  INV_X1 U567 ( .A(G651), .ZN(n523) );
  XOR2_X2 U568 ( .A(KEYINPUT66), .B(n519), .Z(n630) );
  NAND2_X1 U569 ( .A1(G76), .A2(n630), .ZN(n520) );
  NAND2_X1 U570 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U571 ( .A(n522), .B(KEYINPUT5), .ZN(n530) );
  NOR2_X1 U572 ( .A1(G543), .A2(n523), .ZN(n524) );
  XOR2_X1 U573 ( .A(KEYINPUT1), .B(n524), .Z(n634) );
  NAND2_X1 U574 ( .A1(G63), .A2(n634), .ZN(n527) );
  NOR2_X1 U575 ( .A1(G651), .A2(n602), .ZN(n525) );
  XNOR2_X2 U576 ( .A(KEYINPUT64), .B(n525), .ZN(n635) );
  NAND2_X1 U577 ( .A1(G51), .A2(n635), .ZN(n526) );
  NAND2_X1 U578 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U579 ( .A(KEYINPUT6), .B(n528), .Z(n529) );
  NAND2_X1 U580 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U581 ( .A(n531), .B(KEYINPUT7), .ZN(G168) );
  INV_X1 U582 ( .A(G2105), .ZN(n532) );
  NOR2_X1 U583 ( .A1(G2104), .A2(n532), .ZN(n992) );
  NAND2_X1 U584 ( .A1(n992), .A2(G125), .ZN(n535) );
  NAND2_X1 U585 ( .A1(G101), .A2(n995), .ZN(n533) );
  XOR2_X1 U586 ( .A(KEYINPUT23), .B(n533), .Z(n534) );
  NAND2_X1 U587 ( .A1(n535), .A2(n534), .ZN(n540) );
  XOR2_X1 U588 ( .A(KEYINPUT17), .B(n536), .Z(n996) );
  NAND2_X1 U589 ( .A1(G137), .A2(n996), .ZN(n538) );
  AND2_X1 U590 ( .A1(G2104), .A2(G2105), .ZN(n991) );
  NAND2_X1 U591 ( .A1(G113), .A2(n991), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U593 ( .A1(n540), .A2(n539), .ZN(G160) );
  XNOR2_X1 U594 ( .A(KEYINPUT82), .B(G44), .ZN(n541) );
  XNOR2_X1 U595 ( .A(n541), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U596 ( .A1(G64), .A2(n634), .ZN(n543) );
  NAND2_X1 U597 ( .A1(G52), .A2(n635), .ZN(n542) );
  NAND2_X1 U598 ( .A1(n543), .A2(n542), .ZN(n548) );
  NAND2_X1 U599 ( .A1(G90), .A2(n629), .ZN(n545) );
  NAND2_X1 U600 ( .A1(G77), .A2(n630), .ZN(n544) );
  NAND2_X1 U601 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U602 ( .A(KEYINPUT9), .B(n546), .Z(n547) );
  NOR2_X1 U603 ( .A1(n548), .A2(n547), .ZN(G171) );
  AND2_X1 U604 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U605 ( .A(G132), .ZN(G219) );
  INV_X1 U606 ( .A(G82), .ZN(G220) );
  INV_X1 U607 ( .A(G57), .ZN(G237) );
  NAND2_X1 U608 ( .A1(G7), .A2(G661), .ZN(n549) );
  XOR2_X1 U609 ( .A(n549), .B(KEYINPUT10), .Z(n824) );
  NAND2_X1 U610 ( .A1(n824), .A2(G567), .ZN(n550) );
  XOR2_X1 U611 ( .A(KEYINPUT11), .B(n550), .Z(G234) );
  NAND2_X1 U612 ( .A1(G68), .A2(n630), .ZN(n551) );
  XNOR2_X1 U613 ( .A(n551), .B(KEYINPUT68), .ZN(n555) );
  XOR2_X1 U614 ( .A(KEYINPUT12), .B(KEYINPUT67), .Z(n553) );
  NAND2_X1 U615 ( .A1(G81), .A2(n629), .ZN(n552) );
  XNOR2_X1 U616 ( .A(n553), .B(n552), .ZN(n554) );
  NAND2_X1 U617 ( .A1(n555), .A2(n554), .ZN(n557) );
  XNOR2_X1 U618 ( .A(KEYINPUT69), .B(KEYINPUT13), .ZN(n556) );
  XNOR2_X1 U619 ( .A(n557), .B(n556), .ZN(n560) );
  NAND2_X1 U620 ( .A1(n634), .A2(G56), .ZN(n558) );
  XOR2_X1 U621 ( .A(KEYINPUT14), .B(n558), .Z(n559) );
  NOR2_X1 U622 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U623 ( .A(n561), .B(KEYINPUT70), .ZN(n563) );
  NAND2_X1 U624 ( .A1(G43), .A2(n635), .ZN(n562) );
  XOR2_X1 U625 ( .A(G860), .B(KEYINPUT71), .Z(n581) );
  NAND2_X1 U626 ( .A1(n954), .A2(n581), .ZN(G153) );
  INV_X1 U627 ( .A(G171), .ZN(G301) );
  NAND2_X1 U628 ( .A1(G868), .A2(G301), .ZN(n571) );
  NAND2_X1 U629 ( .A1(n634), .A2(G66), .ZN(n568) );
  NAND2_X1 U630 ( .A1(G54), .A2(n635), .ZN(n566) );
  NAND2_X1 U631 ( .A1(G79), .A2(n630), .ZN(n565) );
  NAND2_X1 U632 ( .A1(G92), .A2(n629), .ZN(n564) );
  AND2_X1 U633 ( .A1(n566), .A2(n517), .ZN(n567) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  INV_X1 U635 ( .A(G868), .ZN(n648) );
  NAND2_X1 U636 ( .A1(n1009), .A2(n648), .ZN(n570) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(G284) );
  XOR2_X1 U638 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  AND2_X1 U639 ( .A1(n634), .A2(G65), .ZN(n575) );
  NAND2_X1 U640 ( .A1(G78), .A2(n630), .ZN(n573) );
  NAND2_X1 U641 ( .A1(G53), .A2(n635), .ZN(n572) );
  NAND2_X1 U642 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U643 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U644 ( .A1(n629), .A2(G91), .ZN(n576) );
  NAND2_X1 U645 ( .A1(n577), .A2(n576), .ZN(G299) );
  NOR2_X1 U646 ( .A1(G286), .A2(n648), .ZN(n579) );
  NOR2_X1 U647 ( .A1(G868), .A2(G299), .ZN(n578) );
  NOR2_X1 U648 ( .A1(n579), .A2(n578), .ZN(G297) );
  INV_X1 U649 ( .A(G559), .ZN(n580) );
  NOR2_X1 U650 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U651 ( .A1(n1009), .A2(n582), .ZN(n583) );
  XOR2_X1 U652 ( .A(KEYINPUT16), .B(n583), .Z(G148) );
  INV_X1 U653 ( .A(n954), .ZN(n584) );
  NOR2_X1 U654 ( .A1(G868), .A2(n584), .ZN(n587) );
  INV_X1 U655 ( .A(n1009), .ZN(n737) );
  NAND2_X1 U656 ( .A1(G868), .A2(n737), .ZN(n585) );
  NOR2_X1 U657 ( .A1(G559), .A2(n585), .ZN(n586) );
  NOR2_X1 U658 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U659 ( .A(KEYINPUT73), .B(n588), .Z(G282) );
  NAND2_X1 U660 ( .A1(n992), .A2(G123), .ZN(n589) );
  XNOR2_X1 U661 ( .A(n589), .B(KEYINPUT18), .ZN(n591) );
  NAND2_X1 U662 ( .A1(G135), .A2(n996), .ZN(n590) );
  NAND2_X1 U663 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U664 ( .A(KEYINPUT74), .B(n592), .ZN(n596) );
  NAND2_X1 U665 ( .A1(G99), .A2(n995), .ZN(n594) );
  NAND2_X1 U666 ( .A1(G111), .A2(n991), .ZN(n593) );
  NAND2_X1 U667 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U668 ( .A1(n596), .A2(n595), .ZN(n979) );
  XOR2_X1 U669 ( .A(G2096), .B(n979), .Z(n597) );
  NOR2_X1 U670 ( .A1(G2100), .A2(n597), .ZN(n598) );
  XNOR2_X1 U671 ( .A(KEYINPUT75), .B(n598), .ZN(G156) );
  NAND2_X1 U672 ( .A1(G651), .A2(G74), .ZN(n600) );
  NAND2_X1 U673 ( .A1(G49), .A2(n635), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U675 ( .A(KEYINPUT78), .B(n601), .Z(n606) );
  NAND2_X1 U676 ( .A1(G87), .A2(n602), .ZN(n603) );
  XNOR2_X1 U677 ( .A(KEYINPUT79), .B(n603), .ZN(n604) );
  NOR2_X1 U678 ( .A1(n634), .A2(n604), .ZN(n605) );
  NAND2_X1 U679 ( .A1(n606), .A2(n605), .ZN(G288) );
  NAND2_X1 U680 ( .A1(n634), .A2(G62), .ZN(n607) );
  XNOR2_X1 U681 ( .A(n607), .B(KEYINPUT80), .ZN(n609) );
  NAND2_X1 U682 ( .A1(G50), .A2(n635), .ZN(n608) );
  NAND2_X1 U683 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U684 ( .A(KEYINPUT81), .B(n610), .ZN(n614) );
  NAND2_X1 U685 ( .A1(n630), .A2(G75), .ZN(n612) );
  NAND2_X1 U686 ( .A1(G88), .A2(n629), .ZN(n611) );
  AND2_X1 U687 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U688 ( .A1(n614), .A2(n613), .ZN(G303) );
  INV_X1 U689 ( .A(G303), .ZN(G166) );
  NAND2_X1 U690 ( .A1(G86), .A2(n629), .ZN(n616) );
  NAND2_X1 U691 ( .A1(G61), .A2(n634), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U693 ( .A1(n630), .A2(G73), .ZN(n617) );
  XOR2_X1 U694 ( .A(KEYINPUT2), .B(n617), .Z(n618) );
  NOR2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n621) );
  NAND2_X1 U696 ( .A1(G48), .A2(n635), .ZN(n620) );
  NAND2_X1 U697 ( .A1(n621), .A2(n620), .ZN(G305) );
  NAND2_X1 U698 ( .A1(G60), .A2(n634), .ZN(n623) );
  NAND2_X1 U699 ( .A1(G72), .A2(n630), .ZN(n622) );
  NAND2_X1 U700 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U701 ( .A1(G85), .A2(n629), .ZN(n624) );
  XNOR2_X1 U702 ( .A(KEYINPUT65), .B(n624), .ZN(n625) );
  NOR2_X1 U703 ( .A1(n626), .A2(n625), .ZN(n628) );
  NAND2_X1 U704 ( .A1(G47), .A2(n635), .ZN(n627) );
  NAND2_X1 U705 ( .A1(n628), .A2(n627), .ZN(G290) );
  NAND2_X1 U706 ( .A1(n737), .A2(G559), .ZN(n953) );
  NAND2_X1 U707 ( .A1(G93), .A2(n629), .ZN(n632) );
  NAND2_X1 U708 ( .A1(G80), .A2(n630), .ZN(n631) );
  NAND2_X1 U709 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U710 ( .A(KEYINPUT76), .B(n633), .ZN(n639) );
  NAND2_X1 U711 ( .A1(G67), .A2(n634), .ZN(n637) );
  NAND2_X1 U712 ( .A1(G55), .A2(n635), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U714 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U715 ( .A(KEYINPUT77), .B(n640), .ZN(n956) );
  XNOR2_X1 U716 ( .A(KEYINPUT19), .B(G299), .ZN(n641) );
  XNOR2_X1 U717 ( .A(n641), .B(G288), .ZN(n642) );
  XOR2_X1 U718 ( .A(n956), .B(n642), .Z(n645) );
  XOR2_X1 U719 ( .A(G166), .B(G305), .Z(n643) );
  XNOR2_X1 U720 ( .A(n643), .B(G290), .ZN(n644) );
  XNOR2_X1 U721 ( .A(n645), .B(n644), .ZN(n646) );
  XOR2_X1 U722 ( .A(n954), .B(n646), .Z(n1007) );
  XNOR2_X1 U723 ( .A(n953), .B(n1007), .ZN(n647) );
  NAND2_X1 U724 ( .A1(n647), .A2(G868), .ZN(n650) );
  NAND2_X1 U725 ( .A1(n648), .A2(n956), .ZN(n649) );
  NAND2_X1 U726 ( .A1(n650), .A2(n649), .ZN(G295) );
  NAND2_X1 U727 ( .A1(G2084), .A2(G2078), .ZN(n651) );
  XOR2_X1 U728 ( .A(KEYINPUT20), .B(n651), .Z(n652) );
  NAND2_X1 U729 ( .A1(G2090), .A2(n652), .ZN(n653) );
  XNOR2_X1 U730 ( .A(KEYINPUT21), .B(n653), .ZN(n654) );
  NAND2_X1 U731 ( .A1(n654), .A2(G2072), .ZN(G158) );
  NAND2_X1 U732 ( .A1(G69), .A2(G120), .ZN(n655) );
  NOR2_X1 U733 ( .A1(G237), .A2(n655), .ZN(n656) );
  NAND2_X1 U734 ( .A1(G108), .A2(n656), .ZN(n951) );
  NAND2_X1 U735 ( .A1(G567), .A2(n951), .ZN(n657) );
  XNOR2_X1 U736 ( .A(n657), .B(KEYINPUT83), .ZN(n662) );
  NOR2_X1 U737 ( .A1(G220), .A2(G219), .ZN(n658) );
  XNOR2_X1 U738 ( .A(KEYINPUT22), .B(n658), .ZN(n659) );
  NAND2_X1 U739 ( .A1(n659), .A2(G96), .ZN(n660) );
  OR2_X1 U740 ( .A1(G218), .A2(n660), .ZN(n952) );
  AND2_X1 U741 ( .A1(G2106), .A2(n952), .ZN(n661) );
  NOR2_X1 U742 ( .A1(n662), .A2(n661), .ZN(G319) );
  INV_X1 U743 ( .A(G319), .ZN(n664) );
  NAND2_X1 U744 ( .A1(G483), .A2(G661), .ZN(n663) );
  NOR2_X1 U745 ( .A1(n664), .A2(n663), .ZN(n828) );
  NAND2_X1 U746 ( .A1(n828), .A2(G36), .ZN(G176) );
  NAND2_X1 U747 ( .A1(n995), .A2(G102), .ZN(n665) );
  XNOR2_X1 U748 ( .A(n665), .B(KEYINPUT84), .ZN(n667) );
  NAND2_X1 U749 ( .A1(G138), .A2(n996), .ZN(n666) );
  NAND2_X1 U750 ( .A1(n667), .A2(n666), .ZN(n671) );
  NAND2_X1 U751 ( .A1(G114), .A2(n991), .ZN(n669) );
  NAND2_X1 U752 ( .A1(G126), .A2(n992), .ZN(n668) );
  NAND2_X1 U753 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U754 ( .A1(n671), .A2(n670), .ZN(G164) );
  NAND2_X1 U755 ( .A1(G131), .A2(n996), .ZN(n673) );
  NAND2_X1 U756 ( .A1(G119), .A2(n992), .ZN(n672) );
  NAND2_X1 U757 ( .A1(n673), .A2(n672), .ZN(n677) );
  NAND2_X1 U758 ( .A1(G95), .A2(n995), .ZN(n675) );
  NAND2_X1 U759 ( .A1(G107), .A2(n991), .ZN(n674) );
  NAND2_X1 U760 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U761 ( .A1(n677), .A2(n676), .ZN(n983) );
  INV_X1 U762 ( .A(G1991), .ZN(n974) );
  NOR2_X1 U763 ( .A1(n983), .A2(n974), .ZN(n686) );
  NAND2_X1 U764 ( .A1(G141), .A2(n996), .ZN(n679) );
  NAND2_X1 U765 ( .A1(G129), .A2(n992), .ZN(n678) );
  NAND2_X1 U766 ( .A1(n679), .A2(n678), .ZN(n682) );
  NAND2_X1 U767 ( .A1(n995), .A2(G105), .ZN(n680) );
  XOR2_X1 U768 ( .A(KEYINPUT38), .B(n680), .Z(n681) );
  NOR2_X1 U769 ( .A1(n682), .A2(n681), .ZN(n684) );
  NAND2_X1 U770 ( .A1(n991), .A2(G117), .ZN(n683) );
  NAND2_X1 U771 ( .A1(n684), .A2(n683), .ZN(n984) );
  AND2_X1 U772 ( .A1(G1996), .A2(n984), .ZN(n685) );
  NOR2_X1 U773 ( .A1(n686), .A2(n685), .ZN(n931) );
  NOR2_X1 U774 ( .A1(G164), .A2(G1384), .ZN(n702) );
  INV_X1 U775 ( .A(n702), .ZN(n688) );
  NAND2_X1 U776 ( .A1(G40), .A2(G160), .ZN(n687) );
  XNOR2_X1 U777 ( .A(n687), .B(KEYINPUT85), .ZN(n703) );
  NAND2_X1 U778 ( .A1(n688), .A2(n703), .ZN(n689) );
  NOR2_X1 U779 ( .A1(n931), .A2(n689), .ZN(n797) );
  XNOR2_X1 U780 ( .A(KEYINPUT87), .B(n797), .ZN(n700) );
  INV_X1 U781 ( .A(n689), .ZN(n805) );
  XNOR2_X1 U782 ( .A(KEYINPUT86), .B(KEYINPUT34), .ZN(n693) );
  NAND2_X1 U783 ( .A1(G104), .A2(n995), .ZN(n691) );
  NAND2_X1 U784 ( .A1(G140), .A2(n996), .ZN(n690) );
  NAND2_X1 U785 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U786 ( .A(n693), .B(n692), .ZN(n698) );
  NAND2_X1 U787 ( .A1(G116), .A2(n991), .ZN(n695) );
  NAND2_X1 U788 ( .A1(G128), .A2(n992), .ZN(n694) );
  NAND2_X1 U789 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U790 ( .A(KEYINPUT35), .B(n696), .Z(n697) );
  NOR2_X1 U791 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U792 ( .A(KEYINPUT36), .B(n699), .ZN(n985) );
  XNOR2_X1 U793 ( .A(G2067), .B(KEYINPUT37), .ZN(n802) );
  NOR2_X1 U794 ( .A1(n985), .A2(n802), .ZN(n940) );
  NAND2_X1 U795 ( .A1(n805), .A2(n940), .ZN(n800) );
  NAND2_X1 U796 ( .A1(n700), .A2(n800), .ZN(n701) );
  XNOR2_X1 U797 ( .A(n701), .B(KEYINPUT88), .ZN(n792) );
  XOR2_X1 U798 ( .A(G1981), .B(G305), .Z(n884) );
  NAND2_X1 U799 ( .A1(G8), .A2(n742), .ZN(n786) );
  INV_X1 U800 ( .A(n786), .ZN(n705) );
  NAND2_X1 U801 ( .A1(G288), .A2(G1976), .ZN(n704) );
  XOR2_X1 U802 ( .A(KEYINPUT97), .B(n704), .Z(n898) );
  AND2_X1 U803 ( .A1(n705), .A2(n898), .ZN(n706) );
  NOR2_X1 U804 ( .A1(KEYINPUT33), .A2(n706), .ZN(n709) );
  NOR2_X1 U805 ( .A1(G1976), .A2(G288), .ZN(n774) );
  NAND2_X1 U806 ( .A1(n774), .A2(KEYINPUT33), .ZN(n707) );
  NOR2_X1 U807 ( .A1(n786), .A2(n707), .ZN(n708) );
  NOR2_X1 U808 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U809 ( .A1(n884), .A2(n710), .ZN(n778) );
  NOR2_X1 U810 ( .A1(G2090), .A2(n742), .ZN(n711) );
  XNOR2_X1 U811 ( .A(n711), .B(KEYINPUT96), .ZN(n713) );
  NOR2_X1 U812 ( .A1(n786), .A2(G1971), .ZN(n712) );
  NOR2_X1 U813 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U814 ( .A1(n714), .A2(G303), .ZN(n761) );
  NOR2_X1 U815 ( .A1(G2084), .A2(n742), .ZN(n764) );
  NOR2_X1 U816 ( .A1(G1966), .A2(n786), .ZN(n716) );
  XNOR2_X1 U817 ( .A(n716), .B(n715), .ZN(n766) );
  NAND2_X1 U818 ( .A1(n766), .A2(G8), .ZN(n717) );
  NOR2_X1 U819 ( .A1(n764), .A2(n717), .ZN(n718) );
  XNOR2_X1 U820 ( .A(n718), .B(KEYINPUT30), .ZN(n720) );
  AND2_X1 U821 ( .A1(n720), .A2(n719), .ZN(n724) );
  INV_X1 U822 ( .A(G1961), .ZN(n888) );
  NAND2_X1 U823 ( .A1(n742), .A2(n888), .ZN(n722) );
  INV_X1 U824 ( .A(n742), .ZN(n740) );
  XNOR2_X1 U825 ( .A(G2078), .B(KEYINPUT25), .ZN(n838) );
  NAND2_X1 U826 ( .A1(n740), .A2(n838), .ZN(n721) );
  NAND2_X1 U827 ( .A1(n722), .A2(n721), .ZN(n755) );
  NOR2_X1 U828 ( .A1(G171), .A2(n755), .ZN(n723) );
  NOR2_X1 U829 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U830 ( .A(KEYINPUT31), .B(n725), .Z(n759) );
  INV_X1 U831 ( .A(G1996), .ZN(n969) );
  NOR2_X1 U832 ( .A1(n742), .A2(n969), .ZN(n726) );
  XNOR2_X1 U833 ( .A(n726), .B(KEYINPUT26), .ZN(n728) );
  AND2_X1 U834 ( .A1(n742), .A2(G1341), .ZN(n727) );
  NOR2_X1 U835 ( .A1(n728), .A2(n727), .ZN(n735) );
  AND2_X1 U836 ( .A1(n735), .A2(n737), .ZN(n729) );
  NAND2_X1 U837 ( .A1(n729), .A2(n954), .ZN(n733) );
  NOR2_X1 U838 ( .A1(G2067), .A2(n742), .ZN(n731) );
  NOR2_X1 U839 ( .A1(n740), .A2(G1348), .ZN(n730) );
  NOR2_X1 U840 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U841 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U842 ( .A(n734), .B(KEYINPUT91), .ZN(n739) );
  AND2_X1 U843 ( .A1(n735), .A2(n954), .ZN(n736) );
  NOR2_X1 U844 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U845 ( .A1(n739), .A2(n738), .ZN(n746) );
  NAND2_X1 U846 ( .A1(n740), .A2(G2072), .ZN(n741) );
  XOR2_X1 U847 ( .A(KEYINPUT27), .B(n741), .Z(n744) );
  NAND2_X1 U848 ( .A1(G1956), .A2(n742), .ZN(n743) );
  NAND2_X1 U849 ( .A1(n744), .A2(n743), .ZN(n748) );
  NOR2_X1 U850 ( .A1(G299), .A2(n748), .ZN(n745) );
  NOR2_X1 U851 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U852 ( .A(n747), .B(KEYINPUT92), .ZN(n751) );
  NAND2_X1 U853 ( .A1(G299), .A2(n748), .ZN(n749) );
  XOR2_X1 U854 ( .A(n749), .B(KEYINPUT28), .Z(n750) );
  NOR2_X2 U855 ( .A1(n751), .A2(n750), .ZN(n754) );
  INV_X1 U856 ( .A(KEYINPUT93), .ZN(n752) );
  XNOR2_X1 U857 ( .A(n754), .B(n753), .ZN(n757) );
  NAND2_X1 U858 ( .A1(n755), .A2(G171), .ZN(n756) );
  NAND2_X1 U859 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U860 ( .A1(n759), .A2(n758), .ZN(n767) );
  NAND2_X1 U861 ( .A1(G286), .A2(n767), .ZN(n760) );
  NAND2_X1 U862 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U863 ( .A1(G8), .A2(n762), .ZN(n763) );
  XNOR2_X1 U864 ( .A(KEYINPUT32), .B(n763), .ZN(n772) );
  NAND2_X1 U865 ( .A1(G8), .A2(n764), .ZN(n765) );
  AND2_X1 U866 ( .A1(n766), .A2(n765), .ZN(n769) );
  XNOR2_X1 U867 ( .A(n767), .B(KEYINPUT94), .ZN(n768) );
  AND2_X1 U868 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U869 ( .A(n770), .B(KEYINPUT95), .ZN(n771) );
  NAND2_X1 U870 ( .A1(n772), .A2(n771), .ZN(n781) );
  NOR2_X1 U871 ( .A1(G1971), .A2(G303), .ZN(n773) );
  NOR2_X1 U872 ( .A1(n774), .A2(n773), .ZN(n894) );
  INV_X1 U873 ( .A(KEYINPUT33), .ZN(n775) );
  AND2_X1 U874 ( .A1(n894), .A2(n775), .ZN(n776) );
  NOR2_X1 U875 ( .A1(G2090), .A2(G303), .ZN(n779) );
  NAND2_X1 U876 ( .A1(G8), .A2(n779), .ZN(n780) );
  NAND2_X1 U877 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U878 ( .A1(n782), .A2(n786), .ZN(n788) );
  NOR2_X1 U879 ( .A1(G1981), .A2(G305), .ZN(n783) );
  XNOR2_X1 U880 ( .A(n783), .B(KEYINPUT24), .ZN(n784) );
  XNOR2_X1 U881 ( .A(KEYINPUT89), .B(n784), .ZN(n785) );
  OR2_X1 U882 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U883 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X1 U884 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U885 ( .A(G1986), .B(G290), .ZN(n890) );
  NAND2_X1 U886 ( .A1(n805), .A2(n890), .ZN(n793) );
  NAND2_X1 U887 ( .A1(n794), .A2(n793), .ZN(n809) );
  NOR2_X1 U888 ( .A1(G1996), .A2(n984), .ZN(n933) );
  NOR2_X1 U889 ( .A1(G1986), .A2(G290), .ZN(n795) );
  AND2_X1 U890 ( .A1(n974), .A2(n983), .ZN(n926) );
  NOR2_X1 U891 ( .A1(n795), .A2(n926), .ZN(n796) );
  NOR2_X1 U892 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U893 ( .A1(n933), .A2(n798), .ZN(n799) );
  XNOR2_X1 U894 ( .A(n799), .B(KEYINPUT39), .ZN(n801) );
  NAND2_X1 U895 ( .A1(n801), .A2(n800), .ZN(n803) );
  NAND2_X1 U896 ( .A1(n985), .A2(n802), .ZN(n927) );
  NAND2_X1 U897 ( .A1(n803), .A2(n927), .ZN(n804) );
  XNOR2_X1 U898 ( .A(KEYINPUT98), .B(n804), .ZN(n806) );
  NAND2_X1 U899 ( .A1(n806), .A2(n805), .ZN(n807) );
  XOR2_X1 U900 ( .A(KEYINPUT99), .B(n807), .Z(n808) );
  NAND2_X1 U901 ( .A1(n809), .A2(n808), .ZN(n811) );
  XNOR2_X1 U902 ( .A(KEYINPUT100), .B(KEYINPUT40), .ZN(n810) );
  XNOR2_X1 U903 ( .A(n811), .B(n810), .ZN(G329) );
  XNOR2_X1 U904 ( .A(G2443), .B(G1341), .ZN(n821) );
  XOR2_X1 U905 ( .A(G2451), .B(G2446), .Z(n813) );
  XNOR2_X1 U906 ( .A(G1348), .B(KEYINPUT101), .ZN(n812) );
  XNOR2_X1 U907 ( .A(n813), .B(n812), .ZN(n817) );
  XOR2_X1 U908 ( .A(G2435), .B(G2438), .Z(n815) );
  XNOR2_X1 U909 ( .A(G2454), .B(KEYINPUT102), .ZN(n814) );
  XNOR2_X1 U910 ( .A(n815), .B(n814), .ZN(n816) );
  XOR2_X1 U911 ( .A(n817), .B(n816), .Z(n819) );
  XNOR2_X1 U912 ( .A(G2427), .B(G2430), .ZN(n818) );
  XNOR2_X1 U913 ( .A(n819), .B(n818), .ZN(n820) );
  XNOR2_X1 U914 ( .A(n821), .B(n820), .ZN(n822) );
  NAND2_X1 U915 ( .A1(n822), .A2(G14), .ZN(n1012) );
  XNOR2_X1 U916 ( .A(KEYINPUT103), .B(n1012), .ZN(G401) );
  NAND2_X1 U917 ( .A1(n824), .A2(G2106), .ZN(n823) );
  XNOR2_X1 U918 ( .A(n823), .B(KEYINPUT104), .ZN(G217) );
  INV_X1 U919 ( .A(n824), .ZN(G223) );
  AND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n825) );
  NAND2_X1 U921 ( .A1(G661), .A2(n825), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n826) );
  XOR2_X1 U923 ( .A(KEYINPUT105), .B(n826), .Z(n827) );
  NAND2_X1 U924 ( .A1(n828), .A2(n827), .ZN(G188) );
  NAND2_X1 U926 ( .A1(G100), .A2(n995), .ZN(n830) );
  NAND2_X1 U927 ( .A1(G112), .A2(n991), .ZN(n829) );
  NAND2_X1 U928 ( .A1(n830), .A2(n829), .ZN(n831) );
  XNOR2_X1 U929 ( .A(KEYINPUT108), .B(n831), .ZN(n834) );
  NAND2_X1 U930 ( .A1(n992), .A2(G124), .ZN(n832) );
  XOR2_X1 U931 ( .A(KEYINPUT44), .B(n832), .Z(n833) );
  NOR2_X1 U932 ( .A1(n834), .A2(n833), .ZN(n836) );
  NAND2_X1 U933 ( .A1(n996), .A2(G136), .ZN(n835) );
  NAND2_X1 U934 ( .A1(n836), .A2(n835), .ZN(n837) );
  XNOR2_X1 U935 ( .A(KEYINPUT109), .B(n837), .ZN(G162) );
  XNOR2_X1 U936 ( .A(G27), .B(n838), .ZN(n849) );
  XNOR2_X1 U937 ( .A(KEYINPUT115), .B(G2067), .ZN(n839) );
  XNOR2_X1 U938 ( .A(n839), .B(G26), .ZN(n844) );
  XOR2_X1 U939 ( .A(G25), .B(G1991), .Z(n840) );
  NAND2_X1 U940 ( .A1(n840), .A2(G28), .ZN(n842) );
  XNOR2_X1 U941 ( .A(G33), .B(G2072), .ZN(n841) );
  NOR2_X1 U942 ( .A1(n842), .A2(n841), .ZN(n843) );
  NAND2_X1 U943 ( .A1(n844), .A2(n843), .ZN(n847) );
  XNOR2_X1 U944 ( .A(KEYINPUT116), .B(G1996), .ZN(n845) );
  XNOR2_X1 U945 ( .A(G32), .B(n845), .ZN(n846) );
  NOR2_X1 U946 ( .A1(n847), .A2(n846), .ZN(n848) );
  NAND2_X1 U947 ( .A1(n849), .A2(n848), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n850), .B(KEYINPUT53), .ZN(n853) );
  XOR2_X1 U949 ( .A(G2084), .B(KEYINPUT54), .Z(n851) );
  XNOR2_X1 U950 ( .A(G34), .B(n851), .ZN(n852) );
  NAND2_X1 U951 ( .A1(n853), .A2(n852), .ZN(n855) );
  XNOR2_X1 U952 ( .A(G35), .B(G2090), .ZN(n854) );
  NOR2_X1 U953 ( .A1(n855), .A2(n854), .ZN(n856) );
  XOR2_X1 U954 ( .A(KEYINPUT55), .B(n856), .Z(n857) );
  NOR2_X1 U955 ( .A1(G29), .A2(n857), .ZN(n948) );
  XNOR2_X1 U956 ( .A(KEYINPUT121), .B(G1341), .ZN(n858) );
  XNOR2_X1 U957 ( .A(n858), .B(G19), .ZN(n864) );
  XNOR2_X1 U958 ( .A(KEYINPUT59), .B(G4), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n859), .B(KEYINPUT123), .ZN(n860) );
  XNOR2_X1 U960 ( .A(G1348), .B(n860), .ZN(n862) );
  XNOR2_X1 U961 ( .A(G1956), .B(G20), .ZN(n861) );
  NOR2_X1 U962 ( .A1(n862), .A2(n861), .ZN(n863) );
  NAND2_X1 U963 ( .A1(n864), .A2(n863), .ZN(n867) );
  XNOR2_X1 U964 ( .A(KEYINPUT122), .B(G1981), .ZN(n865) );
  XNOR2_X1 U965 ( .A(G6), .B(n865), .ZN(n866) );
  NOR2_X1 U966 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U967 ( .A(KEYINPUT60), .B(n868), .ZN(n870) );
  XOR2_X1 U968 ( .A(G1961), .B(G5), .Z(n869) );
  NAND2_X1 U969 ( .A1(n870), .A2(n869), .ZN(n880) );
  XOR2_X1 U970 ( .A(G1966), .B(G21), .Z(n878) );
  XNOR2_X1 U971 ( .A(G1971), .B(G22), .ZN(n872) );
  XNOR2_X1 U972 ( .A(G1976), .B(G23), .ZN(n871) );
  NOR2_X1 U973 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U974 ( .A(KEYINPUT124), .B(n873), .Z(n875) );
  XNOR2_X1 U975 ( .A(G1986), .B(G24), .ZN(n874) );
  NOR2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U977 ( .A(n876), .B(KEYINPUT58), .ZN(n877) );
  NAND2_X1 U978 ( .A1(n878), .A2(n877), .ZN(n879) );
  NOR2_X1 U979 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U980 ( .A(KEYINPUT61), .B(n881), .Z(n882) );
  NOR2_X1 U981 ( .A1(G16), .A2(n882), .ZN(n883) );
  XOR2_X1 U982 ( .A(KEYINPUT125), .B(n883), .Z(n911) );
  XNOR2_X1 U983 ( .A(G1966), .B(G168), .ZN(n885) );
  NAND2_X1 U984 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U985 ( .A(n886), .B(KEYINPUT57), .ZN(n903) );
  XOR2_X1 U986 ( .A(G1348), .B(n1009), .Z(n887) );
  XNOR2_X1 U987 ( .A(n887), .B(KEYINPUT118), .ZN(n892) );
  XOR2_X1 U988 ( .A(n888), .B(G301), .Z(n889) );
  NOR2_X1 U989 ( .A1(n890), .A2(n889), .ZN(n891) );
  NAND2_X1 U990 ( .A1(n892), .A2(n891), .ZN(n901) );
  NAND2_X1 U991 ( .A1(G1971), .A2(G303), .ZN(n893) );
  NAND2_X1 U992 ( .A1(n894), .A2(n893), .ZN(n896) );
  XNOR2_X1 U993 ( .A(G1956), .B(G299), .ZN(n895) );
  NOR2_X1 U994 ( .A1(n896), .A2(n895), .ZN(n897) );
  NAND2_X1 U995 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U996 ( .A(KEYINPUT119), .B(n899), .Z(n900) );
  NOR2_X1 U997 ( .A1(n901), .A2(n900), .ZN(n902) );
  NAND2_X1 U998 ( .A1(n903), .A2(n902), .ZN(n905) );
  XOR2_X1 U999 ( .A(G1341), .B(n954), .Z(n904) );
  NOR2_X1 U1000 ( .A1(n905), .A2(n904), .ZN(n908) );
  XNOR2_X1 U1001 ( .A(G16), .B(KEYINPUT117), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(KEYINPUT56), .B(n906), .ZN(n907) );
  NOR2_X1 U1003 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(KEYINPUT120), .B(n909), .ZN(n910) );
  NOR2_X1 U1005 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1006 ( .A(KEYINPUT126), .B(n912), .ZN(n946) );
  NAND2_X1 U1007 ( .A1(G103), .A2(n995), .ZN(n914) );
  NAND2_X1 U1008 ( .A1(G139), .A2(n996), .ZN(n913) );
  NAND2_X1 U1009 ( .A1(n914), .A2(n913), .ZN(n921) );
  XNOR2_X1 U1010 ( .A(KEYINPUT112), .B(KEYINPUT47), .ZN(n919) );
  NAND2_X1 U1011 ( .A1(n991), .A2(G115), .ZN(n917) );
  NAND2_X1 U1012 ( .A1(n992), .A2(G127), .ZN(n915) );
  XOR2_X1 U1013 ( .A(KEYINPUT111), .B(n915), .Z(n916) );
  NAND2_X1 U1014 ( .A1(n917), .A2(n916), .ZN(n918) );
  XOR2_X1 U1015 ( .A(n919), .B(n918), .Z(n920) );
  NOR2_X1 U1016 ( .A1(n921), .A2(n920), .ZN(n1003) );
  XOR2_X1 U1017 ( .A(G2072), .B(n1003), .Z(n923) );
  XOR2_X1 U1018 ( .A(G164), .B(G2078), .Z(n922) );
  NOR2_X1 U1019 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1020 ( .A(KEYINPUT50), .B(n924), .ZN(n938) );
  XOR2_X1 U1021 ( .A(G2084), .B(G160), .Z(n925) );
  NOR2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n928) );
  NAND2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1024 ( .A1(n979), .A2(n929), .ZN(n930) );
  NAND2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n936) );
  XOR2_X1 U1026 ( .A(G2090), .B(G162), .Z(n932) );
  NOR2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1028 ( .A(KEYINPUT51), .B(n934), .ZN(n935) );
  NOR2_X1 U1029 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1030 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1031 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1032 ( .A(KEYINPUT52), .B(n941), .Z(n942) );
  NOR2_X1 U1033 ( .A1(KEYINPUT55), .A2(n942), .ZN(n943) );
  XOR2_X1 U1034 ( .A(KEYINPUT114), .B(n943), .Z(n944) );
  NAND2_X1 U1035 ( .A1(n944), .A2(G29), .ZN(n945) );
  NAND2_X1 U1036 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1037 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1038 ( .A1(n949), .A2(G11), .ZN(n950) );
  XOR2_X1 U1039 ( .A(KEYINPUT62), .B(n950), .Z(G311) );
  XNOR2_X1 U1040 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1041 ( .A(G120), .ZN(G236) );
  INV_X1 U1042 ( .A(G96), .ZN(G221) );
  INV_X1 U1043 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1044 ( .A1(n952), .A2(n951), .ZN(G325) );
  INV_X1 U1045 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1046 ( .A(n954), .B(n953), .Z(n955) );
  NOR2_X1 U1047 ( .A1(n955), .A2(G860), .ZN(n957) );
  XOR2_X1 U1048 ( .A(n957), .B(n956), .Z(G145) );
  XOR2_X1 U1049 ( .A(G2100), .B(G2096), .Z(n959) );
  XNOR2_X1 U1050 ( .A(G2090), .B(KEYINPUT43), .ZN(n958) );
  XNOR2_X1 U1051 ( .A(n959), .B(n958), .ZN(n960) );
  XOR2_X1 U1052 ( .A(n960), .B(G2678), .Z(n962) );
  XNOR2_X1 U1053 ( .A(G2072), .B(KEYINPUT106), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(n962), .B(n961), .ZN(n966) );
  XOR2_X1 U1055 ( .A(KEYINPUT42), .B(G2078), .Z(n964) );
  XNOR2_X1 U1056 ( .A(G2084), .B(G2067), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(n964), .B(n963), .ZN(n965) );
  XNOR2_X1 U1058 ( .A(n966), .B(n965), .ZN(G227) );
  XOR2_X1 U1059 ( .A(G1981), .B(G1971), .Z(n968) );
  XNOR2_X1 U1060 ( .A(G1966), .B(G1956), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(n968), .B(n967), .ZN(n973) );
  XOR2_X1 U1062 ( .A(KEYINPUT107), .B(G2474), .Z(n971) );
  XOR2_X1 U1063 ( .A(n969), .B(G1961), .Z(n970) );
  XNOR2_X1 U1064 ( .A(n971), .B(n970), .ZN(n972) );
  XOR2_X1 U1065 ( .A(n973), .B(n972), .Z(n976) );
  XOR2_X1 U1066 ( .A(G1976), .B(n974), .Z(n975) );
  XNOR2_X1 U1067 ( .A(n976), .B(n975), .ZN(n978) );
  XOR2_X1 U1068 ( .A(G1986), .B(KEYINPUT41), .Z(n977) );
  XNOR2_X1 U1069 ( .A(n978), .B(n977), .ZN(G229) );
  XOR2_X1 U1070 ( .A(KEYINPUT110), .B(KEYINPUT48), .Z(n981) );
  XNOR2_X1 U1071 ( .A(n979), .B(KEYINPUT46), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(n981), .B(n980), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(n983), .B(n982), .ZN(n987) );
  XOR2_X1 U1074 ( .A(n985), .B(n984), .Z(n986) );
  XNOR2_X1 U1075 ( .A(n987), .B(n986), .ZN(n988) );
  XOR2_X1 U1076 ( .A(n988), .B(G162), .Z(n990) );
  XNOR2_X1 U1077 ( .A(G160), .B(G164), .ZN(n989) );
  XNOR2_X1 U1078 ( .A(n990), .B(n989), .ZN(n1005) );
  NAND2_X1 U1079 ( .A1(G118), .A2(n991), .ZN(n994) );
  NAND2_X1 U1080 ( .A1(G130), .A2(n992), .ZN(n993) );
  NAND2_X1 U1081 ( .A1(n994), .A2(n993), .ZN(n1001) );
  NAND2_X1 U1082 ( .A1(G106), .A2(n995), .ZN(n998) );
  NAND2_X1 U1083 ( .A1(G142), .A2(n996), .ZN(n997) );
  NAND2_X1 U1084 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1085 ( .A(KEYINPUT45), .B(n999), .Z(n1000) );
  NOR2_X1 U1086 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1087 ( .A(n1003), .B(n1002), .ZN(n1004) );
  XNOR2_X1 U1088 ( .A(n1005), .B(n1004), .ZN(n1006) );
  NOR2_X1 U1089 ( .A1(G37), .A2(n1006), .ZN(G395) );
  XOR2_X1 U1090 ( .A(G286), .B(G171), .Z(n1008) );
  XNOR2_X1 U1091 ( .A(n1008), .B(n1007), .ZN(n1010) );
  XOR2_X1 U1092 ( .A(n1010), .B(n1009), .Z(n1011) );
  NOR2_X1 U1093 ( .A1(G37), .A2(n1011), .ZN(G397) );
  NAND2_X1 U1094 ( .A1(G319), .A2(n1012), .ZN(n1016) );
  NOR2_X1 U1095 ( .A1(G227), .A2(G229), .ZN(n1013) );
  XOR2_X1 U1096 ( .A(KEYINPUT49), .B(n1013), .Z(n1014) );
  XNOR2_X1 U1097 ( .A(n1014), .B(KEYINPUT113), .ZN(n1015) );
  NOR2_X1 U1098 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  NOR2_X1 U1099 ( .A1(G395), .A2(G397), .ZN(n1017) );
  NAND2_X1 U1100 ( .A1(n1018), .A2(n1017), .ZN(G225) );
  INV_X1 U1101 ( .A(G225), .ZN(G308) );
  INV_X1 U1102 ( .A(G108), .ZN(G238) );
endmodule

