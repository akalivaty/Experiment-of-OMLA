//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 1 0 0 0 0 1 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1300, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT65), .ZN(G353));
  OAI21_X1  g0010(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0011(.A(G1), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G13), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT0), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n220), .B1(new_n203), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  INV_X1    g0025(.A(G77), .ZN(new_n226));
  INV_X1    g0026(.A(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G107), .ZN(new_n228));
  INV_X1    g0028(.A(G264), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n225), .B1(new_n226), .B2(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  OAI22_X1  g0030(.A1(new_n224), .A2(new_n230), .B1(new_n212), .B2(new_n213), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n232), .A2(new_n213), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT66), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n206), .A2(new_n207), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  OAI221_X1 g0036(.A(new_n219), .B1(KEYINPUT1), .B2(new_n231), .C1(new_n234), .C2(new_n236), .ZN(new_n237));
  AOI21_X1  g0037(.A(new_n237), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  INV_X1    g0039(.A(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT2), .B(G226), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G358));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XOR2_X1   g0048(.A(G107), .B(G116), .Z(new_n249));
  XOR2_X1   g0049(.A(new_n248), .B(new_n249), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT67), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n207), .A2(G68), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n203), .A2(G50), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G58), .B(G77), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n251), .B(new_n256), .ZN(G351));
  AND2_X1   g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  OAI211_X1 g0059(.A(G250), .B(G1698), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G283), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  AOI21_X1  g0066(.A(G1698), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT84), .ZN(new_n268));
  AND2_X1   g0068(.A1(KEYINPUT4), .A2(G244), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n271), .B(new_n269), .C1(new_n258), .C2(new_n259), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT84), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n262), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n264), .A2(KEYINPUT77), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT77), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G33), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n263), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  OAI211_X1 g0078(.A(G244), .B(new_n271), .C1(new_n278), .C2(new_n259), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT4), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n274), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n232), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G33), .A2(G41), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT85), .ZN(new_n288));
  INV_X1    g0088(.A(G274), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n289), .B1(new_n283), .B2(new_n284), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT5), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n212), .B(G45), .C1(new_n291), .C2(G41), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT68), .B(G41), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n290), .B(new_n293), .C1(KEYINPUT5), .C2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G41), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT68), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT68), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G41), .ZN(new_n299));
  AOI21_X1  g0099(.A(KEYINPUT5), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n285), .B1(new_n300), .B2(new_n292), .ZN(new_n301));
  INV_X1    g0101(.A(G257), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n295), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n287), .A2(new_n288), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n285), .B1(new_n274), .B2(new_n281), .ZN(new_n306));
  OAI21_X1  g0106(.A(KEYINPUT85), .B1(new_n306), .B2(new_n303), .ZN(new_n307));
  AND3_X1   g0107(.A1(new_n305), .A2(G190), .A3(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n212), .A2(G13), .A3(G20), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n309), .A2(G97), .ZN(new_n310));
  NAND3_X1  g0110(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n232), .ZN(new_n312));
  INV_X1    g0112(.A(new_n309), .ZN(new_n313));
  AOI211_X1 g0113(.A(new_n312), .B(new_n313), .C1(new_n212), .C2(G33), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n310), .B1(new_n314), .B2(G97), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(G20), .A2(G33), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G77), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT6), .ZN(new_n319));
  AND2_X1   g0119(.A1(G97), .A2(G107), .ZN(new_n320));
  NOR2_X1   g0120(.A1(G97), .A2(G107), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(KEYINPUT6), .A2(G97), .ZN(new_n323));
  OAI21_X1  g0123(.A(KEYINPUT83), .B1(new_n323), .B2(G107), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT83), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n325), .A2(new_n228), .A3(KEYINPUT6), .A4(G97), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n322), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G20), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n258), .A2(new_n259), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT7), .B1(new_n329), .B2(new_n213), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT7), .ZN(new_n331));
  NOR3_X1   g0131(.A1(new_n258), .A2(new_n331), .A3(G20), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n275), .A2(new_n277), .A3(new_n263), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT79), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT79), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n332), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n330), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n318), .B(new_n328), .C1(new_n338), .C2(new_n228), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n316), .B1(new_n339), .B2(new_n312), .ZN(new_n340));
  OAI21_X1  g0140(.A(G200), .B1(new_n306), .B2(new_n303), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(G169), .B1(new_n305), .B2(new_n307), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n303), .B1(new_n282), .B2(new_n286), .ZN(new_n344));
  INV_X1    g0144(.A(G179), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n328), .A2(new_n318), .ZN(new_n347));
  INV_X1    g0147(.A(new_n330), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n332), .A2(new_n333), .A3(new_n336), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n336), .B1(new_n332), .B2(new_n333), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n347), .B1(new_n351), .B2(G107), .ZN(new_n352));
  INV_X1    g0152(.A(new_n312), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n315), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n346), .A2(new_n354), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n308), .A2(new_n342), .B1(new_n343), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g0156(.A(KEYINPUT15), .B(G87), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(new_n309), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT77), .B(G33), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n265), .B1(new_n360), .B2(new_n263), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n361), .A2(new_n213), .A3(G68), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n264), .A2(G20), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT19), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n363), .A2(new_n364), .A3(G97), .ZN(new_n365));
  NAND2_X1  g0165(.A1(G33), .A2(G97), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n321), .A2(new_n222), .B1(new_n366), .B2(new_n213), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n365), .B1(new_n367), .B2(new_n364), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n362), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n359), .B1(new_n369), .B2(new_n312), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n314), .A2(new_n358), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n361), .A2(G238), .A3(new_n271), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n275), .A2(new_n277), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G116), .ZN(new_n375));
  OAI211_X1 g0175(.A(G244), .B(G1698), .C1(new_n278), .C2(new_n259), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n373), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n286), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n212), .A2(new_n289), .A3(G45), .ZN(new_n379));
  INV_X1    g0179(.A(G45), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n223), .B1(new_n380), .B2(G1), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n285), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n378), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n372), .B1(new_n384), .B2(G179), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n382), .B1(new_n377), .B2(new_n286), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n386), .A2(G169), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n314), .A2(G87), .ZN(new_n388));
  INV_X1    g0188(.A(G200), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n370), .B(new_n388), .C1(new_n386), .C2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(G190), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n384), .A2(new_n391), .ZN(new_n392));
  OAI22_X1  g0192(.A1(new_n385), .A2(new_n387), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n356), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n297), .A2(new_n299), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n212), .B(G274), .C1(new_n395), .C2(G45), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n212), .B1(G41), .B2(G45), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n285), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n396), .B1(new_n221), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT72), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n285), .A2(new_n397), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G238), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n403), .A2(KEYINPUT72), .A3(new_n396), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n267), .A2(G226), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n265), .A2(new_n266), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(G1698), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n405), .B(new_n366), .C1(new_n240), .C2(new_n407), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n401), .A2(new_n404), .B1(new_n286), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT13), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT73), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n286), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n399), .A2(new_n400), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT72), .B1(new_n403), .B2(new_n396), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT73), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n415), .A2(new_n416), .A3(KEYINPUT13), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n411), .A2(new_n417), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n410), .B(new_n412), .C1(new_n413), .C2(new_n414), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT74), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n409), .A2(KEYINPUT74), .A3(new_n410), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n418), .A2(G179), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n419), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n401), .A2(new_n404), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n410), .B1(new_n425), .B2(new_n412), .ZN(new_n426));
  OAI21_X1  g0226(.A(G169), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT14), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT14), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(G169), .C1(new_n424), .C2(new_n426), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n423), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n313), .A2(new_n203), .ZN(new_n432));
  XNOR2_X1  g0232(.A(new_n432), .B(KEYINPUT12), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n363), .A2(G77), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n317), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n353), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT11), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT70), .B1(new_n313), .B2(new_n312), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT70), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n309), .A2(new_n440), .A3(new_n232), .A4(new_n311), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n212), .A2(G20), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(G68), .A3(new_n443), .ZN(new_n444));
  OR2_X1    g0244(.A1(new_n436), .A2(KEYINPUT11), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n438), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT75), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT75), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n438), .A2(new_n444), .A3(new_n448), .A4(new_n445), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n431), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(G200), .B1(new_n424), .B2(new_n426), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n418), .A2(new_n421), .A3(new_n422), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n453), .B(new_n450), .C1(new_n454), .C2(new_n391), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n452), .A2(KEYINPUT76), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(KEYINPUT76), .B1(new_n452), .B2(new_n455), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n402), .A2(G226), .ZN(new_n458));
  INV_X1    g0258(.A(G223), .ZN(new_n459));
  OAI22_X1  g0259(.A1(new_n407), .A2(new_n459), .B1(new_n226), .B2(new_n406), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n460), .B1(G222), .B2(new_n267), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n396), .B(new_n458), .C1(new_n461), .C2(new_n285), .ZN(new_n462));
  INV_X1    g0262(.A(G169), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n208), .A2(G20), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n317), .A2(G150), .ZN(new_n466));
  XNOR2_X1  g0266(.A(KEYINPUT8), .B(G58), .ZN(new_n467));
  XNOR2_X1  g0267(.A(new_n467), .B(KEYINPUT69), .ZN(new_n468));
  INV_X1    g0268(.A(new_n363), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n465), .B(new_n466), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n312), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n309), .A2(G50), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n353), .A2(new_n443), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n472), .B1(new_n474), .B2(G50), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n464), .B(new_n476), .C1(G179), .C2(new_n462), .ZN(new_n477));
  INV_X1    g0277(.A(new_n467), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n478), .A2(new_n317), .B1(G20), .B2(G77), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n479), .B1(new_n469), .B2(new_n357), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n480), .A2(new_n312), .B1(new_n226), .B2(new_n313), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n442), .A2(G77), .A3(new_n443), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n396), .B1(new_n227), .B2(new_n398), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n267), .A2(G232), .ZN(new_n485));
  OAI221_X1 g0285(.A(new_n485), .B1(new_n228), .B2(new_n406), .C1(new_n221), .C2(new_n407), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n484), .B1(new_n486), .B2(new_n286), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n483), .B1(G190), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n389), .B2(new_n487), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n345), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n483), .B(new_n490), .C1(G169), .C2(new_n487), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n471), .A2(KEYINPUT71), .A3(new_n475), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(KEYINPUT71), .B1(new_n471), .B2(new_n475), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT9), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT71), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n476), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT9), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(new_n499), .A3(new_n493), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT10), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n462), .A2(new_n391), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(G200), .B2(new_n462), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n501), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n502), .B1(new_n501), .B2(new_n504), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n477), .B(new_n492), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n456), .A2(new_n457), .A3(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n204), .B(new_n205), .C1(new_n202), .C2(new_n203), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n509), .A2(G20), .B1(G159), .B2(new_n317), .ZN(new_n510));
  NOR3_X1   g0310(.A1(new_n361), .A2(new_n331), .A3(G20), .ZN(new_n511));
  OAI21_X1  g0311(.A(KEYINPUT78), .B1(new_n278), .B2(new_n259), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT78), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n513), .B(new_n265), .C1(new_n360), .C2(new_n263), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n213), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n511), .B1(new_n516), .B2(new_n331), .ZN(new_n517));
  OAI211_X1 g0317(.A(KEYINPUT16), .B(new_n510), .C1(new_n517), .C2(new_n203), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n510), .B1(new_n338), .B2(new_n203), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT16), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n518), .A2(new_n312), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G33), .A2(G87), .ZN(new_n523));
  XNOR2_X1  g0323(.A(new_n523), .B(KEYINPUT80), .ZN(new_n524));
  AND2_X1   g0324(.A1(G226), .A2(G1698), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n524), .B1(new_n361), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n361), .A2(G223), .A3(new_n271), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n286), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT81), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n285), .A2(G232), .A3(new_n397), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n396), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n530), .B1(new_n396), .B2(new_n531), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n529), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n389), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(G190), .B2(new_n535), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n468), .A2(new_n474), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(new_n309), .B2(new_n468), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n522), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  XOR2_X1   g0341(.A(KEYINPUT82), .B(KEYINPUT17), .Z(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n510), .ZN(new_n544));
  OR3_X1    g0344(.A1(new_n361), .A2(new_n331), .A3(G20), .ZN(new_n545));
  AOI21_X1  g0345(.A(G20), .B1(new_n512), .B2(new_n514), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n546), .B2(KEYINPUT7), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n544), .B1(new_n547), .B2(G68), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n353), .B1(new_n548), .B2(KEYINPUT16), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n539), .B1(new_n549), .B2(new_n521), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT17), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n551), .A2(KEYINPUT82), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n550), .A2(new_n537), .A3(new_n553), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n543), .A2(new_n554), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n529), .A2(new_n534), .A3(G179), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n463), .B1(new_n529), .B2(new_n534), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(KEYINPUT18), .B1(new_n550), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n522), .A2(new_n540), .ZN(new_n560));
  INV_X1    g0360(.A(new_n557), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n529), .A2(new_n534), .A3(G179), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT18), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n560), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n559), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n555), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n508), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(G116), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n311), .A2(new_n232), .B1(G20), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(G20), .B1(G33), .B2(G283), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n264), .A2(G97), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n572), .A2(new_n573), .A3(KEYINPUT87), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT87), .B1(new_n572), .B2(new_n573), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n571), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT20), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(KEYINPUT20), .B(new_n571), .C1(new_n574), .C2(new_n575), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n570), .B1(new_n212), .B2(G33), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n439), .A2(new_n441), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n313), .A2(new_n570), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n302), .A2(new_n271), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n229), .A2(G1698), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n586), .B(new_n587), .C1(new_n278), .C2(new_n259), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n329), .A2(G303), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n286), .ZN(new_n591));
  OAI211_X1 g0391(.A(G270), .B(new_n285), .C1(new_n300), .C2(new_n292), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n592), .A2(new_n295), .A3(KEYINPUT86), .ZN(new_n593));
  AOI21_X1  g0393(.A(KEYINPUT86), .B1(new_n592), .B2(new_n295), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n591), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n585), .B1(new_n595), .B2(G200), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n391), .B2(new_n595), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n285), .B1(new_n588), .B2(new_n589), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n592), .A2(new_n295), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT86), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n592), .A2(new_n295), .A3(KEYINPUT86), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n598), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n603), .A2(G179), .A3(new_n585), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT21), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n463), .B1(new_n580), .B2(new_n584), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n605), .B1(new_n606), .B2(new_n595), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n606), .A2(new_n605), .A3(new_n595), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n597), .B(new_n604), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n314), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT25), .B1(new_n313), .B2(new_n228), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n313), .A2(KEYINPUT25), .A3(new_n228), .ZN(new_n613));
  OAI22_X1  g0413(.A1(new_n611), .A2(new_n228), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT88), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT22), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n213), .A2(G87), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n616), .B1(new_n329), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n228), .A2(G20), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT23), .ZN(new_n620));
  XNOR2_X1  g0420(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n374), .A2(new_n213), .A3(G116), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n618), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n616), .A2(new_n222), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n213), .B(new_n624), .C1(new_n278), .C2(new_n259), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n615), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT24), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n353), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n623), .A2(new_n615), .A3(new_n625), .ZN(new_n629));
  INV_X1    g0429(.A(new_n625), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n618), .A2(new_n621), .A3(new_n622), .ZN(new_n631));
  OAI21_X1  g0431(.A(KEYINPUT88), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n629), .A2(new_n632), .A3(KEYINPUT24), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n614), .B1(new_n628), .B2(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(G264), .B(new_n285), .C1(new_n300), .C2(new_n292), .ZN(new_n635));
  NOR2_X1   g0435(.A1(G250), .A2(G1698), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n636), .B1(new_n302), .B2(G1698), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n361), .A2(new_n637), .B1(G294), .B2(new_n374), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n295), .B(new_n635), .C1(new_n638), .C2(new_n285), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n463), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(G179), .B2(new_n639), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n634), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n628), .A2(new_n633), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n639), .A2(new_n389), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n644), .B1(G190), .B2(new_n639), .ZN(new_n645));
  INV_X1    g0445(.A(new_n614), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n643), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT89), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT89), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n634), .A2(new_n649), .A3(new_n645), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n642), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  AND4_X1   g0451(.A1(new_n394), .A2(new_n569), .A3(new_n610), .A4(new_n651), .ZN(G372));
  OAI21_X1  g0452(.A(new_n604), .B1(new_n608), .B2(new_n607), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT90), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n604), .B(KEYINPUT90), .C1(new_n608), .C2(new_n607), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n642), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n648), .A2(new_n650), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(new_n394), .A3(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n385), .A2(new_n387), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n305), .A2(new_n307), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n463), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n346), .A2(new_n354), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n663), .B1(new_n667), .B2(new_n393), .ZN(new_n668));
  INV_X1    g0468(.A(new_n390), .ZN(new_n669));
  INV_X1    g0469(.A(new_n392), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n386), .A2(new_n345), .B1(new_n370), .B2(new_n371), .ZN(new_n671));
  INV_X1    g0471(.A(new_n387), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n669), .A2(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n343), .A2(new_n355), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(new_n674), .A3(KEYINPUT26), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n662), .B1(new_n668), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n661), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n569), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n477), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n564), .B1(new_n560), .B2(new_n563), .ZN(new_n680));
  AOI211_X1 g0480(.A(KEYINPUT18), .B(new_n558), .C1(new_n522), .C2(new_n540), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n491), .ZN(new_n683));
  AOI22_X1  g0483(.A1(new_n455), .A2(new_n683), .B1(new_n431), .B2(new_n451), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n682), .B1(new_n684), .B2(new_n555), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n505), .A2(new_n506), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n679), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n678), .A2(new_n687), .ZN(G369));
  NOR3_X1   g0488(.A1(new_n215), .A2(G1), .A3(G20), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n690), .A2(KEYINPUT91), .A3(KEYINPUT27), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(KEYINPUT91), .B1(new_n690), .B2(KEYINPUT27), .ZN(new_n693));
  OAI221_X1 g0493(.A(G213), .B1(KEYINPUT27), .B2(new_n690), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(G343), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n585), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n657), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n609), .B1(new_n698), .B2(new_n697), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT92), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n642), .A2(new_n697), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n634), .A2(new_n697), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n660), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n705), .B1(new_n707), .B2(new_n658), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT92), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n700), .A2(new_n709), .A3(new_n701), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n703), .A2(new_n708), .A3(G330), .A4(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n707), .A2(new_n658), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n653), .A2(new_n697), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n705), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n711), .A2(new_n715), .ZN(G399));
  NOR2_X1   g0516(.A1(new_n216), .A2(new_n395), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n235), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n321), .A2(new_n222), .A3(new_n570), .ZN(new_n719));
  OR3_X1    g0519(.A1(new_n717), .A2(new_n212), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n718), .B1(new_n720), .B2(KEYINPUT93), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n721), .B1(KEYINPUT93), .B2(new_n720), .ZN(new_n722));
  XOR2_X1   g0522(.A(new_n722), .B(KEYINPUT28), .Z(new_n723));
  NAND4_X1  g0523(.A1(new_n394), .A2(new_n651), .A3(new_n610), .A4(new_n697), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT30), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n601), .A2(new_n602), .ZN(new_n726));
  INV_X1    g0526(.A(new_n635), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n361), .A2(new_n637), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n374), .A2(G294), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n727), .B1(new_n730), .B2(new_n286), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n598), .A2(new_n345), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n386), .A2(new_n726), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n725), .B1(new_n664), .B2(new_n733), .ZN(new_n734));
  AND4_X1   g0534(.A1(new_n386), .A2(new_n726), .A3(new_n731), .A4(new_n732), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n735), .A2(KEYINPUT30), .A3(new_n307), .A4(new_n305), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n603), .A2(new_n386), .A3(G179), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n639), .B1(new_n306), .B2(new_n303), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT94), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI211_X1 g0540(.A(KEYINPUT94), .B(new_n639), .C1(new_n306), .C2(new_n303), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n737), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n734), .A2(new_n736), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(KEYINPUT31), .B1(new_n743), .B2(new_n696), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n724), .B1(KEYINPUT95), .B2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT95), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n743), .A2(new_n696), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT31), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n743), .A2(KEYINPUT31), .A3(new_n696), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n746), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n745), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G330), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n356), .A2(KEYINPUT96), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n393), .B1(new_n648), .B2(new_n650), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n653), .A2(new_n642), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT96), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n757), .B1(new_n343), .B2(new_n355), .C1(new_n308), .C2(new_n342), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n754), .A2(new_n755), .A3(new_n756), .A4(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n696), .B1(new_n759), .B2(new_n676), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(KEYINPUT29), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n696), .B1(new_n661), .B2(new_n676), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n761), .B1(new_n762), .B2(KEYINPUT29), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n753), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n723), .B1(new_n764), .B2(G1), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT97), .Z(G364));
  NAND3_X1  g0566(.A1(new_n703), .A2(G330), .A3(new_n710), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n215), .A2(G20), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n212), .B1(new_n768), .B2(G45), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n717), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n767), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n703), .A2(new_n710), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G330), .ZN(new_n777));
  OR3_X1    g0577(.A1(KEYINPUT98), .A2(G13), .A3(G33), .ZN(new_n778));
  OAI21_X1  g0578(.A(KEYINPUT98), .B1(G13), .B2(G33), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(G20), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n775), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n216), .A2(new_n329), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n784), .A2(G355), .B1(new_n570), .B2(new_n216), .ZN(new_n785));
  INV_X1    g0585(.A(new_n515), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n216), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n235), .A2(new_n380), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(new_n256), .B2(new_n380), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n785), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n232), .B1(G20), .B2(new_n463), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n782), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n772), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n213), .A2(G179), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n795), .A2(G190), .A3(G200), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n795), .A2(new_n391), .A3(G200), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n222), .A2(new_n796), .B1(new_n797), .B2(new_n228), .ZN(new_n798));
  NOR3_X1   g0598(.A1(new_n391), .A2(G179), .A3(G200), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n213), .ZN(new_n800));
  INV_X1    g0600(.A(G97), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(G20), .A2(G179), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n803), .A2(G190), .A3(G200), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n803), .A2(new_n391), .A3(G200), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n406), .B1(new_n805), .B2(new_n226), .C1(new_n202), .C2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n803), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n809), .A2(new_n391), .A3(G200), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n802), .B(new_n808), .C1(G68), .C2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(G190), .A2(G200), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n795), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(G159), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT32), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n809), .A2(G190), .A3(G200), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n798), .B(new_n818), .C1(G50), .C2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n822), .A2(KEYINPUT99), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n822), .A2(KEYINPUT99), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n796), .B(KEYINPUT100), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(G303), .ZN(new_n826));
  INV_X1    g0626(.A(G311), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n805), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(G322), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n329), .B1(new_n807), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n814), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n828), .B(new_n830), .C1(G329), .C2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n797), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G283), .A2(new_n833), .B1(new_n820), .B2(G326), .ZN(new_n834));
  INV_X1    g0634(.A(new_n800), .ZN(new_n835));
  XNOR2_X1  g0635(.A(KEYINPUT33), .B(G317), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n835), .A2(G294), .B1(new_n811), .B2(new_n836), .ZN(new_n837));
  AND4_X1   g0637(.A1(new_n826), .A2(new_n832), .A3(new_n834), .A4(new_n837), .ZN(new_n838));
  NOR3_X1   g0638(.A1(new_n823), .A2(new_n824), .A3(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n792), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n794), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n774), .A2(new_n777), .B1(new_n783), .B2(new_n841), .ZN(G396));
  AOI22_X1  g0642(.A1(new_n811), .A2(G283), .B1(G116), .B2(new_n804), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT101), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n797), .A2(new_n222), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n845), .B(new_n802), .C1(G303), .C2(new_n820), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n825), .A2(G107), .ZN(new_n847));
  INV_X1    g0647(.A(G294), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n329), .B1(new_n807), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G311), .B2(new_n831), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n844), .A2(new_n846), .A3(new_n847), .A4(new_n850), .ZN(new_n851));
  AOI22_X1  g0651(.A1(G143), .A2(new_n806), .B1(new_n804), .B2(G159), .ZN(new_n852));
  INV_X1    g0652(.A(G137), .ZN(new_n853));
  INV_X1    g0653(.A(G150), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n852), .B1(new_n853), .B2(new_n819), .C1(new_n854), .C2(new_n810), .ZN(new_n855));
  XOR2_X1   g0655(.A(new_n855), .B(KEYINPUT34), .Z(new_n856));
  INV_X1    g0656(.A(G132), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n797), .A2(new_n203), .B1(new_n814), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(G58), .B2(new_n835), .ZN(new_n859));
  INV_X1    g0659(.A(new_n825), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n786), .B(new_n859), .C1(new_n860), .C2(new_n207), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n851), .B1(new_n856), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n792), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n780), .A2(new_n792), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n772), .B1(new_n226), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n483), .A2(new_n696), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n489), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n491), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n683), .A2(new_n697), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n863), .B(new_n865), .C1(new_n871), .C2(new_n781), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT102), .ZN(new_n873));
  OR2_X1    g0673(.A1(new_n762), .A2(new_n871), .ZN(new_n874));
  INV_X1    g0674(.A(new_n341), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n875), .A2(new_n354), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n305), .A2(G190), .A3(new_n307), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n665), .A2(new_n666), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n660), .A2(new_n878), .A3(new_n673), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n642), .B1(new_n655), .B2(new_n656), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n662), .ZN(new_n882));
  NOR3_X1   g0682(.A1(new_n667), .A2(new_n393), .A3(new_n663), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT26), .B1(new_n673), .B2(new_n674), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n697), .B(new_n871), .C1(new_n881), .C2(new_n885), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n874), .A2(G330), .A3(new_n752), .A4(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n873), .B1(new_n887), .B2(new_n772), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n874), .A2(new_n886), .B1(new_n752), .B2(G330), .ZN(new_n889));
  OR2_X1    g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n887), .A2(new_n873), .A3(new_n772), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n872), .B1(new_n890), .B2(new_n891), .ZN(G384));
  NOR2_X1   g0692(.A1(new_n768), .A2(new_n212), .ZN(new_n893));
  INV_X1    g0693(.A(G330), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n510), .B1(new_n517), .B2(new_n203), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n520), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n539), .B1(new_n897), .B2(new_n549), .ZN(new_n898));
  INV_X1    g0698(.A(new_n694), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n563), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n541), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(KEYINPUT103), .A3(KEYINPUT37), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n560), .A2(new_n563), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n560), .A2(new_n899), .ZN(new_n904));
  XOR2_X1   g0704(.A(KEYINPUT104), .B(KEYINPUT37), .Z(new_n905));
  NAND4_X1  g0705(.A1(new_n903), .A2(new_n904), .A3(new_n541), .A4(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT103), .B1(new_n901), .B2(KEYINPUT37), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n898), .A2(new_n694), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n543), .A2(new_n554), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n911), .B1(new_n682), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n895), .B1(new_n909), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT103), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n518), .A2(new_n312), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n548), .A2(KEYINPUT16), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n540), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n558), .A2(new_n694), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n918), .A2(new_n919), .B1(new_n550), .B2(new_n537), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT37), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n915), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(new_n906), .A3(new_n902), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n910), .B1(new_n555), .B2(new_n566), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n923), .A2(KEYINPUT38), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n914), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n451), .A2(new_n696), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n452), .A2(new_n455), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n453), .A2(new_n450), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n421), .A2(new_n422), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n411), .B2(new_n417), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n929), .B1(new_n931), .B2(G190), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n451), .B(new_n696), .C1(new_n932), .C2(new_n431), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n870), .B1(new_n928), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n724), .A2(new_n749), .A3(new_n750), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT40), .B1(new_n926), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n550), .A2(new_n694), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n555), .B2(new_n566), .ZN(new_n939));
  INV_X1    g0739(.A(new_n905), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n541), .B1(new_n550), .B2(new_n558), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n940), .B1(new_n941), .B2(new_n938), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n906), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n895), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n925), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n934), .A2(KEYINPUT40), .A3(new_n935), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n937), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n569), .A2(new_n935), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n894), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n949), .B2(new_n950), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT39), .ZN(new_n953));
  AND3_X1   g0753(.A1(new_n923), .A2(KEYINPUT38), .A3(new_n924), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT38), .B1(new_n939), .B2(new_n943), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n914), .A2(KEYINPUT39), .A3(new_n925), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n452), .A2(new_n696), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n928), .A2(new_n933), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(new_n886), .B2(new_n869), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n926), .A2(new_n962), .B1(new_n566), .B2(new_n694), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n687), .B1(new_n763), .B2(new_n568), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n964), .B(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n893), .B1(new_n952), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n966), .B2(new_n952), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n327), .A2(KEYINPUT35), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n327), .A2(KEYINPUT35), .ZN(new_n970));
  NOR4_X1   g0770(.A1(new_n969), .A2(new_n970), .A3(new_n570), .A4(new_n234), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(KEYINPUT36), .Z(new_n972));
  OAI211_X1 g0772(.A(new_n235), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n252), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n974), .A2(G1), .A3(new_n215), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n968), .A2(new_n972), .A3(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT105), .ZN(G367));
  NAND2_X1  g0777(.A1(new_n370), .A2(new_n388), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n696), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n662), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n980), .B1(new_n393), .B2(new_n979), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT106), .ZN(new_n982));
  XOR2_X1   g0782(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n754), .B(new_n758), .C1(new_n340), .C2(new_n697), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n674), .A2(new_n696), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n660), .A2(new_n706), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n988), .A2(new_n653), .A3(new_n658), .A4(new_n697), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT42), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n667), .B1(new_n985), .B2(new_n658), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n697), .ZN(new_n994));
  OAI21_X1  g0794(.A(KEYINPUT42), .B1(new_n987), .B2(new_n989), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n992), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT109), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n992), .A2(KEYINPUT109), .A3(new_n994), .A4(new_n995), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n982), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(KEYINPUT43), .ZN(new_n1002));
  OR3_X1    g0802(.A1(new_n711), .A2(KEYINPUT108), .A3(new_n987), .ZN(new_n1003));
  OAI21_X1  g0803(.A(KEYINPUT108), .B1(new_n711), .B2(new_n987), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  AND3_X1   g0806(.A1(new_n1000), .A2(new_n1002), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1006), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n984), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n1005), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n984), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1000), .A2(new_n1006), .A3(new_n1002), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n717), .B(KEYINPUT41), .Z(new_n1015));
  INV_X1    g0815(.A(KEYINPUT45), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n989), .A2(new_n704), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1016), .B1(new_n1017), .B2(new_n987), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n985), .A2(new_n986), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n715), .A2(KEYINPUT45), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1017), .A2(KEYINPUT44), .A3(new_n987), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT44), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n715), .B2(new_n1019), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1021), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n711), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1026), .A2(KEYINPUT110), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(KEYINPUT110), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1029), .A2(new_n1021), .A3(new_n1025), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n712), .A2(new_n704), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n713), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n989), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(new_n767), .Z(new_n1034));
  NAND4_X1  g0834(.A1(new_n1028), .A2(new_n764), .A3(new_n1030), .A4(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1015), .B1(new_n1035), .B2(new_n764), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1009), .B(new_n1014), .C1(new_n770), .C2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n793), .B1(new_n217), .B2(new_n357), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n246), .B2(new_n787), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n807), .A2(new_n854), .B1(new_n814), .B2(new_n853), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n329), .B(new_n1040), .C1(G50), .C2(new_n804), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n835), .A2(G68), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n796), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G58), .A2(new_n1043), .B1(new_n811), .B2(G159), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(G77), .A2(new_n833), .B1(new_n820), .B2(G143), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n833), .A2(G97), .ZN(new_n1047));
  INV_X1    g0847(.A(G317), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1047), .B1(new_n1048), .B2(new_n814), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n786), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT111), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT46), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n825), .B2(G116), .ZN(new_n1054));
  NOR3_X1   g0854(.A1(new_n796), .A2(KEYINPUT46), .A3(new_n570), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1052), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(G303), .ZN(new_n1057));
  INV_X1    g0857(.A(G283), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n807), .A2(new_n1057), .B1(new_n805), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G107), .B2(new_n835), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G294), .A2(new_n811), .B1(new_n820), .B2(G311), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1046), .B1(new_n1056), .B2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT47), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n772), .B(new_n1039), .C1(new_n1064), .C2(new_n792), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n782), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1065), .B1(new_n1001), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1037), .A2(new_n1067), .ZN(G387));
  AOI22_X1  g0868(.A1(new_n784), .A2(new_n719), .B1(new_n228), .B2(new_n216), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n243), .A2(new_n380), .ZN(new_n1070));
  AOI211_X1 g0870(.A(G45), .B(new_n719), .C1(G68), .C2(G77), .ZN(new_n1071));
  XOR2_X1   g0871(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n1072));
  OR3_X1    g0872(.A1(new_n1072), .A2(G50), .A3(new_n467), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1072), .B1(G50), .B2(new_n467), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1071), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n787), .A2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1069), .B1(new_n1070), .B2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1077), .A2(KEYINPUT113), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(KEYINPUT113), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n793), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n800), .A2(new_n357), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(G50), .B2(new_n806), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT115), .Z(new_n1083));
  OAI221_X1 g0883(.A(new_n1047), .B1(new_n203), .B2(new_n805), .C1(new_n815), .C2(new_n819), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n468), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1084), .B1(new_n1085), .B2(new_n811), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1043), .A2(G77), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n854), .B2(new_n814), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT114), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1083), .A2(new_n786), .A3(new_n1086), .A4(new_n1089), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G303), .A2(new_n804), .B1(new_n806), .B2(G317), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1091), .B1(new_n827), .B2(new_n810), .C1(new_n829), .C2(new_n819), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT116), .Z(new_n1093));
  INV_X1    g0893(.A(KEYINPUT48), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n835), .A2(G283), .B1(new_n1043), .B2(G294), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1097), .A2(KEYINPUT49), .A3(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n797), .A2(new_n570), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1100), .B(new_n786), .C1(G326), .C2(new_n831), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(KEYINPUT49), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1090), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT117), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n771), .B1(new_n1078), .B2(new_n1080), .C1(new_n1105), .C2(new_n840), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n1031), .B2(new_n782), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n770), .B2(new_n1034), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1034), .A2(new_n764), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1034), .A2(new_n764), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n717), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1108), .B1(new_n1109), .B2(new_n1111), .ZN(G393));
  NOR2_X1   g0912(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n711), .B1(new_n1021), .B2(new_n1025), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1110), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1115), .A2(new_n1035), .A3(new_n717), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n987), .A2(new_n782), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n793), .B1(new_n801), .B2(new_n217), .C1(new_n788), .C2(new_n250), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n771), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n796), .A2(new_n203), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n845), .B(new_n1121), .C1(G143), .C2(new_n831), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n786), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT118), .Z(new_n1124));
  OAI22_X1  g0924(.A1(new_n807), .A2(new_n815), .B1(new_n819), .B2(new_n854), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT51), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n811), .A2(G50), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n835), .A2(G77), .B1(new_n478), .B2(new_n804), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1124), .A2(new_n1126), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  OR2_X1    g0929(.A1(new_n1129), .A2(KEYINPUT119), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n820), .A2(G317), .B1(G311), .B2(new_n806), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT52), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n329), .B1(new_n814), .B2(new_n829), .C1(new_n805), .C2(new_n848), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n797), .A2(new_n228), .B1(new_n810), .B2(new_n1057), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n800), .A2(new_n570), .B1(new_n796), .B2(new_n1058), .ZN(new_n1135));
  OR4_X1    g0935(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1129), .A2(KEYINPUT119), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1130), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1120), .B1(new_n1138), .B2(new_n792), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1117), .A2(new_n770), .B1(new_n1118), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1116), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(KEYINPUT120), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT120), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1116), .A2(new_n1140), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1142), .A2(new_n1144), .ZN(G390));
  NAND2_X1  g0945(.A1(new_n935), .A2(G330), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n934), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n886), .A2(new_n869), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n958), .B1(new_n1150), .B2(new_n960), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n956), .B2(new_n957), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n958), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n869), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(new_n760), .B2(new_n868), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1153), .B1(new_n1155), .B2(new_n961), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n907), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n913), .B1(new_n1157), .B2(new_n922), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n955), .B1(new_n1158), .B2(KEYINPUT38), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1149), .B1(new_n1152), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1150), .A2(new_n960), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n1153), .ZN(new_n1163));
  AOI21_X1  g0963(.A(KEYINPUT38), .B1(new_n923), .B2(new_n924), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n954), .A2(new_n1164), .A3(new_n953), .ZN(new_n1165));
  AOI21_X1  g0965(.A(KEYINPUT39), .B1(new_n945), .B2(new_n925), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1163), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n752), .A2(new_n960), .A3(G330), .A4(new_n871), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1161), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1147), .A2(new_n567), .A3(new_n508), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1172), .B(new_n687), .C1(new_n763), .C2(new_n568), .ZN(new_n1173));
  OAI211_X1 g0973(.A(G330), .B(new_n871), .C1(new_n745), .C2(new_n751), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n961), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n1148), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n1150), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n961), .B1(new_n1146), .B2(new_n870), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1168), .A2(new_n1155), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1173), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1171), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1161), .A2(new_n1170), .A3(new_n1180), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1182), .A2(new_n717), .A3(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1161), .A2(new_n1170), .A3(new_n770), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n780), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n864), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n771), .B1(new_n1085), .B2(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(KEYINPUT54), .B(G143), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n807), .A2(new_n857), .B1(new_n805), .B2(new_n1189), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n329), .B(new_n1190), .C1(G125), .C2(new_n831), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n796), .A2(new_n854), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT53), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(G50), .A2(new_n833), .B1(new_n811), .B2(G137), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n835), .A2(G159), .B1(new_n820), .B2(G128), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1191), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G107), .A2(new_n811), .B1(new_n820), .B2(G283), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n835), .A2(G77), .B1(new_n833), .B2(G68), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n406), .B1(new_n804), .B2(G97), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n831), .A2(G294), .B1(new_n806), .B2(G116), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n860), .A2(new_n222), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1196), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1188), .B1(new_n1203), .B2(new_n792), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1186), .A2(new_n1204), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n1185), .A2(KEYINPUT121), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(KEYINPUT121), .B1(new_n1185), .B2(new_n1205), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1184), .B1(new_n1206), .B2(new_n1207), .ZN(G378));
  OAI21_X1  g1008(.A(new_n936), .B1(new_n954), .B2(new_n1164), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT40), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n894), .B1(new_n946), .B2(new_n948), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n686), .A2(new_n477), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n694), .B1(new_n498), .B2(new_n493), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1214), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n686), .A2(new_n477), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1215), .A2(new_n1217), .A3(new_n1219), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1211), .A2(new_n1212), .A3(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1223), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n964), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1223), .ZN(new_n1227));
  OAI21_X1  g1027(.A(G330), .B1(new_n1159), .B2(new_n947), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1227), .B1(new_n1228), .B2(new_n937), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1211), .A2(new_n1212), .A3(new_n1223), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1229), .A2(new_n959), .A3(new_n963), .A4(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1226), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1227), .A2(new_n780), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1187), .A2(G50), .ZN(new_n1234));
  INV_X1    g1034(.A(G125), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n1235), .A2(new_n819), .B1(new_n810), .B2(new_n857), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(G128), .A2(new_n806), .B1(new_n804), .B2(G137), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n796), .B2(new_n1189), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n1236), .B(new_n1238), .C1(G150), .C2(new_n835), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  OR2_X1    g1040(.A1(new_n1240), .A2(KEYINPUT59), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(KEYINPUT59), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n833), .A2(G159), .ZN(new_n1243));
  AOI211_X1 g1043(.A(G33), .B(G41), .C1(new_n831), .C2(G124), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .A4(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n833), .A2(G58), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n1246), .B1(new_n801), .B2(new_n810), .C1(new_n570), .C2(new_n819), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n358), .A2(new_n804), .B1(new_n806), .B2(G107), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n1058), .B2(new_n814), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1042), .A2(new_n1087), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1247), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n786), .A2(new_n395), .ZN(new_n1252));
  AND2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(KEYINPUT58), .ZN(new_n1254));
  OR2_X1    g1054(.A1(new_n1253), .A2(KEYINPUT58), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n207), .B1(G33), .B2(G41), .C1(new_n786), .C2(new_n395), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1245), .A2(new_n1254), .A3(new_n1255), .A4(new_n1256), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n772), .B(new_n1234), .C1(new_n1257), .C2(new_n792), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1232), .A2(new_n770), .B1(new_n1233), .B2(new_n1258), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1224), .A2(new_n1225), .A3(new_n964), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1229), .A2(new_n1230), .B1(new_n959), .B2(new_n963), .ZN(new_n1261));
  OAI21_X1  g1061(.A(KEYINPUT57), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1173), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1183), .A2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n717), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1183), .A2(new_n1263), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT57), .B1(new_n1232), .B2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1259), .B1(new_n1265), .B2(new_n1267), .ZN(G375));
  NOR2_X1   g1068(.A1(new_n1180), .A2(new_n1015), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1269), .B1(new_n1263), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n961), .A2(new_n780), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n771), .B1(new_n1187), .B2(G68), .ZN(new_n1273));
  OAI22_X1  g1073(.A1(new_n800), .A2(new_n207), .B1(new_n805), .B2(new_n854), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1274), .B(KEYINPUT123), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n831), .A2(G128), .B1(new_n806), .B2(G137), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1246), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n857), .A2(new_n819), .B1(new_n810), .B2(new_n1189), .ZN(new_n1278));
  NOR3_X1   g1078(.A1(new_n1277), .A2(new_n515), .A3(new_n1278), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1275), .B(new_n1279), .C1(new_n815), .C2(new_n860), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n819), .A2(new_n848), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n1281), .B(new_n1081), .C1(G116), .C2(new_n811), .ZN(new_n1282));
  OAI22_X1  g1082(.A1(new_n807), .A2(new_n1058), .B1(new_n814), .B2(new_n1057), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1283), .B1(G107), .B2(new_n804), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1282), .B(new_n1284), .C1(new_n801), .C2(new_n860), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n329), .B1(new_n797), .B2(new_n226), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(new_n1286), .B(KEYINPUT122), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1280), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1273), .B1(new_n1288), .B2(new_n792), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n1270), .A2(new_n770), .B1(new_n1272), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1271), .A2(new_n1290), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1291), .B(KEYINPUT124), .ZN(G381));
  NOR4_X1   g1092(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1185), .A2(new_n1205), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1184), .A2(new_n1295), .ZN(new_n1296));
  AND4_X1   g1096(.A1(new_n1037), .A2(new_n1067), .A3(new_n1142), .A4(new_n1144), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1293), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  OR2_X1    g1098(.A1(new_n1298), .A2(G375), .ZN(G407));
  NAND2_X1  g1099(.A1(new_n1296), .A2(new_n695), .ZN(new_n1300));
  OAI211_X1 g1100(.A(G407), .B(G213), .C1(G375), .C2(new_n1300), .ZN(G409));
  XNOR2_X1  g1101(.A(G393), .B(G396), .ZN(new_n1302));
  AOI22_X1  g1102(.A1(new_n1037), .A2(new_n1067), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1302), .B1(new_n1297), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(G387), .A2(G390), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1302), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1037), .A2(new_n1142), .A3(new_n1067), .A4(new_n1144), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1305), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1304), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT61), .ZN(new_n1310));
  AND2_X1   g1110(.A1(new_n695), .A2(G213), .ZN(new_n1311));
  OAI211_X1 g1111(.A(G378), .B(new_n1259), .C1(new_n1265), .C2(new_n1267), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1232), .A2(new_n1266), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1313), .A2(new_n1015), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1232), .A2(new_n770), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1233), .A2(new_n1258), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1296), .B1(new_n1314), .B2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1311), .B1(new_n1312), .B2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT60), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1320), .B1(new_n1270), .B2(new_n1263), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1177), .A2(new_n1173), .A3(new_n1179), .A4(KEYINPUT60), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1321), .A2(new_n1181), .A3(new_n717), .A4(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(new_n1290), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT125), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(G384), .A2(new_n1325), .ZN(new_n1326));
  OAI211_X1 g1126(.A(KEYINPUT125), .B(new_n872), .C1(new_n890), .C2(new_n891), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1324), .A2(new_n1326), .A3(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(G384), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1329), .A2(new_n1323), .A3(KEYINPUT125), .A4(new_n1290), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1328), .A2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1311), .A2(G2897), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1328), .A2(new_n1330), .A3(G2897), .A4(new_n1311), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1310), .B1(new_n1319), .B2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT62), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1337), .B1(new_n1319), .B2(new_n1331), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1336), .A2(new_n1338), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1319), .A2(new_n1337), .A3(new_n1331), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1309), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  OAI211_X1 g1141(.A(new_n1309), .B(new_n1310), .C1(new_n1319), .C2(new_n1335), .ZN(new_n1342));
  AOI21_X1  g1142(.A(KEYINPUT63), .B1(new_n1319), .B2(new_n1331), .ZN(new_n1343));
  AND3_X1   g1143(.A1(new_n1319), .A2(KEYINPUT63), .A3(new_n1331), .ZN(new_n1344));
  NOR3_X1   g1144(.A1(new_n1342), .A2(new_n1343), .A3(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(KEYINPUT126), .B1(new_n1341), .B2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1336), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1343), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1319), .A2(KEYINPUT63), .A3(new_n1331), .ZN(new_n1349));
  NAND4_X1  g1149(.A1(new_n1347), .A2(new_n1348), .A3(new_n1309), .A4(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT126), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1340), .ZN(new_n1352));
  NOR3_X1   g1152(.A1(new_n1352), .A2(new_n1336), .A3(new_n1338), .ZN(new_n1353));
  OAI211_X1 g1153(.A(new_n1350), .B(new_n1351), .C1(new_n1353), .C2(new_n1309), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1346), .A2(new_n1354), .ZN(G405));
  NAND2_X1  g1155(.A1(G375), .A2(new_n1296), .ZN(new_n1356));
  AOI21_X1  g1156(.A(KEYINPUT127), .B1(new_n1356), .B2(new_n1312), .ZN(new_n1357));
  NOR2_X1   g1157(.A1(new_n1357), .A2(new_n1331), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1356), .A2(KEYINPUT127), .A3(new_n1312), .ZN(new_n1359));
  OR2_X1    g1159(.A1(new_n1358), .A2(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1358), .A2(new_n1359), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1360), .A2(new_n1361), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1362), .A2(new_n1309), .ZN(new_n1363));
  NAND4_X1  g1163(.A1(new_n1360), .A2(new_n1308), .A3(new_n1304), .A4(new_n1361), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1363), .A2(new_n1364), .ZN(G402));
endmodule


