//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 0 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  AOI21_X1  g004(.A(KEYINPUT16), .B1(new_n190), .B2(G125), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT82), .ZN(new_n192));
  INV_X1    g006(.A(G125), .ZN(new_n193));
  OAI211_X1 g007(.A(new_n192), .B(G140), .C1(new_n193), .C2(KEYINPUT81), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT82), .B1(new_n190), .B2(G125), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT81), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(new_n190), .A3(G125), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n195), .A3(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n191), .B1(new_n198), .B2(KEYINPUT16), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  OR2_X1    g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G125), .B(G140), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(new_n200), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n204));
  INV_X1    g018(.A(G119), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G128), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT23), .A3(G119), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n206), .B(new_n208), .C1(G119), .C2(new_n207), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT83), .B(G110), .ZN(new_n210));
  XNOR2_X1  g024(.A(G119), .B(G128), .ZN(new_n211));
  XOR2_X1   g025(.A(KEYINPUT24), .B(G110), .Z(new_n212));
  OAI22_X1  g026(.A1(new_n209), .A2(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n201), .A2(new_n203), .A3(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n199), .B(new_n200), .ZN(new_n215));
  INV_X1    g029(.A(G110), .ZN(new_n216));
  XOR2_X1   g030(.A(new_n209), .B(KEYINPUT80), .Z(new_n217));
  OAI21_X1  g031(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n212), .A2(new_n211), .ZN(new_n219));
  XOR2_X1   g033(.A(new_n219), .B(KEYINPUT79), .Z(new_n220));
  OAI21_X1  g034(.A(new_n214), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G953), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(G221), .A3(G234), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n223), .B(KEYINPUT22), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n224), .B(G137), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n221), .B(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT25), .ZN(new_n228));
  NOR3_X1   g042(.A1(new_n227), .A2(new_n228), .A3(G902), .ZN(new_n229));
  AOI21_X1  g043(.A(KEYINPUT25), .B1(new_n226), .B2(new_n188), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n189), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n189), .A2(G902), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n226), .A2(new_n232), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT74), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT32), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT73), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT66), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n239));
  INV_X1    g053(.A(G134), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n239), .B1(new_n240), .B2(G137), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT11), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(G137), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT11), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n239), .B(new_n244), .C1(new_n240), .C2(G137), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G131), .ZN(new_n247));
  INV_X1    g061(.A(G131), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n242), .A2(new_n248), .A3(new_n243), .A4(new_n245), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G143), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n251), .A2(G146), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(KEYINPUT64), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT64), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G143), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n252), .B1(new_n256), .B2(G146), .ZN(new_n257));
  AND2_X1   g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n253), .A2(new_n255), .A3(new_n200), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n200), .A2(G143), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(KEYINPUT0), .A2(G128), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n257), .A2(new_n258), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n243), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n240), .A2(G137), .ZN(new_n267));
  OAI21_X1  g081(.A(G131), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n249), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n252), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n207), .A2(KEYINPUT1), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT64), .B(G143), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n270), .B(new_n271), .C1(new_n272), .C2(new_n200), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n260), .B1(new_n272), .B2(new_n200), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT1), .B1(new_n251), .B2(G146), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G128), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n273), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n250), .A2(new_n265), .B1(new_n269), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n238), .B1(new_n279), .B2(KEYINPUT30), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT30), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n270), .B(new_n258), .C1(new_n272), .C2(new_n200), .ZN(new_n282));
  INV_X1    g096(.A(new_n264), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n282), .B1(new_n274), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n284), .B1(new_n247), .B2(new_n249), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n249), .A2(new_n268), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n262), .A2(new_n276), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n286), .B1(new_n287), .B2(new_n273), .ZN(new_n288));
  OAI211_X1 g102(.A(KEYINPUT66), .B(new_n281), .C1(new_n285), .C2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n280), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n200), .B1(new_n253), .B2(new_n255), .ZN(new_n291));
  INV_X1    g105(.A(new_n271), .ZN(new_n292));
  NOR3_X1   g106(.A1(new_n291), .A2(new_n252), .A3(new_n292), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n259), .A2(new_n261), .B1(G128), .B2(new_n275), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT70), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT70), .B1(new_n287), .B2(new_n273), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n269), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n250), .A2(new_n265), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(KEYINPUT30), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT71), .ZN(new_n301));
  NOR2_X1   g115(.A1(KEYINPUT2), .A2(G113), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT69), .ZN(new_n304));
  NAND2_X1  g118(.A1(KEYINPUT2), .A2(G113), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n305), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT69), .B1(new_n307), .B2(new_n302), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT68), .ZN(new_n310));
  INV_X1    g124(.A(G116), .ZN(new_n311));
  NOR3_X1   g125(.A1(new_n310), .A2(new_n311), .A3(G119), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n311), .A2(G119), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT68), .B1(new_n205), .B2(G116), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n312), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT67), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n309), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n313), .A2(KEYINPUT68), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n310), .B1(new_n311), .B2(G119), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n319), .B1(new_n313), .B2(new_n320), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n321), .A2(KEYINPUT67), .A3(new_n308), .A4(new_n306), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n295), .B1(new_n293), .B2(new_n294), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n287), .A2(KEYINPUT70), .A3(new_n273), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n326), .A2(new_n269), .B1(new_n250), .B2(new_n265), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT71), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(new_n328), .A3(KEYINPUT30), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n290), .A2(new_n301), .A3(new_n323), .A4(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n323), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n298), .A2(new_n299), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT72), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n327), .A2(KEYINPUT72), .A3(new_n331), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G237), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(new_n222), .A3(G210), .ZN(new_n338));
  XOR2_X1   g152(.A(new_n338), .B(KEYINPUT27), .Z(new_n339));
  XNOR2_X1  g153(.A(new_n339), .B(KEYINPUT26), .ZN(new_n340));
  INV_X1    g154(.A(G101), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n340), .B(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n330), .A2(new_n336), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT31), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n330), .A2(KEYINPUT31), .A3(new_n336), .A4(new_n342), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT28), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n332), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n279), .A2(new_n331), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n350), .B1(new_n334), .B2(new_n335), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n349), .B1(new_n351), .B2(new_n348), .ZN(new_n352));
  INV_X1    g166(.A(new_n342), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n347), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(G472), .A2(G902), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n237), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n345), .A2(new_n346), .B1(new_n353), .B2(new_n352), .ZN(new_n358));
  INV_X1    g172(.A(new_n356), .ZN(new_n359));
  NOR3_X1   g173(.A1(new_n358), .A2(KEYINPUT73), .A3(new_n359), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n235), .B(new_n236), .C1(new_n357), .C2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n355), .A2(new_n237), .A3(new_n356), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT73), .B1(new_n358), .B2(new_n359), .ZN(new_n363));
  AOI21_X1  g177(.A(KEYINPUT32), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n358), .A2(new_n359), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT74), .B1(new_n365), .B2(KEYINPUT32), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n361), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT77), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n349), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(KEYINPUT28), .B1(new_n327), .B2(new_n331), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n370), .A2(KEYINPUT77), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT72), .B1(new_n327), .B2(new_n331), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n286), .B1(new_n324), .B2(new_n325), .ZN(new_n373));
  NOR4_X1   g187(.A1(new_n373), .A2(new_n285), .A3(new_n333), .A4(new_n323), .ZN(new_n374));
  OAI22_X1  g188(.A1(new_n372), .A2(new_n374), .B1(new_n327), .B2(new_n331), .ZN(new_n375));
  AOI211_X1 g189(.A(new_n369), .B(new_n371), .C1(new_n375), .C2(KEYINPUT28), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT29), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n353), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(G902), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n330), .A2(new_n336), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n353), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT76), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n380), .A2(KEYINPUT76), .A3(new_n353), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n342), .B(new_n349), .C1(new_n351), .C2(new_n348), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT75), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n383), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n377), .B1(new_n385), .B2(KEYINPUT75), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n379), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n389), .A2(KEYINPUT78), .A3(G472), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT78), .B1(new_n389), .B2(G472), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n234), .B1(new_n367), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(G214), .B1(G237), .B2(G902), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G952), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n396), .A2(KEYINPUT101), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n396), .A2(KEYINPUT101), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n222), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n399), .B1(G234), .B2(G237), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT21), .B(G898), .ZN(new_n401));
  AOI211_X1 g215(.A(new_n188), .B(new_n222), .C1(G234), .C2(G237), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n265), .A2(new_n193), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n278), .A2(G125), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G224), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n407), .A2(G953), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n406), .B(new_n409), .ZN(new_n410));
  XOR2_X1   g224(.A(G110), .B(G122), .Z(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G104), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT3), .B1(new_n413), .B2(G107), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT3), .ZN(new_n415));
  INV_X1    g229(.A(G107), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n416), .A3(G104), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n413), .A2(G107), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n414), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  XOR2_X1   g233(.A(KEYINPUT86), .B(KEYINPUT4), .Z(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(G101), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n419), .A2(G101), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT84), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n414), .A2(new_n417), .A3(new_n341), .A4(new_n418), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n424), .A2(KEYINPUT85), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(KEYINPUT85), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n423), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT4), .B1(new_n422), .B2(KEYINPUT84), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n323), .B(new_n421), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n414), .A2(new_n417), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT85), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n430), .A2(new_n431), .A3(new_n341), .A4(new_n418), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n424), .A2(KEYINPUT85), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n416), .A2(G104), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n418), .A2(new_n434), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n432), .A2(new_n433), .B1(G101), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G113), .ZN(new_n437));
  XOR2_X1   g251(.A(KEYINPUT94), .B(KEYINPUT5), .Z(new_n438));
  AOI21_X1  g252(.A(new_n437), .B1(new_n438), .B2(new_n313), .ZN(new_n439));
  XNOR2_X1  g253(.A(KEYINPUT94), .B(KEYINPUT5), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n319), .B(new_n440), .C1(new_n313), .C2(new_n320), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT95), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n316), .A2(new_n303), .A3(new_n305), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n439), .A2(new_n441), .A3(KEYINPUT95), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n436), .A2(new_n444), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n412), .B1(new_n429), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT6), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT97), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT97), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n448), .A2(new_n452), .A3(new_n449), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n429), .A2(new_n412), .A3(new_n447), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(new_n448), .ZN(new_n456));
  AOI21_X1  g270(.A(KEYINPUT96), .B1(new_n456), .B2(KEYINPUT6), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT96), .ZN(new_n458));
  NOR4_X1   g272(.A1(new_n455), .A2(new_n448), .A3(new_n458), .A4(new_n449), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n410), .B(new_n454), .C1(new_n457), .C2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n406), .A2(KEYINPUT7), .A3(new_n409), .ZN(new_n461));
  XOR2_X1   g275(.A(new_n461), .B(KEYINPUT99), .Z(new_n462));
  NAND2_X1  g276(.A1(new_n316), .A2(KEYINPUT5), .ZN(new_n463));
  XOR2_X1   g277(.A(new_n463), .B(KEYINPUT98), .Z(new_n464));
  INV_X1    g278(.A(new_n439), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n445), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n436), .ZN(new_n467));
  XOR2_X1   g281(.A(new_n411), .B(KEYINPUT8), .Z(new_n468));
  NAND3_X1  g282(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n467), .B(new_n468), .C1(new_n436), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n409), .A2(KEYINPUT7), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n471), .B1(new_n404), .B2(new_n405), .ZN(new_n472));
  INV_X1    g286(.A(new_n455), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n462), .A2(new_n470), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n460), .A2(new_n188), .A3(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(G210), .B1(G237), .B2(G902), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n460), .A2(new_n188), .A3(new_n476), .A4(new_n474), .ZN(new_n479));
  AOI211_X1 g293(.A(new_n395), .B(new_n403), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n199), .B(G146), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n251), .A2(new_n337), .A3(new_n222), .A4(G214), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n337), .A2(new_n222), .A3(G214), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n482), .B1(new_n256), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n484), .A2(new_n248), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT17), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n484), .B(new_n248), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n481), .B(new_n486), .C1(KEYINPUT17), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n485), .A2(KEYINPUT18), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n198), .A2(G146), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n203), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT18), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n484), .B1(new_n492), .B2(new_n248), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n489), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(G113), .B(G122), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(new_n413), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n488), .A2(new_n497), .A3(new_n494), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n188), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(G475), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n198), .A2(KEYINPUT19), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n202), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n487), .B(new_n201), .C1(G146), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n494), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n498), .ZN(new_n510));
  AOI21_X1  g324(.A(G475), .B1(new_n500), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n188), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n512), .A2(KEYINPUT20), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT20), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n514), .B1(new_n511), .B2(new_n188), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n503), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT13), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n256), .A2(new_n518), .A3(G128), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n207), .A2(G143), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n520), .B1(new_n272), .B2(new_n207), .ZN(new_n521));
  OAI211_X1 g335(.A(G134), .B(new_n519), .C1(new_n521), .C2(new_n518), .ZN(new_n522));
  XNOR2_X1  g336(.A(G116), .B(G122), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n523), .B(new_n416), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n522), .B(new_n524), .C1(G134), .C2(new_n521), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n521), .B(new_n240), .ZN(new_n526));
  OR2_X1    g340(.A1(new_n311), .A2(G122), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n416), .B1(new_n527), .B2(KEYINPUT14), .ZN(new_n528));
  XOR2_X1   g342(.A(new_n528), .B(new_n523), .Z(new_n529));
  OAI21_X1  g343(.A(new_n525), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  XOR2_X1   g344(.A(KEYINPUT9), .B(G234), .Z(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n532), .A2(new_n187), .A3(G953), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n530), .A2(new_n534), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n188), .ZN(new_n539));
  INV_X1    g353(.A(G478), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n540), .A2(KEYINPUT15), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n539), .B(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n480), .A2(new_n517), .A3(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(G221), .B1(new_n532), .B2(G902), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n326), .A2(KEYINPUT10), .A3(new_n436), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n432), .A2(new_n433), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n207), .B1(new_n259), .B2(KEYINPUT1), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n273), .B1(new_n549), .B2(new_n257), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n435), .A2(G101), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  XOR2_X1   g366(.A(KEYINPUT87), .B(KEYINPUT10), .Z(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT88), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT88), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n552), .A2(new_n557), .A3(new_n554), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n547), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT89), .ZN(new_n560));
  INV_X1    g374(.A(new_n250), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n265), .B(new_n421), .C1(new_n427), .C2(new_n428), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n559), .A2(new_n560), .A3(new_n561), .A4(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n326), .A2(KEYINPUT10), .A3(new_n436), .ZN(new_n564));
  AOI211_X1 g378(.A(KEYINPUT88), .B(new_n553), .C1(new_n436), .C2(new_n550), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n557), .B1(new_n552), .B2(new_n554), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n562), .B(new_n564), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT89), .B1(new_n567), .B2(new_n250), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(G110), .B(G140), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n222), .A2(G227), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n570), .B(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT92), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n567), .A2(new_n250), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n569), .A2(KEYINPUT92), .A3(new_n572), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  OR2_X1    g392(.A1(new_n436), .A2(new_n278), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n561), .B1(new_n579), .B2(new_n552), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT90), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT91), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT91), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT12), .B1(new_n580), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g399(.A1(new_n563), .A2(new_n568), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n582), .A2(KEYINPUT91), .A3(KEYINPUT12), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n572), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n578), .A2(G469), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(G469), .A2(G902), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n583), .A2(new_n585), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n569), .A2(new_n572), .A3(new_n593), .A4(new_n587), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT93), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n569), .A2(new_n576), .ZN(new_n596));
  INV_X1    g410(.A(new_n572), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT93), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n586), .A2(new_n599), .A3(new_n572), .A4(new_n587), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n595), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(G469), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n602), .A3(new_n188), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n546), .B1(new_n592), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n544), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n393), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(new_n341), .ZN(G3));
  INV_X1    g421(.A(new_n480), .ZN(new_n608));
  OR2_X1    g422(.A1(new_n537), .A2(KEYINPUT33), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n537), .A2(KEYINPUT33), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n609), .A2(G478), .A3(new_n188), .A4(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n539), .A2(new_n540), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n516), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n608), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n362), .A2(new_n363), .ZN(new_n616));
  OAI21_X1  g430(.A(G472), .B1(new_n358), .B2(G902), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n616), .A2(new_n234), .A3(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n615), .A2(new_n604), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT34), .B(G104), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G6));
  NAND2_X1  g436(.A1(new_n503), .A2(KEYINPUT102), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT102), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n502), .A2(new_n624), .A3(G475), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n512), .B(KEYINPUT20), .ZN(new_n627));
  INV_X1    g441(.A(new_n403), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n626), .A2(new_n627), .A3(new_n542), .A4(new_n628), .ZN(new_n629));
  OR2_X1    g443(.A1(new_n629), .A2(KEYINPUT103), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n395), .B1(new_n478), .B2(new_n479), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(KEYINPUT103), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n633), .A2(new_n604), .A3(new_n619), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT35), .B(G107), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G9));
  NAND2_X1  g450(.A1(new_n616), .A2(new_n617), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n232), .ZN(new_n639));
  INV_X1    g453(.A(new_n225), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(KEYINPUT36), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n221), .B(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n231), .B1(new_n639), .B2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n544), .A2(new_n604), .A3(new_n638), .A4(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT104), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT37), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(new_n216), .ZN(G12));
  INV_X1    g462(.A(KEYINPUT78), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n371), .B1(new_n375), .B2(KEYINPUT28), .ZN(new_n650));
  INV_X1    g464(.A(new_n369), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n378), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n188), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT75), .ZN(new_n655));
  INV_X1    g469(.A(new_n350), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n656), .B1(new_n372), .B2(new_n374), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n370), .B1(new_n657), .B2(KEYINPUT28), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n655), .B1(new_n658), .B2(new_n342), .ZN(new_n659));
  AOI21_X1  g473(.A(KEYINPUT76), .B1(new_n380), .B2(new_n353), .ZN(new_n660));
  AOI211_X1 g474(.A(new_n382), .B(new_n342), .C1(new_n330), .C2(new_n336), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n388), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n654), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(G472), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n649), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n389), .A2(KEYINPUT78), .A3(G472), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n236), .B1(new_n357), .B2(new_n360), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n365), .A2(KEYINPUT32), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n235), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n668), .A2(new_n672), .A3(new_n361), .ZN(new_n673));
  INV_X1    g487(.A(G900), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n400), .B1(new_n674), .B2(new_n402), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  AND4_X1   g490(.A1(new_n627), .A2(new_n626), .A3(new_n542), .A4(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n631), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT105), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n631), .A2(new_n677), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n673), .A2(new_n682), .A3(new_n604), .A4(new_n644), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G128), .ZN(G30));
  XNOR2_X1  g498(.A(new_n675), .B(KEYINPUT39), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n604), .A2(new_n686), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n687), .A2(KEYINPUT40), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(KEYINPUT40), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n478), .A2(new_n479), .ZN(new_n690));
  XOR2_X1   g504(.A(new_n690), .B(KEYINPUT38), .Z(new_n691));
  NOR2_X1   g505(.A1(new_n543), .A2(new_n517), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n691), .A2(new_n395), .A3(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n688), .A2(new_n689), .A3(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n343), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n696), .B1(new_n353), .B2(new_n375), .ZN(new_n697));
  OAI21_X1  g511(.A(G472), .B1(new_n697), .B2(G902), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n672), .A2(new_n361), .A3(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n644), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n695), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n256), .ZN(G45));
  NAND4_X1  g517(.A1(new_n673), .A2(new_n604), .A3(new_n631), .A4(new_n644), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n613), .A2(new_n516), .A3(new_n676), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n200), .ZN(G48));
  NAND2_X1  g521(.A1(new_n601), .A2(new_n188), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(G469), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n603), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n710), .A2(new_n546), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n673), .A2(new_n234), .A3(new_n615), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT41), .B(G113), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT106), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n712), .B(new_n714), .ZN(G15));
  NAND4_X1  g529(.A1(new_n673), .A2(new_n234), .A3(new_n633), .A4(new_n711), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  NAND4_X1  g531(.A1(new_n673), .A2(new_n544), .A3(new_n644), .A4(new_n711), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G119), .ZN(G21));
  INV_X1    g533(.A(new_n234), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n347), .B1(new_n376), .B2(new_n342), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n356), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n617), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n711), .A2(new_n724), .A3(new_n480), .A4(new_n692), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n705), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n613), .A2(new_n516), .A3(KEYINPUT107), .A4(new_n676), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n731), .A2(new_n700), .A3(new_n723), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n711), .A3(new_n631), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G125), .ZN(G27));
  OAI21_X1  g548(.A(new_n236), .B1(new_n358), .B2(new_n359), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n668), .A2(new_n670), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n234), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n603), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n590), .A2(new_n591), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n545), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(KEYINPUT108), .B1(new_n690), .B2(new_n395), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n478), .A2(new_n743), .A3(new_n394), .A4(new_n479), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n730), .A2(KEYINPUT42), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n741), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n741), .A2(new_n745), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n748), .A2(new_n673), .A3(new_n234), .A4(new_n730), .ZN(new_n749));
  XOR2_X1   g563(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n750));
  AOI22_X1  g564(.A1(new_n738), .A2(new_n747), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n248), .ZN(G33));
  AND4_X1   g566(.A1(new_n673), .A2(new_n748), .A3(new_n234), .A4(new_n677), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n240), .ZN(G36));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n755));
  AOI21_X1  g569(.A(KEYINPUT92), .B1(new_n569), .B2(new_n572), .ZN(new_n756));
  AOI211_X1 g570(.A(new_n574), .B(new_n597), .C1(new_n563), .C2(new_n568), .ZN(new_n757));
  INV_X1    g571(.A(new_n576), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n755), .B1(new_n759), .B2(new_n588), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n578), .A2(KEYINPUT45), .A3(new_n589), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(G469), .A3(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(KEYINPUT46), .A3(new_n591), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT110), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n764), .A3(new_n603), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n764), .B1(new_n763), .B2(new_n603), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n762), .A2(new_n591), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT46), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n546), .B1(new_n768), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n517), .A2(new_n613), .ZN(new_n773));
  XOR2_X1   g587(.A(new_n773), .B(KEYINPUT43), .Z(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(new_n637), .A3(new_n644), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT44), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n775), .B(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n745), .B(KEYINPUT111), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n772), .A2(new_n686), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G137), .ZN(G39));
  NAND2_X1  g595(.A1(new_n763), .A2(new_n603), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT110), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n771), .A3(new_n765), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n545), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT47), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT112), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n786), .A2(KEYINPUT112), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n673), .A2(new_n234), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n790), .B1(new_n784), .B2(new_n545), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n745), .A2(new_n705), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n791), .A2(new_n792), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G140), .ZN(G42));
  NAND2_X1  g611(.A1(new_n710), .A2(KEYINPUT49), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n798), .A2(new_n234), .A3(new_n545), .A4(new_n394), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n710), .A2(KEYINPUT49), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n799), .A2(new_n773), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n699), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(new_n802), .A3(new_n691), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n683), .B(new_n733), .C1(new_n704), .C2(new_n705), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n741), .A2(new_n675), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n692), .A2(new_n690), .A3(new_n394), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n805), .A2(new_n700), .A3(new_n699), .A4(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(KEYINPUT52), .B1(new_n804), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n683), .A2(new_n733), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n604), .B(new_n644), .C1(new_n367), .C2(new_n392), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n705), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n631), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n811), .A2(new_n815), .A3(new_n816), .A4(new_n807), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n809), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n749), .A2(new_n750), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n747), .A2(new_n234), .A3(new_n736), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n753), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n543), .A2(new_n676), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n742), .A2(new_n744), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(new_n627), .A3(new_n626), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n812), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT113), .ZN(new_n826));
  INV_X1    g640(.A(new_n614), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n826), .B1(new_n480), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n542), .A2(new_n627), .A3(new_n503), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n829), .B1(new_n614), .B2(KEYINPUT113), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n830), .A2(new_n631), .A3(new_n628), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n604), .B(new_n619), .C1(new_n828), .C2(new_n831), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n645), .B(new_n832), .C1(new_n393), .C2(new_n605), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n825), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n748), .A2(new_n732), .ZN(new_n835));
  AND4_X1   g649(.A1(new_n712), .A2(new_n716), .A3(new_n718), .A4(new_n725), .ZN(new_n836));
  AND4_X1   g650(.A1(new_n821), .A2(new_n834), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n818), .A2(new_n837), .A3(KEYINPUT53), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n809), .A2(new_n817), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n821), .A2(new_n834), .A3(new_n835), .A4(new_n836), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT54), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n838), .A2(new_n845), .A3(new_n842), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n774), .A2(new_n400), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n848), .A2(new_n711), .A3(new_n724), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n631), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n848), .A2(new_n711), .A3(new_n823), .ZN(new_n851));
  XOR2_X1   g665(.A(new_n851), .B(KEYINPUT115), .Z(new_n852));
  AND2_X1   g666(.A1(new_n852), .A2(new_n738), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n853), .A2(KEYINPUT48), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(KEYINPUT48), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n711), .A2(new_n823), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n234), .A2(new_n400), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n856), .A2(new_n699), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n399), .B1(new_n858), .B2(new_n827), .ZN(new_n859));
  AND4_X1   g673(.A1(new_n850), .A2(new_n854), .A3(new_n855), .A4(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n847), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n858), .A2(new_n517), .A3(new_n612), .A4(new_n611), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n862), .A2(KEYINPUT116), .ZN(new_n863));
  INV_X1    g677(.A(new_n723), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n852), .A2(new_n644), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n862), .A2(KEYINPUT116), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n849), .A2(new_n395), .A3(new_n691), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n867), .A2(KEYINPUT50), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n863), .A2(new_n865), .A3(new_n866), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n867), .A2(KEYINPUT50), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n848), .A2(new_n724), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n789), .B1(new_n785), .B2(new_n787), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n793), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n710), .A2(new_n545), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n779), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n869), .B(new_n870), .C1(new_n871), .C2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT51), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n876), .A2(KEYINPUT114), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n877), .B1(new_n876), .B2(KEYINPUT114), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n861), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(G952), .A2(G953), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n803), .B1(new_n880), .B2(new_n881), .ZN(G75));
  NAND2_X1  g696(.A1(new_n396), .A2(G953), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT117), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT53), .B1(new_n818), .B2(new_n837), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n840), .A2(new_n841), .A3(new_n839), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(new_n188), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT56), .B1(new_n889), .B2(G210), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n454), .B1(new_n457), .B2(new_n459), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(new_n410), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT55), .Z(new_n893));
  OR2_X1    g707(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n890), .A2(new_n893), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n885), .B1(new_n894), .B2(new_n895), .ZN(G51));
  NOR3_X1   g710(.A1(new_n888), .A2(new_n188), .A3(new_n762), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT119), .Z(new_n898));
  NAND3_X1  g712(.A1(new_n844), .A2(KEYINPUT118), .A3(new_n846), .ZN(new_n899));
  OR3_X1    g713(.A1(new_n843), .A2(KEYINPUT118), .A3(KEYINPUT54), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n591), .B(KEYINPUT57), .Z(new_n901));
  NAND3_X1  g715(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n601), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n885), .B1(new_n898), .B2(new_n903), .ZN(G54));
  NAND3_X1  g718(.A1(new_n889), .A2(KEYINPUT58), .A3(G475), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n500), .A2(new_n510), .ZN(new_n906));
  OR2_X1    g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n905), .A2(new_n906), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n885), .B1(new_n907), .B2(new_n908), .ZN(G60));
  INV_X1    g723(.A(KEYINPUT120), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n609), .A2(new_n610), .ZN(new_n911));
  NAND2_X1  g725(.A1(G478), .A2(G902), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT59), .Z(new_n913));
  NOR2_X1   g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n899), .A2(new_n900), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n913), .B1(new_n844), .B2(new_n846), .ZN(new_n916));
  INV_X1    g730(.A(new_n911), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n884), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n910), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n911), .B1(new_n847), .B2(new_n913), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n899), .A2(new_n900), .A3(new_n914), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n920), .A2(KEYINPUT120), .A3(new_n884), .A4(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n919), .A2(new_n922), .ZN(G63));
  NAND2_X1  g737(.A1(G217), .A2(G902), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT60), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n886), .B2(new_n887), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n885), .B1(new_n927), .B2(new_n227), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT121), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT61), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n925), .B1(new_n838), .B2(new_n842), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n884), .B1(new_n931), .B2(new_n226), .ZN(new_n932));
  AOI211_X1 g746(.A(new_n643), .B(new_n925), .C1(new_n838), .C2(new_n842), .ZN(new_n933));
  OAI21_X1  g747(.A(KEYINPUT122), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n933), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT122), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n928), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n930), .A2(new_n934), .A3(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT61), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n929), .B(new_n884), .C1(new_n931), .C2(new_n226), .ZN(new_n940));
  AOI22_X1  g754(.A1(new_n937), .A2(new_n934), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n938), .A2(new_n941), .ZN(G66));
  INV_X1    g756(.A(new_n833), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n836), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT123), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n222), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT124), .Z(new_n947));
  OAI21_X1  g761(.A(G953), .B1(new_n401), .B2(new_n407), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n891), .B1(G898), .B2(new_n222), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n949), .B(new_n950), .ZN(G69));
  AOI21_X1  g765(.A(new_n222), .B1(G227), .B2(G900), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n290), .A2(new_n301), .A3(new_n329), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(new_n507), .ZN(new_n954));
  INV_X1    g768(.A(new_n804), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n784), .A2(new_n545), .A3(new_n686), .A4(new_n806), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n821), .B(new_n955), .C1(new_n956), .C2(new_n737), .ZN(new_n957));
  INV_X1    g771(.A(new_n779), .ZN(new_n958));
  NOR4_X1   g772(.A1(new_n785), .A2(new_n777), .A3(new_n958), .A4(new_n685), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(G953), .B1(new_n960), .B2(new_n796), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n222), .A2(G900), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n792), .ZN(new_n965));
  INV_X1    g779(.A(new_n795), .ZN(new_n966));
  NOR4_X1   g780(.A1(new_n872), .A2(new_n965), .A3(new_n793), .A4(new_n966), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n751), .A2(new_n804), .A3(new_n753), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n772), .A2(new_n686), .A3(new_n738), .A4(new_n806), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n968), .A2(new_n780), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n222), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n963), .ZN(new_n972));
  AOI21_X1  g786(.A(KEYINPUT126), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n954), .B1(new_n964), .B2(new_n973), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n829), .A2(new_n614), .ZN(new_n975));
  NOR4_X1   g789(.A1(new_n393), .A2(new_n687), .A3(new_n745), .A4(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT62), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n977), .B1(new_n702), .B2(new_n804), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n955), .B(KEYINPUT62), .C1(new_n701), .C2(new_n695), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n976), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n980), .A2(new_n780), .A3(new_n796), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n954), .A2(G953), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n974), .A2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT125), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n952), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n954), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n962), .B1(new_n961), .B2(new_n963), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n971), .A2(KEYINPUT126), .A3(new_n972), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n987), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n983), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n985), .B(new_n952), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n986), .A2(new_n993), .ZN(G72));
  NAND2_X1  g808(.A1(G472), .A2(G902), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT63), .Z(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(KEYINPUT127), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n997), .B1(new_n981), .B2(new_n945), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n998), .A2(new_n342), .ZN(new_n999));
  OR3_X1    g813(.A1(new_n945), .A2(new_n967), .A3(new_n970), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n380), .B1(new_n1000), .B2(new_n997), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n343), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n383), .A2(new_n384), .A3(new_n343), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n843), .A2(new_n996), .A3(new_n1003), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n1002), .A2(new_n884), .A3(new_n1004), .ZN(G57));
endmodule


