//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0 0 1 1 0 1 1 1 0 1 1 1 1 1 0 1 0 0 0 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 0 0 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n995,
    new_n996;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G226gat), .ZN(new_n206));
  INV_X1    g005(.A(G233gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT25), .ZN(new_n209));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(KEYINPUT24), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G183gat), .B(G190gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT24), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G169gat), .ZN(new_n216));
  INV_X1    g015(.A(G176gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n218), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT66), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n224), .B(new_n218), .C1(new_n220), .C2(new_n221), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n215), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n216), .A2(new_n217), .A3(KEYINPUT23), .ZN(new_n227));
  NAND2_X1  g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT67), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n227), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n232), .B(KEYINPUT68), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n209), .B1(new_n226), .B2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n227), .A2(new_n209), .A3(new_n228), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n215), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n223), .A2(new_n225), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n228), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n239), .B1(KEYINPUT26), .B2(new_n218), .ZN(new_n240));
  OR2_X1    g039(.A1(new_n218), .A2(KEYINPUT26), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT27), .B(G183gat), .ZN(new_n243));
  INV_X1    g042(.A(G190gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n243), .A2(KEYINPUT28), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT28), .B1(new_n243), .B2(new_n244), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n242), .B(new_n210), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n238), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n208), .B1(new_n234), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n215), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n237), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n232), .B(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT25), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n247), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(new_n245), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n240), .A2(new_n241), .B1(G183gat), .B2(G190gat), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n257), .A2(new_n258), .B1(new_n236), .B2(new_n237), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT29), .B1(new_n255), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n250), .B1(new_n260), .B2(new_n208), .ZN(new_n261));
  XNOR2_X1  g060(.A(G197gat), .B(G204gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT72), .B(G218gat), .ZN(new_n263));
  INV_X1    g062(.A(G211gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n262), .B1(new_n265), .B2(KEYINPUT22), .ZN(new_n266));
  XNOR2_X1  g065(.A(G211gat), .B(G218gat), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n262), .B(new_n267), .C1(new_n265), .C2(KEYINPUT22), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n261), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n250), .B(new_n271), .C1(new_n260), .C2(new_n208), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n205), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n272), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n277), .A2(new_n274), .A3(new_n204), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n276), .A2(KEYINPUT30), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT30), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n277), .A2(new_n280), .A3(new_n274), .A4(new_n204), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G155gat), .ZN(new_n283));
  INV_X1    g082(.A(G162gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G155gat), .A2(G162gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XOR2_X1   g086(.A(G141gat), .B(G148gat), .Z(new_n288));
  INV_X1    g087(.A(KEYINPUT2), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT73), .ZN(new_n292));
  INV_X1    g091(.A(G141gat), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n292), .B1(new_n293), .B2(G148gat), .ZN(new_n294));
  INV_X1    g093(.A(G148gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n295), .A2(KEYINPUT73), .A3(G141gat), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n294), .B(new_n296), .C1(G141gat), .C2(new_n295), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n286), .B1(new_n285), .B2(KEYINPUT2), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(KEYINPUT74), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT74), .B1(new_n297), .B2(new_n298), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n291), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  XOR2_X1   g101(.A(G127gat), .B(G134gat), .Z(new_n303));
  XNOR2_X1  g102(.A(G113gat), .B(G120gat), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n303), .B1(KEYINPUT1), .B2(new_n304), .ZN(new_n305));
  XOR2_X1   g104(.A(G113gat), .B(G120gat), .Z(new_n306));
  INV_X1    g105(.A(KEYINPUT1), .ZN(new_n307));
  XNOR2_X1  g106(.A(G127gat), .B(G134gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT4), .B1(new_n302), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n297), .A2(new_n298), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT74), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n290), .B1(new_n314), .B2(new_n299), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT4), .ZN(new_n316));
  INV_X1    g115(.A(new_n310), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n311), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n302), .A2(KEYINPUT3), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT3), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n315), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n310), .B(KEYINPUT75), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n320), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G225gat), .A2(G233gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n319), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n315), .A2(new_n317), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT75), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n310), .B(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n327), .B1(new_n329), .B2(new_n315), .ZN(new_n330));
  INV_X1    g129(.A(new_n325), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n326), .A2(KEYINPUT5), .A3(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G57gat), .B(G85gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n334), .B(KEYINPUT77), .ZN(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G1gat), .B(G29gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n337), .B(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n311), .A2(KEYINPUT78), .A3(new_n318), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT78), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n327), .A2(new_n342), .A3(KEYINPUT4), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n331), .A2(KEYINPUT5), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n341), .A2(new_n343), .A3(new_n324), .A4(new_n344), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n333), .A2(KEYINPUT79), .A3(new_n340), .A4(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT6), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n345), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n339), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n340), .B1(new_n333), .B2(new_n345), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT79), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n333), .A2(new_n340), .A3(new_n345), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n282), .B(new_n351), .C1(KEYINPUT6), .C2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G228gat), .A2(G233gat), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT29), .B1(new_n269), .B2(new_n270), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n302), .B1(new_n358), .B2(KEYINPUT3), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT80), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n357), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT29), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n362), .B1(new_n302), .B2(KEYINPUT3), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(new_n272), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n359), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n364), .B(new_n359), .C1(new_n360), .C2(new_n357), .ZN(new_n367));
  AOI21_X1  g166(.A(G22gat), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n366), .A2(G22gat), .A3(new_n367), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  XOR2_X1   g170(.A(G78gat), .B(G106gat), .Z(new_n372));
  XNOR2_X1  g171(.A(KEYINPUT31), .B(G50gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n372), .B(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n374), .B1(new_n368), .B2(KEYINPUT81), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n369), .A2(KEYINPUT81), .A3(new_n370), .A4(new_n374), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n356), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT70), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n234), .A2(new_n249), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n380), .B1(new_n381), .B2(new_n317), .ZN(new_n382));
  OAI211_X1 g181(.A(KEYINPUT70), .B(new_n310), .C1(new_n234), .C2(new_n249), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(KEYINPUT69), .A3(new_n317), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n255), .A2(new_n259), .A3(new_n317), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT69), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n382), .A2(new_n383), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT34), .ZN(new_n389));
  NAND2_X1  g188(.A1(G227gat), .A2(G233gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(KEYINPUT64), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n388), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n382), .A2(new_n383), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n384), .A2(new_n387), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n394), .A2(new_n390), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n396), .A2(KEYINPUT71), .A3(KEYINPUT34), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT71), .B1(new_n396), .B2(KEYINPUT34), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n393), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(KEYINPUT32), .B1(new_n388), .B2(new_n392), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT33), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n402), .B1(new_n388), .B2(new_n392), .ZN(new_n403));
  XOR2_X1   g202(.A(G15gat), .B(G43gat), .Z(new_n404));
  XNOR2_X1  g203(.A(G71gat), .B(G99gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n404), .B(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n401), .A2(new_n403), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n406), .ZN(new_n408));
  OAI221_X1 g207(.A(KEYINPUT32), .B1(new_n402), .B2(new_n408), .C1(new_n388), .C2(new_n392), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n400), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT34), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT71), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n397), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n415), .A2(new_n407), .A3(new_n409), .A4(new_n393), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n411), .A2(new_n416), .A3(KEYINPUT36), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT36), .B1(new_n411), .B2(new_n416), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n379), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n351), .B1(new_n355), .B2(KEYINPUT6), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT37), .B1(new_n273), .B2(new_n275), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT37), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n277), .A2(new_n422), .A3(new_n274), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n423), .A3(new_n205), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT38), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT83), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n424), .A2(KEYINPUT83), .A3(KEYINPUT38), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT38), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n421), .A2(new_n429), .A3(new_n423), .A4(new_n205), .ZN(new_n430));
  AND2_X1   g229(.A1(new_n430), .A2(new_n278), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n420), .A2(new_n427), .A3(new_n428), .A4(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n341), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n324), .A2(new_n343), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n331), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n435), .B(KEYINPUT39), .C1(new_n331), .C2(new_n330), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT39), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n437), .B(new_n331), .C1(new_n433), .C2(new_n434), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT82), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n438), .A2(new_n439), .A3(new_n340), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n439), .B1(new_n438), .B2(new_n340), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n436), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT40), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n282), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n436), .B(KEYINPUT40), .C1(new_n440), .C2(new_n441), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n444), .A2(new_n445), .A3(new_n350), .A4(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n378), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n432), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n419), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT84), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n400), .A2(new_n410), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n415), .A2(new_n393), .B1(new_n407), .B2(new_n409), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT35), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n376), .A2(new_n455), .A3(new_n377), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n356), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT85), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n411), .A2(new_n416), .A3(KEYINPUT84), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n454), .A2(new_n457), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n454), .A2(new_n457), .A3(new_n459), .ZN(new_n461));
  INV_X1    g260(.A(new_n356), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n462), .A2(new_n448), .A3(new_n416), .A4(new_n411), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n461), .A2(KEYINPUT85), .B1(new_n463), .B2(KEYINPUT35), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n450), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(G229gat), .A2(G233gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(G29gat), .A2(G36gat), .ZN(new_n467));
  INV_X1    g266(.A(G50gat), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT15), .B1(new_n468), .B2(G43gat), .ZN(new_n469));
  INV_X1    g268(.A(G43gat), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n470), .A2(G50gat), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n467), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT15), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT87), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(new_n468), .B2(G43gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n468), .A2(G43gat), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n470), .A2(KEYINPUT87), .A3(G50gat), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n472), .B1(new_n473), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT88), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT86), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT14), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT14), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT86), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(G29gat), .A2(G36gat), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n482), .A2(new_n486), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n480), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n486), .B1(new_n482), .B2(new_n484), .ZN(new_n491));
  AOI211_X1 g290(.A(G29gat), .B(G36gat), .C1(new_n481), .C2(KEYINPUT14), .ZN(new_n492));
  NOR3_X1   g291(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT88), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n479), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n467), .B1(new_n491), .B2(new_n492), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n469), .A2(new_n471), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(G15gat), .B(G22gat), .ZN(new_n499));
  INV_X1    g298(.A(G1gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT16), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n499), .A2(G1gat), .ZN(new_n504));
  OAI21_X1  g303(.A(G8gat), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(G8gat), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n502), .B(new_n506), .C1(G1gat), .C2(new_n499), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n498), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n494), .A2(KEYINPUT17), .A3(new_n497), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n505), .A2(new_n507), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT88), .B1(new_n491), .B2(new_n492), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT86), .B(KEYINPUT14), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n480), .B(new_n489), .C1(new_n514), .C2(new_n486), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g315(.A1(new_n516), .A2(new_n479), .B1(new_n495), .B2(new_n496), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n517), .A2(KEYINPUT17), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n466), .B(new_n509), .C1(new_n512), .C2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT89), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT18), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n520), .B1(new_n519), .B2(new_n521), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n466), .B(KEYINPUT13), .Z(new_n525));
  NOR2_X1   g324(.A1(new_n498), .A2(new_n508), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n511), .A2(new_n517), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(new_n519), .B2(new_n521), .ZN(new_n529));
  XNOR2_X1  g328(.A(G113gat), .B(G141gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(G197gat), .ZN(new_n531));
  XOR2_X1   g330(.A(KEYINPUT11), .B(G169gat), .Z(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n533), .B(KEYINPUT12), .Z(new_n534));
  NOR2_X1   g333(.A1(new_n529), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n508), .B1(new_n517), .B2(KEYINPUT17), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT17), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n498), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n527), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n539), .A2(KEYINPUT18), .A3(new_n466), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n519), .A2(new_n521), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(new_n541), .A3(new_n528), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n524), .A2(new_n535), .B1(new_n542), .B2(new_n534), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n465), .A2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G57gat), .B(G64gat), .Z(new_n545));
  OR2_X1    g344(.A1(G71gat), .A2(G78gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(G71gat), .A2(G78gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT9), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n545), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G57gat), .B(G64gat), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n547), .B(new_n546), .C1(new_n552), .C2(new_n549), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT21), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(G231gat), .A2(G233gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(G127gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n554), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n508), .B1(KEYINPUT21), .B2(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n560), .B(new_n562), .Z(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(new_n283), .ZN(new_n565));
  XNOR2_X1  g364(.A(G183gat), .B(G211gat), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n565), .B(new_n566), .Z(new_n567));
  NAND2_X1  g366(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n560), .B(new_n562), .ZN(new_n569));
  INV_X1    g368(.A(new_n567), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G99gat), .B(G106gat), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT7), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT90), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT90), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT7), .ZN(new_n578));
  AND2_X1   g377(.A1(G85gat), .A2(G92gat), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n576), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G99gat), .A2(G106gat), .ZN(new_n581));
  INV_X1    g380(.A(G85gat), .ZN(new_n582));
  INV_X1    g381(.A(G92gat), .ZN(new_n583));
  AOI22_X1  g382(.A1(KEYINPUT8), .A2(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n579), .B1(new_n576), .B2(new_n578), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n574), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n576), .A2(new_n578), .ZN(new_n588));
  INV_X1    g387(.A(new_n579), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n590), .A2(new_n573), .A3(new_n580), .A4(new_n584), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  AND2_X1   g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593));
  AOI22_X1  g392(.A1(new_n498), .A2(new_n592), .B1(KEYINPUT41), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n587), .A2(new_n591), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n510), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n594), .B1(new_n596), .B2(new_n518), .ZN(new_n597));
  XOR2_X1   g396(.A(G190gat), .B(G218gat), .Z(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n593), .A2(KEYINPUT41), .ZN(new_n600));
  XNOR2_X1  g399(.A(G134gat), .B(G162gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n598), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n594), .B(new_n603), .C1(new_n596), .C2(new_n518), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n599), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n602), .B1(new_n599), .B2(new_n604), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT92), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n551), .A2(new_n553), .A3(KEYINPUT10), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n592), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT92), .B1(new_n595), .B2(new_n610), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT91), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n591), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n595), .A2(new_n561), .A3(new_n616), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n591), .B(new_n587), .C1(new_n554), .C2(new_n615), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT10), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(G230gat), .ZN(new_n620));
  OAI22_X1  g419(.A1(new_n614), .A2(new_n619), .B1(new_n620), .B2(new_n207), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n207), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n617), .A2(new_n622), .A3(new_n618), .ZN(new_n623));
  XNOR2_X1  g422(.A(G120gat), .B(G148gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(G176gat), .B(G204gat), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n624), .B(new_n625), .Z(new_n626));
  NAND3_X1  g425(.A1(new_n621), .A2(new_n623), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n626), .B1(new_n621), .B2(new_n623), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n572), .A2(new_n608), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n544), .A2(new_n420), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(KEYINPUT93), .B(G1gat), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(G1324gat));
  XOR2_X1   g434(.A(KEYINPUT16), .B(G8gat), .Z(new_n636));
  NAND4_X1  g435(.A1(new_n544), .A2(new_n445), .A3(new_n632), .A4(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT94), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT42), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n638), .B1(new_n637), .B2(new_n639), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n461), .A2(KEYINPUT85), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n463), .A2(KEYINPUT35), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n643), .A2(new_n460), .A3(new_n644), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n419), .A2(new_n449), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT18), .B1(new_n539), .B2(new_n466), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n534), .B1(new_n529), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n541), .A2(KEYINPUT89), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n534), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n540), .A2(new_n653), .A3(new_n528), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n649), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n647), .A2(new_n655), .A3(new_n445), .A4(new_n632), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(G8gat), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(KEYINPUT95), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT95), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n656), .A2(new_n659), .A3(G8gat), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n661), .B1(new_n639), .B2(new_n637), .ZN(new_n662));
  OAI21_X1  g461(.A(KEYINPUT96), .B1(new_n642), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n637), .A2(new_n639), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n664), .B1(new_n658), .B2(new_n660), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT96), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n665), .B(new_n666), .C1(new_n641), .C2(new_n640), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n663), .A2(new_n667), .ZN(G1325gat));
  NAND2_X1  g467(.A1(new_n544), .A2(new_n632), .ZN(new_n669));
  OR2_X1    g468(.A1(new_n417), .A2(new_n418), .ZN(new_n670));
  OAI21_X1  g469(.A(G15gat), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n454), .ZN(new_n672));
  INV_X1    g471(.A(new_n459), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n675), .A2(G15gat), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n671), .B1(new_n669), .B2(new_n676), .ZN(G1326gat));
  OR3_X1    g476(.A1(new_n669), .A2(KEYINPUT97), .A3(new_n448), .ZN(new_n678));
  OAI21_X1  g477(.A(KEYINPUT97), .B1(new_n669), .B2(new_n448), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT43), .B(G22gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1327gat));
  XOR2_X1   g481(.A(new_n572), .B(KEYINPUT98), .Z(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n630), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n684), .A2(new_n543), .A3(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(KEYINPUT99), .A2(KEYINPUT44), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n687), .B1(new_n647), .B2(new_n607), .ZN(new_n688));
  XOR2_X1   g487(.A(KEYINPUT99), .B(KEYINPUT44), .Z(new_n689));
  AOI211_X1 g488(.A(new_n608), .B(new_n689), .C1(new_n645), .C2(new_n646), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n420), .B(new_n686), .C1(new_n688), .C2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT100), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI22_X1  g492(.A1(new_n465), .A2(new_n608), .B1(KEYINPUT99), .B2(KEYINPUT44), .ZN(new_n694));
  INV_X1    g493(.A(new_n689), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n647), .A2(new_n607), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n697), .A2(KEYINPUT100), .A3(new_n420), .A4(new_n686), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n693), .A2(G29gat), .A3(new_n698), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n572), .A2(new_n608), .A3(new_n685), .ZN(new_n700));
  INV_X1    g499(.A(new_n420), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(G29gat), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n544), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT45), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT101), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n699), .A2(new_n704), .A3(KEYINPUT101), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(G1328gat));
  NAND2_X1  g508(.A1(new_n544), .A2(new_n700), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n710), .A2(G36gat), .A3(new_n282), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT46), .ZN(new_n712));
  INV_X1    g511(.A(G36gat), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n697), .A2(new_n686), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n714), .A2(new_n445), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n712), .B1(new_n713), .B2(new_n715), .ZN(G1329gat));
  NAND4_X1  g515(.A1(new_n544), .A2(new_n470), .A3(new_n674), .A4(new_n700), .ZN(new_n717));
  INV_X1    g516(.A(new_n670), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  OAI211_X1 g518(.A(KEYINPUT47), .B(new_n717), .C1(new_n719), .C2(new_n470), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT47), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n470), .B1(new_n714), .B2(new_n718), .ZN(new_n722));
  INV_X1    g521(.A(new_n717), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n720), .A2(new_n724), .ZN(G1330gat));
  INV_X1    g524(.A(KEYINPUT48), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n697), .A2(new_n378), .A3(new_n686), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(new_n468), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n378), .A2(new_n468), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n710), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n726), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  OAI221_X1 g530(.A(KEYINPUT48), .B1(new_n710), .B2(new_n729), .C1(new_n727), .C2(new_n468), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(G1331gat));
  NAND3_X1  g532(.A1(new_n572), .A2(new_n608), .A3(new_n685), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n465), .A2(new_n655), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n420), .ZN(new_n736));
  XOR2_X1   g535(.A(KEYINPUT102), .B(G57gat), .Z(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1332gat));
  INV_X1    g537(.A(KEYINPUT49), .ZN(new_n739));
  INV_X1    g538(.A(G64gat), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n445), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT103), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n735), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n739), .A2(new_n740), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1333gat));
  INV_X1    g544(.A(G71gat), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n735), .A2(new_n746), .A3(new_n674), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n735), .A2(new_n718), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n748), .B2(new_n746), .ZN(new_n749));
  XNOR2_X1  g548(.A(KEYINPUT104), .B(KEYINPUT50), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(G1334gat));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n378), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g552(.A1(new_n572), .A2(new_n655), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n685), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n755), .B(KEYINPUT105), .Z(new_n756));
  AND2_X1   g555(.A1(new_n697), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n420), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(G85gat), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n465), .A2(new_n608), .ZN(new_n760));
  AOI22_X1  g559(.A1(new_n760), .A2(new_n754), .B1(KEYINPUT106), .B2(KEYINPUT51), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT107), .ZN(new_n763));
  XOR2_X1   g562(.A(KEYINPUT106), .B(KEYINPUT51), .Z(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n760), .A2(new_n754), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n762), .A2(new_n763), .A3(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n763), .B1(new_n762), .B2(new_n766), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n685), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n420), .A2(new_n582), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n759), .B1(new_n770), .B2(new_n771), .ZN(G1336gat));
  INV_X1    g571(.A(new_n766), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n773), .A2(new_n761), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n282), .A2(new_n630), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n583), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n697), .A2(new_n445), .A3(new_n756), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(new_n583), .ZN(new_n779));
  OAI21_X1  g578(.A(KEYINPUT52), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781));
  OAI221_X1 g580(.A(new_n781), .B1(new_n778), .B2(new_n583), .C1(new_n774), .C2(new_n776), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(G1337gat));
  NAND2_X1  g582(.A1(new_n757), .A2(new_n718), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G99gat), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n675), .A2(G99gat), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n770), .B2(new_n786), .ZN(G1338gat));
  NOR3_X1   g586(.A1(new_n448), .A2(G106gat), .A3(new_n630), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n788), .B1(new_n773), .B2(new_n761), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n697), .A2(new_n378), .A3(new_n756), .ZN(new_n790));
  INV_X1    g589(.A(G106gat), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT53), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n789), .B(new_n794), .C1(new_n790), .C2(new_n791), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(G1339gat));
  NAND2_X1  g595(.A1(new_n617), .A2(new_n618), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT10), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n612), .A2(new_n613), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n799), .A2(new_n622), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT108), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n799), .A2(KEYINPUT108), .A3(new_n622), .A4(new_n800), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n803), .A2(KEYINPUT54), .A3(new_n621), .A4(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n622), .B1(new_n799), .B2(new_n800), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n626), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n805), .A2(KEYINPUT55), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n627), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT55), .B1(new_n805), .B2(new_n808), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n810), .A2(new_n543), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n524), .A2(new_n535), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n539), .A2(new_n466), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n526), .A2(new_n527), .A3(new_n525), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n533), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n817), .A2(new_n630), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n608), .B1(new_n812), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT109), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n813), .A2(new_n607), .A3(new_n816), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n821), .A2(new_n810), .A3(new_n811), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n819), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n805), .A2(new_n808), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n827), .A2(new_n655), .A3(new_n627), .A4(new_n809), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n685), .A2(new_n813), .A3(new_n816), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n607), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT109), .B1(new_n830), .B2(new_n822), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n824), .A2(new_n683), .A3(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n631), .A2(new_n655), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n832), .A2(KEYINPUT110), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT110), .B1(new_n832), .B2(new_n834), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n835), .A2(new_n836), .A3(new_n701), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n448), .A2(new_n416), .A3(new_n411), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n837), .A2(new_n282), .A3(new_n839), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(KEYINPUT112), .ZN(new_n841));
  INV_X1    g640(.A(G113gat), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(new_n842), .A3(new_n655), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n701), .A2(new_n445), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n674), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n835), .A2(new_n836), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(KEYINPUT111), .A3(new_n448), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n834), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT110), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n832), .A2(KEYINPUT110), .A3(new_n834), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(new_n448), .A3(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT111), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n845), .B1(new_n847), .B2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(G113gat), .B1(new_n856), .B2(new_n543), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n843), .A2(new_n857), .ZN(G1340gat));
  NOR2_X1   g657(.A1(new_n630), .A2(G120gat), .ZN(new_n859));
  XOR2_X1   g658(.A(new_n859), .B(KEYINPUT113), .Z(new_n860));
  NAND2_X1  g659(.A1(new_n841), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(G120gat), .B1(new_n856), .B2(new_n630), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(G1341gat));
  NAND3_X1  g662(.A1(new_n855), .A2(G127gat), .A3(new_n684), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n837), .A2(new_n282), .A3(new_n839), .A4(new_n572), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT114), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n559), .B1(new_n865), .B2(new_n866), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n864), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT115), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n864), .B(new_n871), .C1(new_n867), .C2(new_n868), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(G1342gat));
  OAI21_X1  g672(.A(G134gat), .B1(new_n856), .B2(new_n608), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n837), .A2(new_n839), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n445), .A2(new_n608), .ZN(new_n876));
  INV_X1    g675(.A(G134gat), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT56), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  OR3_X1    g678(.A1(new_n875), .A2(KEYINPUT56), .A3(new_n878), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n874), .A2(new_n879), .A3(new_n880), .ZN(G1343gat));
  NAND2_X1  g680(.A1(new_n819), .A2(new_n823), .ZN(new_n882));
  INV_X1    g681(.A(new_n572), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n833), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n884), .A2(new_n885), .A3(new_n448), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n850), .A2(new_n378), .A3(new_n851), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(new_n885), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n670), .A2(new_n844), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n888), .A2(new_n543), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT118), .B1(new_n890), .B2(new_n293), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n670), .A2(new_n378), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n892), .B1(new_n837), .B2(KEYINPUT116), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n850), .A2(new_n420), .A3(new_n851), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT116), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n655), .A2(new_n293), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT117), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n893), .A2(new_n282), .A3(new_n896), .A4(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n899), .B1(new_n890), .B2(new_n293), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT58), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n891), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  OAI221_X1 g701(.A(new_n899), .B1(KEYINPUT118), .B2(KEYINPUT58), .C1(new_n890), .C2(new_n293), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n902), .A2(new_n903), .ZN(G1344gat));
  NOR3_X1   g703(.A1(new_n888), .A2(new_n630), .A3(new_n889), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n905), .A2(KEYINPUT59), .A3(new_n295), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n850), .A2(KEYINPUT57), .A3(new_n378), .A4(new_n851), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n882), .A2(KEYINPUT119), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n572), .B1(new_n882), .B2(KEYINPUT119), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n833), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n885), .B1(new_n911), .B2(new_n448), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n913), .A2(new_n670), .A3(new_n685), .A4(new_n844), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n907), .B1(new_n914), .B2(G148gat), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n893), .A2(new_n282), .A3(new_n896), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n685), .A2(new_n295), .ZN(new_n917));
  OAI22_X1  g716(.A1(new_n906), .A2(new_n915), .B1(new_n916), .B2(new_n917), .ZN(G1345gat));
  INV_X1    g717(.A(KEYINPUT120), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n888), .A2(new_n683), .A3(new_n889), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n920), .A2(new_n283), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n572), .A2(new_n283), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n916), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n919), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  OAI221_X1 g723(.A(KEYINPUT120), .B1(new_n916), .B2(new_n922), .C1(new_n283), .C2(new_n920), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1346gat));
  NAND4_X1  g725(.A1(new_n893), .A2(new_n284), .A3(new_n876), .A4(new_n896), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n888), .A2(new_n608), .A3(new_n889), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n928), .B2(new_n284), .ZN(G1347gat));
  NOR3_X1   g728(.A1(new_n835), .A2(new_n836), .A3(new_n420), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(new_n445), .A3(new_n839), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT121), .ZN(new_n932));
  AOI21_X1  g731(.A(G169gat), .B1(new_n932), .B2(new_n655), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n420), .A2(new_n282), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT122), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n674), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n936), .B1(new_n847), .B2(new_n854), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n543), .A2(new_n216), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n933), .B1(new_n937), .B2(new_n938), .ZN(G1348gat));
  NAND3_X1  g738(.A1(new_n932), .A2(new_n217), .A3(new_n685), .ZN(new_n940));
  INV_X1    g739(.A(new_n936), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT111), .B1(new_n846), .B2(new_n448), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n852), .A2(new_n853), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(G176gat), .B1(new_n944), .B2(new_n630), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n940), .A2(new_n945), .ZN(G1349gat));
  OAI21_X1  g745(.A(G183gat), .B1(new_n944), .B2(new_n683), .ZN(new_n947));
  INV_X1    g746(.A(new_n243), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n931), .A2(new_n948), .A3(new_n883), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n947), .A2(new_n950), .A3(new_n951), .A4(KEYINPUT60), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n951), .A2(KEYINPUT60), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(KEYINPUT60), .ZN(new_n954));
  INV_X1    g753(.A(G183gat), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n955), .B1(new_n937), .B2(new_n684), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n953), .B(new_n954), .C1(new_n956), .C2(new_n949), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n952), .A2(new_n957), .ZN(G1350gat));
  NAND3_X1  g757(.A1(new_n932), .A2(new_n244), .A3(new_n607), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n937), .A2(new_n607), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n960), .B1(new_n961), .B2(G190gat), .ZN(new_n962));
  AOI211_X1 g761(.A(KEYINPUT61), .B(new_n244), .C1(new_n937), .C2(new_n607), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(G1351gat));
  NAND3_X1  g763(.A1(new_n930), .A2(new_n378), .A3(new_n670), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n965), .A2(new_n282), .ZN(new_n966));
  XNOR2_X1  g765(.A(KEYINPUT124), .B(G197gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n966), .A2(new_n655), .A3(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(new_n967), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n935), .A2(new_n670), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n908), .A2(KEYINPUT125), .A3(new_n912), .ZN(new_n971));
  INV_X1    g770(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g771(.A(KEYINPUT125), .B1(new_n908), .B2(new_n912), .ZN(new_n973));
  OAI211_X1 g772(.A(new_n655), .B(new_n970), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT126), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n969), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(new_n970), .ZN(new_n977));
  INV_X1    g776(.A(new_n973), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n977), .B1(new_n978), .B2(new_n971), .ZN(new_n979));
  AOI21_X1  g778(.A(KEYINPUT126), .B1(new_n979), .B2(new_n655), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n968), .B1(new_n976), .B2(new_n980), .ZN(G1352gat));
  NAND2_X1  g780(.A1(new_n979), .A2(new_n685), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(G204gat), .ZN(new_n983));
  AOI21_X1  g782(.A(G204gat), .B1(KEYINPUT127), .B2(KEYINPUT62), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n775), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n965), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g785(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n987));
  XOR2_X1   g786(.A(new_n986), .B(new_n987), .Z(new_n988));
  NAND2_X1  g787(.A1(new_n983), .A2(new_n988), .ZN(G1353gat));
  NAND3_X1  g788(.A1(new_n913), .A2(new_n572), .A3(new_n970), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(G211gat), .ZN(new_n991));
  XOR2_X1   g790(.A(new_n991), .B(KEYINPUT63), .Z(new_n992));
  NAND3_X1  g791(.A1(new_n966), .A2(new_n264), .A3(new_n572), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n992), .A2(new_n993), .ZN(G1354gat));
  AOI21_X1  g793(.A(G218gat), .B1(new_n966), .B2(new_n607), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n608), .A2(new_n263), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n995), .B1(new_n979), .B2(new_n996), .ZN(G1355gat));
endmodule


