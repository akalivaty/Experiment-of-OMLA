//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0 0 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1265, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1322, new_n1323,
    new_n1324;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n208), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n202), .A2(G50), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n210), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n213), .B1(new_n216), .B2(new_n217), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT2), .B(G226), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G264), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XOR2_X1   g0035(.A(G107), .B(G116), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  NAND3_X1  g0041(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(new_n214), .ZN(new_n243));
  INV_X1    g0043(.A(KEYINPUT67), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NOR2_X1   g0045(.A1(G20), .A2(G33), .ZN(new_n246));
  INV_X1    g0046(.A(G68), .ZN(new_n247));
  AOI22_X1  g0047(.A1(new_n246), .A2(G50), .B1(G20), .B2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G77), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n208), .A2(G33), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AND2_X1   g0051(.A1(new_n245), .A2(new_n251), .ZN(new_n252));
  OR2_X1    g0052(.A1(new_n252), .A2(KEYINPUT11), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n207), .A2(G13), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(new_n208), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(new_n243), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n207), .A2(G20), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(G68), .A3(new_n257), .ZN(new_n258));
  XOR2_X1   g0058(.A(new_n258), .B(KEYINPUT74), .Z(new_n259));
  NAND2_X1  g0059(.A1(new_n252), .A2(KEYINPUT11), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n255), .A2(new_n247), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n261), .B(KEYINPUT12), .ZN(new_n262));
  AND4_X1   g0062(.A1(new_n253), .A2(new_n259), .A3(new_n260), .A4(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G232), .A3(G1698), .ZN(new_n269));
  INV_X1    g0069(.A(G1698), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n268), .A2(G226), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G97), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n214), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT13), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT64), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(KEYINPUT64), .A2(G33), .A3(G41), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(new_n274), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G41), .ZN(new_n284));
  INV_X1    g0084(.A(G45), .ZN(new_n285));
  AOI21_X1  g0085(.A(G1), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n283), .A2(G274), .A3(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n286), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n283), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G238), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n278), .A2(new_n279), .A3(new_n287), .A4(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(G1698), .B1(new_n266), .B2(new_n267), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n293), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n276), .B1(new_n294), .B2(new_n269), .ZN(new_n295));
  INV_X1    g0095(.A(G238), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n287), .B1(new_n289), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT13), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT14), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(new_n300), .A3(G169), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n292), .A2(new_n298), .A3(G179), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n300), .B1(new_n299), .B2(G169), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT75), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n304), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT75), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n306), .A2(new_n307), .A3(new_n302), .A4(new_n301), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n263), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT8), .B(G58), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT68), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n310), .B(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n312), .B1(new_n207), .B2(G20), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n245), .A2(new_n255), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n313), .A2(new_n314), .B1(new_n312), .B2(new_n255), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT16), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT7), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(new_n268), .B2(G20), .ZN(new_n318));
  AND2_X1   g0118(.A1(KEYINPUT3), .A2(G33), .ZN(new_n319));
  NOR2_X1   g0119(.A1(KEYINPUT3), .A2(G33), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n321), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n247), .B1(new_n318), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G58), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n324), .A2(new_n247), .ZN(new_n325));
  OAI21_X1  g0125(.A(G20), .B1(new_n325), .B2(new_n201), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n246), .A2(G159), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n316), .B1(new_n323), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT7), .B1(new_n321), .B2(new_n208), .ZN(new_n330));
  NOR4_X1   g0130(.A1(new_n319), .A2(new_n320), .A3(new_n317), .A4(G20), .ZN(new_n331));
  OAI21_X1  g0131(.A(G68), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n328), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(KEYINPUT16), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n329), .A2(new_n243), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n315), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT76), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT76), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n315), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n270), .B1(new_n266), .B2(new_n267), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n340), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n293), .A2(G223), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n276), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G232), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n287), .B1(new_n289), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(G169), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n341), .A2(new_n342), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n277), .ZN(new_n348));
  INV_X1    g0148(.A(new_n345), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G179), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n346), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n337), .A2(new_n339), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT18), .ZN(new_n354));
  INV_X1    g0154(.A(G190), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n355), .A2(KEYINPUT77), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n355), .A2(KEYINPUT77), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n348), .A2(new_n349), .A3(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(G200), .B1(new_n343), .B2(new_n345), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n315), .A2(new_n335), .A3(new_n360), .A4(new_n361), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n362), .B(KEYINPUT17), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT18), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n337), .A2(new_n364), .A3(new_n339), .A4(new_n352), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n354), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n263), .B1(new_n355), .B2(new_n299), .ZN(new_n367));
  INV_X1    g0167(.A(G200), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(new_n292), .B2(new_n298), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  OR3_X1    g0170(.A1(new_n309), .A2(new_n366), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT73), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n293), .A2(G222), .B1(new_n321), .B2(G77), .ZN(new_n373));
  INV_X1    g0173(.A(new_n340), .ZN(new_n374));
  XNOR2_X1  g0174(.A(KEYINPUT65), .B(G223), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OR2_X1    g0176(.A1(new_n376), .A2(KEYINPUT66), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(KEYINPUT66), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n378), .A3(new_n277), .ZN(new_n379));
  INV_X1    g0179(.A(new_n287), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n380), .B1(G226), .B2(new_n290), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G169), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G150), .ZN(new_n385));
  INV_X1    g0185(.A(new_n246), .ZN(new_n386));
  OAI22_X1  g0186(.A1(new_n312), .A2(new_n250), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n387), .A2(KEYINPUT69), .ZN(new_n388));
  OAI21_X1  g0188(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n387), .B2(KEYINPUT69), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n245), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(G50), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n392), .B1(new_n207), .B2(G20), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n314), .A2(new_n393), .B1(new_n392), .B2(new_n255), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n379), .A2(new_n351), .A3(new_n381), .ZN(new_n396));
  AND3_X1   g0196(.A1(new_n384), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  XNOR2_X1  g0198(.A(new_n395), .B(KEYINPUT9), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n368), .B1(new_n379), .B2(new_n381), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT10), .B1(new_n400), .B2(KEYINPUT72), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n382), .A2(new_n355), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n402), .A2(new_n400), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n399), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n401), .B1(new_n399), .B2(new_n403), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n398), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n268), .A2(G232), .A3(new_n270), .ZN(new_n408));
  INV_X1    g0208(.A(G107), .ZN(new_n409));
  OAI221_X1 g0209(.A(new_n408), .B1(new_n409), .B2(new_n268), .C1(new_n374), .C2(new_n296), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n277), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n290), .A2(G244), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n287), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n383), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n255), .A2(new_n249), .ZN(new_n415));
  INV_X1    g0215(.A(new_n256), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n257), .A2(G77), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n310), .B1(KEYINPUT70), .B2(new_n386), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(KEYINPUT70), .B2(new_n386), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G20), .A2(G77), .ZN(new_n421));
  XNOR2_X1  g0221(.A(KEYINPUT15), .B(G87), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT71), .ZN(new_n423));
  XNOR2_X1  g0223(.A(new_n422), .B(new_n423), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n420), .B(new_n421), .C1(new_n424), .C2(new_n250), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n418), .B1(new_n425), .B2(new_n243), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n414), .B(new_n427), .C1(G179), .C2(new_n413), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n413), .A2(G200), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(new_n426), .C1(new_n355), .C2(new_n413), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n372), .B1(new_n407), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n399), .A2(new_n403), .ZN(new_n433));
  INV_X1    g0233(.A(new_n401), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n404), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n428), .A2(new_n430), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n436), .A2(KEYINPUT73), .A3(new_n398), .A4(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n371), .B1(new_n432), .B2(new_n438), .ZN(new_n439));
  OAI211_X1 g0239(.A(G244), .B(new_n270), .C1(new_n319), .C2(new_n320), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT4), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT78), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n440), .A2(KEYINPUT78), .A3(new_n441), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n293), .A2(KEYINPUT4), .A3(G244), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n340), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n444), .A2(new_n445), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n277), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n285), .A2(G1), .ZN(new_n450));
  XNOR2_X1  g0250(.A(KEYINPUT5), .B(G41), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n283), .A2(G274), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  AND2_X1   g0252(.A1(KEYINPUT5), .A2(G41), .ZN(new_n453));
  NOR2_X1   g0253(.A1(KEYINPUT5), .A2(G41), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n450), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n283), .A2(new_n455), .A3(G257), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT79), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n452), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n457), .B1(new_n452), .B2(new_n456), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n449), .A2(new_n460), .A3(G190), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT81), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT81), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n449), .A2(new_n460), .A3(new_n463), .A4(G190), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NOR3_X1   g0265(.A1(new_n458), .A2(new_n459), .A3(KEYINPUT80), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT80), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n452), .A2(new_n456), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT79), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n452), .A2(new_n456), .A3(new_n457), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n467), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n449), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G200), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n207), .A2(G33), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n314), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G97), .ZN(new_n476));
  OAI21_X1  g0276(.A(G107), .B1(new_n330), .B2(new_n331), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT6), .ZN(new_n478));
  AND2_X1   g0278(.A1(G97), .A2(G107), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n478), .B1(new_n479), .B2(new_n204), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n409), .A2(KEYINPUT6), .A3(G97), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n482), .A2(G20), .B1(G77), .B2(new_n246), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(G97), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n484), .A2(new_n243), .B1(new_n485), .B2(new_n255), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n476), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n465), .A2(new_n473), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT82), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n487), .B1(new_n462), .B2(new_n464), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(KEYINPUT82), .A3(new_n473), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n449), .A2(new_n460), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n383), .A2(new_n495), .B1(new_n476), .B2(new_n486), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n351), .B(new_n449), .C1(new_n466), .C2(new_n471), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AND3_X1   g0298(.A1(KEYINPUT64), .A2(G33), .A3(G41), .ZN(new_n499));
  AOI21_X1  g0299(.A(KEYINPUT64), .B1(G33), .B2(G41), .ZN(new_n500));
  NOR3_X1   g0300(.A1(new_n499), .A2(new_n500), .A3(new_n214), .ZN(new_n501));
  INV_X1    g0301(.A(G250), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(new_n285), .B2(G1), .ZN(new_n503));
  INV_X1    g0303(.A(G274), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n207), .A2(new_n504), .A3(G45), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(KEYINPUT83), .B1(new_n501), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT83), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n283), .A2(new_n508), .A3(new_n503), .A4(new_n505), .ZN(new_n509));
  OAI211_X1 g0309(.A(G238), .B(new_n270), .C1(new_n319), .C2(new_n320), .ZN(new_n510));
  OAI211_X1 g0310(.A(G244), .B(G1698), .C1(new_n319), .C2(new_n320), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G116), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n507), .A2(new_n509), .B1(new_n513), .B2(new_n277), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n514), .A2(G190), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n514), .A2(new_n368), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT19), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n208), .B1(new_n272), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(G87), .B2(new_n205), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n518), .B1(new_n250), .B2(new_n485), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n268), .A2(new_n208), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n520), .B(new_n521), .C1(new_n522), .C2(new_n247), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n243), .ZN(new_n524));
  XNOR2_X1  g0324(.A(new_n243), .B(KEYINPUT67), .ZN(new_n525));
  INV_X1    g0325(.A(new_n254), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G20), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n525), .A2(G87), .A3(new_n527), .A4(new_n474), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n424), .A2(new_n255), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n524), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n507), .A2(new_n509), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n513), .A2(new_n277), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n532), .A2(new_n533), .A3(G179), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n383), .B2(new_n514), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n314), .A2(new_n474), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n524), .B(new_n529), .C1(new_n536), .C2(new_n424), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n517), .A2(new_n531), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n494), .A2(new_n498), .A3(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n512), .A2(G20), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT23), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n208), .B2(G107), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n409), .A2(KEYINPUT23), .A3(G20), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT22), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n321), .A2(G20), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n545), .B1(new_n546), .B2(G87), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n268), .A2(new_n545), .A3(new_n208), .A4(G87), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n544), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT86), .ZN(new_n551));
  XOR2_X1   g0351(.A(KEYINPUT85), .B(KEYINPUT24), .Z(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n552), .ZN(new_n554));
  INV_X1    g0354(.A(new_n544), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n268), .A2(new_n208), .A3(G87), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(KEYINPUT22), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n555), .B1(new_n557), .B2(new_n548), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n554), .B1(new_n558), .B2(KEYINPUT86), .ZN(new_n559));
  AOI211_X1 g0359(.A(new_n551), .B(new_n555), .C1(new_n557), .C2(new_n548), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n553), .B(new_n243), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n255), .A2(KEYINPUT25), .A3(new_n409), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT87), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT25), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n527), .B2(G107), .ZN(new_n565));
  XNOR2_X1  g0365(.A(new_n563), .B(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n314), .A2(G107), .A3(new_n474), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n561), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n283), .A2(new_n455), .A3(G264), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT88), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT88), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n283), .A2(new_n455), .A3(new_n573), .A4(G264), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n268), .A2(G257), .A3(G1698), .ZN(new_n576));
  NAND2_X1  g0376(.A1(G33), .A2(G294), .ZN(new_n577));
  OAI211_X1 g0377(.A(G250), .B(new_n270), .C1(new_n319), .C2(new_n320), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n277), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n575), .A2(new_n452), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT89), .B1(new_n581), .B2(G169), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(KEYINPUT89), .A3(G169), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n351), .B2(new_n581), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n570), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n572), .A2(new_n574), .B1(new_n579), .B2(new_n277), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n586), .A2(KEYINPUT90), .A3(new_n355), .A4(new_n452), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT90), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(new_n581), .B2(new_n368), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n581), .A2(G190), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n587), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n550), .A2(new_n551), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n558), .A2(KEYINPUT86), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n592), .A2(new_n593), .A3(new_n554), .ZN(new_n594));
  INV_X1    g0394(.A(new_n243), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n557), .A2(new_n548), .ZN(new_n596));
  AOI21_X1  g0396(.A(KEYINPUT86), .B1(new_n596), .B2(new_n544), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n595), .B1(new_n597), .B2(new_n552), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n568), .B1(new_n594), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n591), .A2(new_n599), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n585), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(G116), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n242), .A2(new_n214), .B1(G20), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(G33), .A2(G283), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n604), .B(new_n208), .C1(G33), .C2(new_n485), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT20), .ZN(new_n607));
  OAI21_X1  g0407(.A(KEYINPUT84), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT84), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n603), .A2(new_n610), .A3(new_n605), .A4(KEYINPUT20), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n602), .A2(G20), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n254), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n602), .B1(new_n207), .B2(G33), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n614), .B1(new_n256), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n268), .A2(G264), .A3(G1698), .ZN(new_n618));
  OAI211_X1 g0418(.A(G257), .B(new_n270), .C1(new_n319), .C2(new_n320), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n321), .A2(G303), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n277), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n283), .A2(new_n455), .A3(G270), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n622), .A2(new_n452), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n617), .A2(new_n624), .A3(G169), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT21), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n624), .A2(new_n351), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n617), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n621), .A2(new_n277), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n452), .A2(new_n623), .ZN(new_n631));
  OAI21_X1  g0431(.A(G200), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n612), .A2(new_n616), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n622), .A2(new_n359), .A3(new_n452), .A4(new_n623), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n617), .A2(new_n624), .A3(KEYINPUT21), .A4(G169), .ZN(new_n636));
  AND4_X1   g0436(.A1(new_n627), .A2(new_n629), .A3(new_n635), .A4(new_n636), .ZN(new_n637));
  AND4_X1   g0437(.A1(new_n439), .A2(new_n539), .A3(new_n601), .A4(new_n637), .ZN(G372));
  NAND2_X1  g0438(.A1(new_n305), .A2(new_n308), .ZN(new_n639));
  INV_X1    g0439(.A(new_n263), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n428), .B2(new_n370), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n642), .A2(new_n363), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n336), .A2(new_n352), .A3(KEYINPUT95), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT95), .B1(new_n336), .B2(new_n352), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n364), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n336), .A2(new_n352), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT95), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n336), .A2(new_n352), .A3(KEYINPUT95), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(KEYINPUT18), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n436), .B1(new_n643), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n398), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n439), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT91), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n532), .A2(new_n533), .A3(G179), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n383), .B1(new_n532), .B2(new_n533), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n534), .B(KEYINPUT91), .C1(new_n383), .C2(new_n514), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n537), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n663), .A2(KEYINPUT93), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(KEYINPUT93), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n538), .A2(KEYINPUT26), .A3(new_n497), .A4(new_n496), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n667), .A2(KEYINPUT94), .ZN(new_n668));
  INV_X1    g0468(.A(new_n498), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n515), .A2(new_n516), .A3(new_n530), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n670), .B1(new_n662), .B2(new_n537), .ZN(new_n671));
  AOI21_X1  g0471(.A(KEYINPUT26), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n667), .A2(KEYINPUT94), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n666), .B(new_n668), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n671), .A2(new_n600), .A3(new_n498), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n492), .A2(KEYINPUT82), .A3(new_n473), .ZN(new_n676));
  AOI21_X1  g0476(.A(KEYINPUT82), .B1(new_n492), .B2(new_n473), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n627), .A2(new_n629), .A3(new_n636), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n678), .A2(KEYINPUT92), .B1(new_n585), .B2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT92), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n675), .B(new_n681), .C1(new_n676), .C2(new_n677), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n674), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n655), .B1(new_n656), .B2(new_n683), .ZN(G369));
  OR3_X1    g0484(.A1(new_n254), .A2(KEYINPUT27), .A3(G20), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT27), .B1(new_n254), .B2(G20), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G213), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G343), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n601), .B1(new_n599), .B2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n585), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n689), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n617), .A2(new_n689), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n637), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n679), .B2(new_n695), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n694), .A2(G330), .A3(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n679), .A2(new_n689), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n601), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n692), .A2(new_n690), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n698), .A2(new_n703), .ZN(G399));
  INV_X1    g0504(.A(new_n211), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G41), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(G1), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n217), .B2(new_n707), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n585), .A2(new_n679), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT98), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT98), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n585), .A2(new_n714), .A3(new_n679), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n494), .A2(new_n713), .A3(new_n675), .A4(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT26), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n538), .A2(new_n717), .A3(new_n497), .A4(new_n496), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n664), .A2(new_n665), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n717), .B1(new_n669), .B2(new_n671), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n689), .B1(new_n716), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT29), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(KEYINPUT97), .B1(new_n683), .B2(new_n689), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n672), .A2(new_n673), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n664), .B(new_n665), .C1(KEYINPUT94), .C2(new_n667), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n671), .A2(new_n600), .A3(new_n498), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n491), .B2(new_n493), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n712), .B1(new_n730), .B2(new_n681), .ZN(new_n731));
  INV_X1    g0531(.A(new_n682), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n728), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT97), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(new_n734), .A3(new_n690), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n725), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT29), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n724), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G330), .ZN(new_n739));
  AND4_X1   g0539(.A1(new_n585), .A2(new_n637), .A3(new_n600), .A4(new_n690), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n494), .A2(new_n740), .A3(new_n498), .A4(new_n538), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n514), .A2(G179), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n472), .A2(new_n581), .A3(new_n624), .A4(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT96), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(KEYINPUT30), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n586), .A2(new_n514), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n628), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n745), .B1(new_n747), .B2(new_n495), .ZN(new_n748));
  INV_X1    g0548(.A(new_n495), .ZN(new_n749));
  INV_X1    g0549(.A(new_n745), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n749), .A2(new_n628), .A3(new_n750), .A4(new_n746), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n743), .A2(new_n748), .A3(new_n751), .ZN(new_n752));
  AND3_X1   g0552(.A1(new_n752), .A2(KEYINPUT31), .A3(new_n689), .ZN(new_n753));
  AOI21_X1  g0553(.A(KEYINPUT31), .B1(new_n752), .B2(new_n689), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n739), .B1(new_n741), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n738), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n711), .B1(new_n757), .B2(G1), .ZN(G364));
  INV_X1    g0558(.A(G13), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n207), .B1(new_n760), .B2(G45), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n706), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(new_n697), .B2(G330), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n764), .B1(G330), .B2(new_n697), .ZN(new_n765));
  INV_X1    g0565(.A(new_n763), .ZN(new_n766));
  OAI21_X1  g0566(.A(G20), .B1(KEYINPUT100), .B2(G169), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(KEYINPUT100), .A2(G169), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n214), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n208), .A2(new_n351), .A3(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n355), .ZN(new_n773));
  INV_X1    g0573(.A(G311), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n355), .A2(G179), .A3(G200), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n208), .ZN(new_n776));
  INV_X1    g0576(.A(G294), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n773), .A2(new_n774), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n358), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G326), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n779), .A2(G190), .ZN(new_n784));
  XNOR2_X1  g0584(.A(KEYINPUT33), .B(G317), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n778), .B(new_n783), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n208), .A2(G190), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n787), .A2(new_n351), .A3(new_n368), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n268), .B1(new_n789), .B2(G329), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n359), .A2(new_n772), .ZN(new_n791));
  INV_X1    g0591(.A(G322), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OR3_X1    g0593(.A1(new_n368), .A2(KEYINPUT101), .A3(G179), .ZN(new_n794));
  OAI21_X1  g0594(.A(KEYINPUT101), .B1(new_n368), .B2(G179), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n208), .A2(new_n355), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n793), .B1(G303), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G283), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n794), .A2(new_n787), .A3(new_n795), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n786), .B(new_n799), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n791), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n803), .A2(G58), .B1(G50), .B2(new_n780), .ZN(new_n804));
  INV_X1    g0604(.A(G159), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n788), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT32), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n806), .A2(new_n807), .B1(new_n773), .B2(new_n249), .ZN(new_n808));
  INV_X1    g0608(.A(new_n784), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n776), .A2(new_n485), .B1(new_n809), .B2(new_n247), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n321), .B1(new_n806), .B2(new_n807), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n801), .A2(new_n409), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(G87), .B2(new_n798), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n804), .A2(new_n811), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n771), .B1(new_n802), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(G13), .A2(G33), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(G20), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n770), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n211), .A2(new_n268), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n821), .B(KEYINPUT99), .Z(new_n822));
  INV_X1    g0622(.A(G355), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n822), .A2(new_n823), .B1(G116), .B2(new_n211), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n705), .A2(new_n268), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(G45), .B2(new_n217), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(G45), .B2(new_n240), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n766), .B(new_n816), .C1(new_n820), .C2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n819), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n829), .B1(new_n697), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n765), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G396));
  INV_X1    g0633(.A(KEYINPUT102), .ZN(new_n834));
  OR3_X1    g0634(.A1(new_n428), .A2(new_n834), .A3(new_n690), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n834), .B1(new_n428), .B2(new_n690), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n427), .A2(new_n689), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n835), .A2(new_n836), .B1(new_n437), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(new_n725), .B2(new_n735), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n690), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n678), .A2(KEYINPUT92), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n842), .A2(new_n682), .A3(new_n712), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n841), .B1(new_n843), .B2(new_n728), .ZN(new_n844));
  OR3_X1    g0644(.A1(new_n840), .A2(new_n756), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n756), .B1(new_n840), .B2(new_n844), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n845), .A2(new_n766), .A3(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT103), .ZN(new_n848));
  INV_X1    g0648(.A(new_n773), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n780), .A2(G137), .B1(new_n849), .B2(G159), .ZN(new_n850));
  INV_X1    g0650(.A(G143), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n850), .B1(new_n851), .B2(new_n791), .C1(new_n385), .C2(new_n809), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT34), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n852), .A2(new_n853), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n801), .A2(new_n247), .ZN(new_n856));
  INV_X1    g0656(.A(G132), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n268), .B1(new_n788), .B2(new_n857), .C1(new_n776), .C2(new_n324), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n856), .B(new_n858), .C1(G50), .C2(new_n798), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n854), .A2(new_n855), .A3(new_n859), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n321), .B1(new_n788), .B2(new_n774), .C1(new_n776), .C2(new_n485), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(G107), .B2(new_n798), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n803), .A2(G294), .B1(G283), .B2(new_n784), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n780), .A2(G303), .B1(new_n849), .B2(G116), .ZN(new_n864));
  INV_X1    g0664(.A(new_n801), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(G87), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n862), .A2(new_n863), .A3(new_n864), .A4(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n771), .B1(new_n860), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n770), .A2(new_n817), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n868), .B1(new_n249), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n839), .B2(new_n818), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n763), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n847), .A2(new_n848), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n848), .B1(new_n847), .B2(new_n872), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(G384));
  NOR2_X1   g0675(.A1(new_n760), .A2(new_n207), .ZN(new_n876));
  INV_X1    g0676(.A(new_n370), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n263), .A2(new_n690), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n641), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n878), .B1(new_n309), .B2(new_n370), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n838), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n741), .A2(new_n755), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT106), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n882), .A2(KEYINPUT106), .A3(new_n883), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT40), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n649), .A2(new_n362), .A3(new_n650), .ZN(new_n889));
  INV_X1    g0689(.A(new_n687), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n337), .A2(new_n339), .A3(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT37), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT37), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n362), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n353), .A2(new_n891), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n646), .A2(new_n651), .A3(new_n363), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n892), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT38), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n329), .A2(new_n245), .A3(new_n334), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n315), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n890), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n366), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n903), .A2(new_n352), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n907), .A2(new_n904), .A3(new_n362), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT37), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n896), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n906), .A2(KEYINPUT38), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n888), .B1(new_n901), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n886), .A2(new_n887), .A3(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n906), .A2(new_n910), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT38), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n911), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n914), .B1(new_n884), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n913), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n439), .A2(new_n883), .ZN(new_n922));
  OR2_X1    g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n922), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n923), .A2(G330), .A3(new_n924), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n925), .B(KEYINPUT107), .Z(new_n926));
  AOI21_X1  g0726(.A(new_n654), .B1(new_n738), .B2(new_n439), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n428), .A2(new_n689), .ZN(new_n928));
  INV_X1    g0728(.A(new_n841), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n928), .B1(new_n733), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n879), .B1(new_n641), .B2(new_n877), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n309), .A2(new_n370), .A3(new_n878), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n930), .A2(new_n933), .A3(new_n919), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT39), .ZN(new_n935));
  AOI221_X4 g0735(.A(new_n916), .B1(new_n896), .B2(new_n909), .C1(new_n366), .C2(new_n905), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n935), .B1(new_n900), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n917), .A2(KEYINPUT39), .A3(new_n911), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n641), .A2(new_n689), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n652), .A2(new_n687), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n934), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n927), .B(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n876), .B1(new_n926), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n926), .B2(new_n944), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n602), .B(new_n216), .C1(new_n482), .C2(KEYINPUT35), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(KEYINPUT35), .B2(new_n482), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT36), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n217), .A2(new_n249), .A3(new_n325), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT104), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n950), .A2(new_n951), .B1(new_n392), .B2(G68), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n951), .B2(new_n950), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(G1), .A3(new_n759), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n946), .A2(new_n949), .A3(new_n954), .ZN(G367));
  INV_X1    g0755(.A(new_n825), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n820), .B1(new_n211), .B2(new_n424), .C1(new_n956), .C2(new_n233), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT110), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n776), .A2(new_n247), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n791), .A2(new_n385), .B1(new_n805), .B2(new_n809), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n959), .B(new_n960), .C1(G50), .C2(new_n849), .ZN(new_n961));
  INV_X1    g0761(.A(G137), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n268), .B1(new_n788), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n801), .A2(new_n249), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n963), .B(new_n964), .C1(G143), .C2(new_n780), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n961), .B(new_n965), .C1(new_n324), .C2(new_n797), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n801), .A2(new_n485), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n268), .B(new_n967), .C1(G317), .C2(new_n789), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n969), .A2(KEYINPUT112), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n773), .A2(new_n800), .B1(new_n776), .B2(new_n409), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n803), .A2(G303), .B1(G311), .B2(new_n780), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n777), .B2(new_n809), .ZN(new_n973));
  NOR3_X1   g0773(.A1(new_n970), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(KEYINPUT112), .B2(new_n969), .ZN(new_n975));
  AOI21_X1  g0775(.A(KEYINPUT111), .B1(new_n798), .B2(G116), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT46), .Z(new_n977));
  OAI21_X1  g0777(.A(new_n966), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT47), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n766), .B(new_n958), .C1(new_n979), .C2(new_n770), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT113), .Z(new_n981));
  NOR2_X1   g0781(.A1(new_n531), .A2(new_n690), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n982), .B(new_n670), .C1(new_n662), .C2(new_n537), .ZN(new_n983));
  INV_X1    g0783(.A(new_n666), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n983), .B1(new_n984), .B2(new_n982), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n981), .B1(new_n819), .B2(new_n985), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n498), .B1(new_n488), .B2(new_n690), .C1(new_n676), .C2(new_n677), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n498), .A2(new_n690), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT108), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT109), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n692), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n689), .B1(new_n992), .B2(new_n498), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT43), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n700), .B1(new_n987), .B2(new_n989), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT42), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n994), .A2(new_n995), .A3(new_n985), .A4(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n698), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n991), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n985), .A2(new_n995), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n985), .A2(new_n995), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n997), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1001), .B(new_n1002), .C1(new_n993), .C2(new_n1003), .ZN(new_n1004));
  AND3_X1   g0804(.A1(new_n998), .A2(new_n1000), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1000), .B1(new_n998), .B2(new_n1004), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n990), .A2(new_n703), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT45), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n990), .A2(KEYINPUT45), .A3(new_n703), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n987), .A2(new_n702), .A3(new_n989), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT44), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1013), .B(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n999), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1012), .A2(new_n1015), .A3(new_n698), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n700), .B1(new_n694), .B2(new_n699), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n697), .A2(G330), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1020), .B(new_n1021), .Z(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n757), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n706), .B(KEYINPUT41), .Z(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n761), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n986), .B1(new_n1007), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(G387));
  OAI21_X1  g0830(.A(new_n1023), .B1(new_n738), .B2(new_n756), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n756), .ZN(new_n1032));
  AOI21_X1  g0832(.A(KEYINPUT29), .B1(new_n725), .B2(new_n735), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1022), .B(new_n1032), .C1(new_n1033), .C2(new_n724), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n706), .B(KEYINPUT117), .Z(new_n1035));
  NAND3_X1  g0835(.A1(new_n1031), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n691), .A2(new_n693), .A3(new_n819), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n825), .B1(new_n230), .B2(new_n285), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n708), .B2(new_n822), .ZN(new_n1039));
  OR3_X1    g0839(.A1(new_n310), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1040));
  OAI21_X1  g0840(.A(KEYINPUT50), .B1(new_n310), .B2(G50), .ZN(new_n1041));
  AOI21_X1  g0841(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1040), .A2(new_n708), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n1039), .A2(new_n1043), .B1(new_n409), .B2(new_n705), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n820), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n763), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n321), .B1(new_n789), .B2(G150), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n247), .B2(new_n773), .C1(new_n791), .C2(new_n392), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n967), .B1(G77), .B2(new_n798), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n424), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n776), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1049), .B(new_n1052), .C1(new_n312), .C2(new_n809), .ZN(new_n1053));
  OAI21_X1  g0853(.A(KEYINPUT114), .B1(new_n781), .B2(new_n805), .ZN(new_n1054));
  OR3_X1    g0854(.A1(new_n781), .A2(KEYINPUT114), .A3(new_n805), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1048), .B(new_n1053), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT115), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n268), .B1(new_n789), .B2(G326), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n780), .A2(G322), .B1(G311), .B2(new_n784), .ZN(new_n1059));
  INV_X1    g0859(.A(G303), .ZN(new_n1060));
  INV_X1    g0860(.A(G317), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1059), .B1(new_n1060), .B2(new_n773), .C1(new_n1061), .C2(new_n791), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT116), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1064), .A2(KEYINPUT48), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(KEYINPUT48), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n798), .A2(G294), .B1(new_n1051), .B2(G283), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT49), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1058), .B1(new_n602), .B2(new_n801), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1068), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1071), .A2(KEYINPUT49), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1057), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1046), .B1(new_n1073), .B2(new_n770), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n1022), .A2(new_n762), .B1(new_n1037), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1036), .A2(new_n1075), .ZN(G393));
  NAND3_X1  g0876(.A1(new_n1017), .A2(new_n762), .A3(new_n1018), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n825), .A2(new_n237), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n820), .B1(new_n485), .B2(new_n211), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n763), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n781), .A2(new_n1061), .B1(new_n791), .B2(new_n774), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT52), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n268), .B(new_n813), .C1(G322), .C2(new_n789), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1082), .B(new_n1083), .C1(new_n800), .C2(new_n797), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G294), .A2(new_n849), .B1(new_n1051), .B2(G116), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n1060), .B2(new_n809), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT118), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n866), .B1(new_n247), .B2(new_n797), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n268), .B1(new_n788), .B2(new_n851), .C1(new_n776), .C2(new_n249), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n773), .A2(new_n310), .B1(new_n809), .B2(new_n392), .ZN(new_n1090));
  OR3_X1    g0890(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n803), .A2(G159), .B1(G150), .B2(new_n780), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT51), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n1084), .A2(new_n1087), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1080), .B1(new_n1094), .B2(new_n770), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n991), .B2(new_n830), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1077), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT119), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1077), .A2(KEYINPUT119), .A3(new_n1096), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OR2_X1    g0901(.A1(new_n1034), .A2(new_n1019), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1034), .A2(new_n1019), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1102), .A2(new_n1103), .A3(new_n1035), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1101), .A2(new_n1104), .ZN(G390));
  NAND2_X1  g0905(.A1(new_n882), .A2(new_n756), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1107), .A2(KEYINPUT120), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n937), .A2(new_n938), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n933), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n844), .B2(new_n928), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n939), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1109), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n722), .A2(new_n839), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n928), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n933), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1112), .B1(new_n900), .B2(new_n936), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT120), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n1116), .A2(new_n1117), .B1(new_n1118), .B2(new_n1106), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1108), .B1(new_n1113), .B2(new_n1119), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n689), .B(new_n838), .C1(new_n716), .C2(new_n721), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1110), .B1(new_n1121), .B2(new_n928), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1117), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1122), .A2(new_n1123), .B1(new_n1107), .B2(KEYINPUT120), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1108), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1115), .B1(new_n683), .B2(new_n841), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n939), .B1(new_n1126), .B2(new_n1110), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1124), .B(new_n1125), .C1(new_n1127), .C2(new_n1109), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1120), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n762), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n766), .B1(new_n312), .B2(new_n869), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n321), .B1(new_n789), .B2(G125), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n962), .B2(new_n809), .ZN(new_n1133));
  XOR2_X1   g0933(.A(KEYINPUT54), .B(G143), .Z(new_n1134));
  AOI22_X1  g0934(.A1(new_n780), .A2(G128), .B1(new_n849), .B2(new_n1134), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1135), .B1(new_n857), .B2(new_n791), .C1(new_n805), .C2(new_n776), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1133), .B(new_n1136), .C1(G50), .C2(new_n865), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n797), .A2(new_n385), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT53), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n781), .A2(new_n800), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n791), .A2(new_n602), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n773), .A2(new_n485), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n809), .A2(new_n409), .ZN(new_n1143));
  NOR4_X1   g0943(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n321), .B1(new_n788), .B2(new_n777), .C1(new_n776), .C2(new_n249), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n856), .B(new_n1145), .C1(G87), .C2(new_n798), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1137), .A2(new_n1139), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1131), .B1(new_n771), .B2(new_n1147), .C1(new_n1109), .C2(new_n818), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1130), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1035), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT122), .ZN(new_n1151));
  AOI211_X1 g0951(.A(KEYINPUT97), .B(new_n689), .C1(new_n843), .C2(new_n728), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n734), .B1(new_n733), .B2(new_n690), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n737), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1154), .A2(new_n439), .A3(new_n723), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n439), .A2(new_n756), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1155), .A2(new_n655), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n756), .A2(new_n839), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n1160), .A2(new_n933), .B1(new_n756), .B2(new_n882), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT121), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1159), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n739), .B(new_n838), .C1(new_n741), .C2(new_n755), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1106), .B1(new_n1164), .B2(new_n1110), .ZN(new_n1165));
  OAI21_X1  g0965(.A(KEYINPUT121), .B1(new_n1165), .B2(new_n1158), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1161), .A2(new_n930), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1163), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1151), .B1(new_n1157), .B2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1150), .B1(new_n1169), .B2(new_n1129), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n1165), .A2(KEYINPUT121), .A3(new_n1158), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1167), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1162), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1171), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n927), .A2(new_n1174), .A3(new_n1156), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1175), .A2(new_n1151), .A3(new_n1120), .A4(new_n1128), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1149), .B1(new_n1170), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(G378));
  INV_X1    g0978(.A(new_n869), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n763), .B1(new_n1179), .B2(G50), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n395), .A2(new_n890), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n436), .B2(new_n398), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1183), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n397), .B(new_n1185), .C1(new_n435), .C2(new_n404), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1182), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n407), .A2(new_n1185), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n436), .A2(new_n398), .A3(new_n1183), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1188), .A2(new_n1189), .A3(new_n1181), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1187), .A2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1191), .A2(new_n818), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n268), .A2(G41), .ZN(new_n1193));
  AOI211_X1 g0993(.A(G50), .B(new_n1193), .C1(new_n265), .C2(new_n284), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n781), .A2(new_n602), .B1(new_n485), .B2(new_n809), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(G107), .B2(new_n803), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1193), .B1(new_n800), .B2(new_n788), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n959), .B(new_n1197), .C1(G77), .C2(new_n798), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1050), .A2(new_n849), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n865), .A2(G58), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1196), .A2(new_n1198), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT58), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1194), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  AOI211_X1 g1003(.A(G33), .B(G41), .C1(new_n789), .C2(G124), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n780), .A2(G125), .B1(new_n1051), .B2(G150), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT123), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n803), .A2(G128), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n857), .B2(new_n809), .C1(new_n962), .C2(new_n773), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1206), .B(new_n1208), .C1(new_n798), .C2(new_n1134), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT59), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1204), .B1(new_n805), .B2(new_n801), .C1(new_n1209), .C2(new_n1210), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1203), .B1(new_n1202), .B2(new_n1201), .C1(new_n1211), .C2(new_n1212), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1180), .B(new_n1192), .C1(new_n770), .C2(new_n1213), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n913), .A2(G330), .A3(new_n920), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1191), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n934), .B2(new_n942), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1126), .A2(new_n1110), .A3(new_n918), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1218), .A2(new_n1191), .A3(new_n940), .A4(new_n941), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1215), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1217), .A2(new_n1215), .A3(new_n1219), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1214), .B1(new_n1223), .B2(new_n762), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1129), .A2(new_n1174), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1157), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(KEYINPUT57), .B1(new_n1227), .B2(new_n1223), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1217), .A2(new_n1219), .A3(new_n1215), .ZN(new_n1229));
  OAI21_X1  g1029(.A(KEYINPUT57), .B1(new_n1229), .B2(new_n1220), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1157), .B1(new_n1129), .B2(new_n1174), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1035), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1224), .B1(new_n1228), .B2(new_n1232), .ZN(G375));
  XOR2_X1   g1033(.A(new_n761), .B(KEYINPUT125), .Z(new_n1234));
  OR2_X1    g1034(.A1(new_n1168), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n933), .A2(new_n817), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n763), .B1(new_n1179), .B2(G68), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n803), .A2(G137), .B1(new_n784), .B2(new_n1134), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1239), .B1(new_n392), .B2(new_n776), .C1(new_n857), .C2(new_n781), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n798), .A2(G159), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n849), .A2(G150), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n321), .B1(new_n789), .B2(G128), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1200), .A2(new_n1241), .A3(new_n1242), .A4(new_n1243), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n321), .B1(new_n788), .B2(new_n1060), .C1(new_n773), .C2(new_n409), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1245), .A2(new_n964), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1246), .B(new_n1052), .C1(new_n485), .C2(new_n797), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n780), .A2(G294), .B1(G116), .B2(new_n784), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n800), .B2(new_n791), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n1240), .A2(new_n1244), .B1(new_n1247), .B2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1238), .B1(new_n1250), .B2(new_n770), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1236), .B1(new_n1237), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1157), .A2(new_n1168), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(KEYINPUT124), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT124), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1157), .A2(new_n1255), .A3(new_n1168), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1254), .A2(new_n1026), .A3(new_n1175), .A4(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1252), .A2(new_n1257), .ZN(G381));
  INV_X1    g1058(.A(G384), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1036), .A2(new_n832), .A3(new_n1075), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1029), .A2(new_n1259), .A3(new_n1260), .A4(new_n1262), .ZN(new_n1263));
  OR4_X1    g1063(.A1(G378), .A2(new_n1263), .A3(G375), .A4(G381), .ZN(G407));
  NAND2_X1  g1064(.A1(new_n1177), .A2(new_n688), .ZN(new_n1265));
  OAI211_X1 g1065(.A(G407), .B(G213), .C1(G375), .C2(new_n1265), .ZN(G409));
  AOI21_X1  g1066(.A(new_n832), .B1(new_n1036), .B2(new_n1075), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1260), .B1(new_n1262), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1267), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1269), .A2(G390), .A3(new_n1261), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1268), .A2(new_n1029), .A3(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1029), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1272));
  OR2_X1    g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(KEYINPUT60), .B1(new_n1157), .B2(new_n1168), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1254), .A2(new_n1256), .A3(new_n1274), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1157), .A2(new_n1168), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1150), .B1(new_n1276), .B2(KEYINPUT60), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1278), .A2(G384), .A3(new_n1252), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G384), .B1(new_n1278), .B2(new_n1252), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1229), .A2(new_n1220), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1168), .B1(new_n1120), .B2(new_n1128), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1026), .B1(new_n1283), .B2(new_n1157), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1282), .B1(new_n1284), .B2(new_n1234), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1177), .B1(new_n1214), .B2(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1286), .B1(G375), .B2(new_n1177), .ZN(new_n1287));
  INV_X1    g1087(.A(G213), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1288), .A2(G343), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1281), .A2(new_n1287), .A3(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(KEYINPUT62), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT62), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1281), .A2(new_n1287), .A3(new_n1293), .A4(new_n1290), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT61), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1289), .A2(G2897), .ZN(new_n1297));
  XOR2_X1   g1097(.A(new_n1297), .B(KEYINPUT127), .Z(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1299), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1278), .A2(new_n1252), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1259), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1278), .A2(G384), .A3(new_n1252), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1302), .A2(new_n1303), .A3(new_n1298), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1300), .A2(new_n1304), .ZN(new_n1305));
  OAI211_X1 g1105(.A(G378), .B(new_n1224), .C1(new_n1228), .C2(new_n1232), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1289), .B1(new_n1306), .B2(new_n1286), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1296), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1273), .B1(new_n1295), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1287), .A2(new_n1290), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(KEYINPUT126), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT126), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1287), .A2(new_n1312), .A3(new_n1290), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1311), .A2(new_n1313), .A3(new_n1304), .A4(new_n1300), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1281), .A2(new_n1287), .A3(KEYINPUT63), .A4(new_n1290), .ZN(new_n1315));
  NOR3_X1   g1115(.A1(new_n1271), .A2(new_n1272), .A3(KEYINPUT61), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT63), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1291), .A2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1314), .A2(new_n1317), .A3(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1309), .A2(new_n1320), .ZN(G405));
  NAND2_X1  g1121(.A1(G375), .A2(new_n1177), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1306), .A2(new_n1322), .ZN(new_n1323));
  XNOR2_X1  g1123(.A(new_n1323), .B(new_n1281), .ZN(new_n1324));
  XNOR2_X1  g1124(.A(new_n1324), .B(new_n1273), .ZN(G402));
endmodule


