//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(G217), .ZN(new_n189));
  NOR3_X1   g003(.A1(new_n188), .A2(new_n189), .A3(G953), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  INV_X1    g005(.A(G122), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT14), .B1(new_n192), .B2(G116), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT86), .B(G122), .ZN(new_n194));
  INV_X1    g008(.A(G116), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n193), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT14), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n192), .A2(G116), .ZN(new_n198));
  AOI22_X1  g012(.A1(new_n196), .A2(KEYINPUT87), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT87), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n200), .B(new_n193), .C1(new_n194), .C2(new_n195), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n191), .B1(new_n199), .B2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n192), .A2(KEYINPUT86), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT86), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G122), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n195), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  NOR3_X1   g020(.A1(new_n206), .A2(G107), .A3(new_n198), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  AND2_X1   g022(.A1(KEYINPUT65), .A2(G134), .ZN(new_n209));
  NOR2_X1   g023(.A1(KEYINPUT65), .A2(G134), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G128), .ZN(new_n213));
  INV_X1    g027(.A(G128), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G143), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n211), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(new_n215), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n218));
  INV_X1    g032(.A(G134), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT65), .A2(G134), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n216), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n208), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT88), .B1(new_n202), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n193), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT87), .B1(new_n206), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n198), .A2(new_n197), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(new_n201), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G107), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT88), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n231), .A2(new_n232), .A3(new_n208), .A4(new_n224), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n226), .A2(new_n233), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n213), .A2(new_n215), .A3(KEYINPUT13), .ZN(new_n235));
  OAI21_X1  g049(.A(G134), .B1(new_n213), .B2(KEYINPUT13), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n216), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(G107), .B1(new_n206), .B2(new_n198), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n237), .B1(new_n208), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n190), .B1(new_n234), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n190), .ZN(new_n242));
  AOI211_X1 g056(.A(new_n239), .B(new_n242), .C1(new_n226), .C2(new_n233), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n187), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT89), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G478), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(KEYINPUT15), .ZN(new_n248));
  OAI211_X1 g062(.A(KEYINPUT89), .B(new_n187), .C1(new_n241), .C2(new_n243), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n246), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  OR2_X1    g064(.A1(new_n244), .A2(new_n248), .ZN(new_n251));
  INV_X1    g065(.A(G953), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n252), .A2(G952), .ZN(new_n253));
  NAND2_X1  g067(.A1(G234), .A2(G237), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n254), .A2(G902), .A3(G953), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT21), .B(G898), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n256), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n250), .A2(new_n251), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(KEYINPUT18), .A2(G131), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G237), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT67), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT67), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G237), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  AND4_X1   g083(.A1(G143), .A2(new_n269), .A3(G214), .A4(new_n252), .ZN(new_n270));
  AOI21_X1  g084(.A(G953), .B1(new_n266), .B2(new_n268), .ZN(new_n271));
  AOI21_X1  g085(.A(G143), .B1(new_n271), .B2(G214), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n264), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G140), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G125), .ZN(new_n275));
  INV_X1    g089(.A(G125), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G140), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G146), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n278), .B(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n269), .A2(G214), .A3(new_n252), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n212), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n271), .A2(G143), .A3(G214), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n283), .A3(new_n263), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n273), .A2(new_n280), .A3(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(G131), .B1(new_n270), .B2(new_n272), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT17), .ZN(new_n287));
  INV_X1    g101(.A(G131), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n282), .A2(new_n288), .A3(new_n283), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n286), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  OAI211_X1 g104(.A(KEYINPUT17), .B(G131), .C1(new_n270), .C2(new_n272), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n275), .A2(new_n277), .A3(KEYINPUT16), .ZN(new_n292));
  OR3_X1    g106(.A1(new_n276), .A2(KEYINPUT16), .A3(G140), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n292), .A2(new_n293), .A3(KEYINPUT73), .A4(G146), .ZN(new_n294));
  AOI21_X1  g108(.A(G146), .B1(new_n292), .B2(new_n293), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT73), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n292), .A2(new_n293), .A3(G146), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n291), .A2(new_n294), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n285), .B1(new_n290), .B2(new_n299), .ZN(new_n300));
  XOR2_X1   g114(.A(G113), .B(G122), .Z(new_n301));
  XOR2_X1   g115(.A(KEYINPUT83), .B(G104), .Z(new_n302));
  XOR2_X1   g116(.A(new_n301), .B(new_n302), .Z(new_n303));
  NAND2_X1  g117(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n303), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n285), .B(new_n305), .C1(new_n290), .C2(new_n299), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n187), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n308), .A2(G475), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT85), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT84), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n273), .A2(new_n280), .A3(new_n284), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n275), .A2(new_n277), .A3(KEYINPUT19), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT19), .B1(new_n275), .B2(new_n277), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n297), .B1(new_n316), .B2(G146), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n317), .B1(new_n286), .B2(new_n289), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n303), .B1(new_n313), .B2(new_n318), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n306), .A2(new_n312), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n312), .B1(new_n306), .B2(new_n319), .ZN(new_n321));
  NOR2_X1   g135(.A1(G475), .A2(G902), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NOR3_X1   g137(.A1(new_n320), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT20), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n311), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n306), .A2(new_n319), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT84), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n306), .A2(new_n312), .A3(new_n319), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n322), .A3(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(KEYINPUT85), .A3(KEYINPUT20), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n327), .A2(new_n325), .A3(new_n322), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n326), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n262), .A2(new_n310), .A3(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(G214), .B1(G237), .B2(G902), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(G210), .B1(G237), .B2(G902), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT6), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT2), .B(G113), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(G116), .B(G119), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n341), .A2(KEYINPUT5), .ZN(new_n343));
  INV_X1    g157(.A(G119), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G116), .ZN(new_n345));
  OAI21_X1  g159(.A(G113), .B1(new_n345), .B2(KEYINPUT5), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n342), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G104), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT3), .B1(new_n348), .B2(G107), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT3), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(new_n191), .A3(G104), .ZN(new_n351));
  INV_X1    g165(.A(G101), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n348), .A2(G107), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n349), .A2(new_n351), .A3(new_n352), .A4(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n348), .A2(G107), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n191), .A2(G104), .ZN(new_n356));
  OAI21_X1  g170(.A(G101), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n347), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n341), .B(new_n339), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n349), .A2(new_n351), .A3(new_n353), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G101), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n354), .A2(KEYINPUT4), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n360), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT4), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n361), .A2(new_n365), .A3(G101), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT77), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n361), .A2(KEYINPUT77), .A3(new_n365), .A4(G101), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n359), .B1(new_n364), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(G110), .B(G122), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT81), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n372), .B(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n338), .B1(new_n371), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n359), .ZN(new_n376));
  INV_X1    g190(.A(new_n370), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n363), .A2(new_n362), .ZN(new_n378));
  INV_X1    g192(.A(new_n360), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n376), .B1(new_n377), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n372), .B(KEYINPUT81), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n375), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n214), .A2(KEYINPUT1), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n279), .A2(G143), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n212), .A2(G146), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n212), .A2(KEYINPUT1), .A3(G146), .ZN(new_n389));
  XNOR2_X1  g203(.A(G143), .B(G146), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n388), .B(new_n389), .C1(G128), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n276), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT0), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n214), .ZN(new_n394));
  NAND2_X1  g208(.A1(KEYINPUT0), .A2(G128), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n386), .A2(new_n387), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n386), .A2(new_n387), .A3(new_n395), .ZN(new_n397));
  OAI21_X1  g211(.A(G125), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n392), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT82), .ZN(new_n400));
  INV_X1    g214(.A(G224), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n401), .A2(G953), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT82), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n392), .A2(new_n398), .A3(new_n403), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n400), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n402), .B1(new_n400), .B2(new_n404), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n381), .A2(new_n338), .A3(new_n382), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n384), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT7), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n402), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n399), .B(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT8), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n374), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n382), .A2(KEYINPUT8), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n347), .A2(new_n358), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n416), .B1(new_n376), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n371), .A2(new_n374), .ZN(new_n420));
  AOI21_X1  g234(.A(G902), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n337), .B1(new_n409), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n409), .A2(new_n337), .A3(new_n421), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n336), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n426));
  INV_X1    g240(.A(G469), .ZN(new_n427));
  INV_X1    g241(.A(G137), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT11), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT64), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT64), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT11), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n222), .A2(new_n428), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n220), .A2(G137), .A3(new_n221), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n428), .A2(KEYINPUT11), .A3(G134), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(G131), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n430), .A2(new_n432), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n438), .B1(new_n211), .B2(G137), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n428), .A2(KEYINPUT11), .A3(G134), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n440), .B1(new_n211), .B2(G137), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(new_n441), .A3(new_n288), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n388), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n389), .B1(new_n390), .B2(G128), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT78), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI211_X1 g261(.A(KEYINPUT78), .B(new_n389), .C1(new_n390), .C2(G128), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n358), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n354), .A2(new_n357), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n450), .A2(new_n391), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n443), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT12), .ZN(new_n453));
  OR2_X1    g267(.A1(new_n453), .A2(KEYINPUT80), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(KEYINPUT80), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n452), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT79), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n391), .A2(KEYINPUT10), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n457), .B1(new_n458), .B2(new_n358), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n450), .A2(KEYINPUT79), .A3(KEYINPUT10), .A4(new_n391), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(G128), .B1(new_n386), .B2(new_n387), .ZN(new_n462));
  INV_X1    g276(.A(new_n389), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n446), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(new_n388), .A3(new_n448), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n450), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT10), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(KEYINPUT66), .B1(new_n396), .B2(new_n397), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n386), .A2(new_n387), .A3(new_n395), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT66), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n394), .A2(new_n395), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n470), .B(new_n471), .C1(new_n472), .C2(new_n390), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n370), .A2(new_n474), .A3(new_n378), .ZN(new_n475));
  INV_X1    g289(.A(new_n443), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n461), .A2(new_n468), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  OR2_X1    g291(.A1(new_n450), .A2(new_n391), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n466), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n479), .A2(KEYINPUT80), .A3(new_n453), .A4(new_n443), .ZN(new_n480));
  XNOR2_X1  g294(.A(G110), .B(G140), .ZN(new_n481));
  INV_X1    g295(.A(G227), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(G953), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n481), .B(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n456), .A2(new_n477), .A3(new_n480), .A4(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n461), .A2(new_n475), .A3(new_n468), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n443), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n485), .B1(new_n489), .B2(new_n477), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n427), .B(new_n187), .C1(new_n487), .C2(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n427), .A2(new_n187), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n456), .A2(new_n477), .A3(new_n480), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n484), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n489), .A2(new_n485), .A3(new_n477), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(G469), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n491), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n425), .A2(new_n426), .A3(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n334), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT30), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n396), .A2(new_n397), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n502), .B1(new_n437), .B2(new_n442), .ZN(new_n503));
  NOR3_X1   g317(.A1(new_n433), .A2(new_n436), .A3(G131), .ZN(new_n504));
  AOI21_X1  g318(.A(G137), .B1(new_n220), .B2(new_n221), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n428), .A2(G134), .ZN(new_n506));
  OAI21_X1  g320(.A(G131), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n391), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n501), .B1(new_n503), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n288), .B1(new_n439), .B2(new_n441), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n474), .B1(new_n504), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n442), .A2(new_n507), .A3(new_n391), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(KEYINPUT30), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n510), .A2(new_n514), .A3(new_n379), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n512), .A2(new_n360), .A3(new_n513), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n271), .A2(G210), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT27), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT26), .B(G101), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n519), .B(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT29), .B1(new_n517), .B2(new_n522), .ZN(new_n523));
  XOR2_X1   g337(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n379), .B1(new_n503), .B2(new_n509), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n525), .B1(new_n526), .B2(new_n516), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT28), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n516), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n528), .A2(new_n521), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n523), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT70), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT70), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n523), .A2(new_n534), .A3(new_n531), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT71), .ZN(new_n536));
  AOI22_X1  g350(.A1(new_n437), .A2(new_n442), .B1(new_n469), .B2(new_n473), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n537), .A2(new_n509), .A3(new_n379), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n360), .B1(new_n512), .B2(new_n513), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n536), .B(KEYINPUT28), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n530), .A2(KEYINPUT71), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n379), .B1(new_n537), .B2(new_n509), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n529), .B1(new_n542), .B2(new_n516), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n540), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  AND2_X1   g358(.A1(new_n521), .A2(KEYINPUT29), .ZN(new_n545));
  AOI21_X1  g359(.A(G902), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n533), .A2(new_n535), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n515), .A2(new_n521), .A3(new_n516), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT31), .ZN(new_n549));
  INV_X1    g363(.A(new_n530), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n522), .B1(new_n550), .B2(new_n527), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT31), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n515), .A2(new_n552), .A3(new_n521), .A4(new_n516), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n549), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(G472), .A2(G902), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(KEYINPUT69), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT32), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT32), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n554), .A2(new_n559), .A3(new_n556), .ZN(new_n560));
  AOI22_X1  g374(.A1(G472), .A2(new_n547), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT76), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n278), .A2(new_n279), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n297), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n214), .A2(G119), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n344), .A2(G128), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT24), .B(G110), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT23), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n570), .B1(new_n344), .B2(G128), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n214), .A2(KEYINPUT23), .A3(G119), .ZN(new_n572));
  INV_X1    g386(.A(G110), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n571), .A2(new_n572), .A3(new_n573), .A4(new_n566), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT74), .B1(new_n564), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n297), .A3(new_n563), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT74), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n297), .A2(new_n296), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n292), .A2(new_n293), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n279), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n580), .A2(new_n294), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n571), .A2(new_n572), .A3(new_n566), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(G110), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT72), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT72), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n584), .A2(new_n587), .A3(G110), .ZN(new_n588));
  OR2_X1    g402(.A1(new_n567), .A2(new_n568), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  OAI22_X1  g404(.A1(new_n576), .A2(new_n579), .B1(new_n583), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(KEYINPUT22), .B(G137), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n252), .A2(G221), .A3(G234), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n580), .A2(new_n294), .A3(new_n582), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n597), .A2(new_n588), .A3(new_n589), .A4(new_n586), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n598), .B(new_n594), .C1(new_n576), .C2(new_n579), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n189), .B1(G234), .B2(new_n187), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n600), .A2(G902), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n596), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT75), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT75), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n596), .A2(new_n604), .A3(new_n599), .A4(new_n601), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n596), .A2(new_n187), .A3(new_n599), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT25), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT25), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n596), .A2(new_n610), .A3(new_n187), .A4(new_n599), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n611), .A3(new_n600), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n562), .B1(new_n607), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n607), .A2(new_n562), .A3(new_n612), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n561), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n500), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G101), .ZN(G3));
  NAND3_X1  g433(.A1(new_n246), .A2(new_n247), .A3(new_n249), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n247), .A2(G902), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n241), .A2(new_n243), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n241), .A2(new_n243), .A3(KEYINPUT33), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n621), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI22_X1  g440(.A1(new_n333), .A2(new_n310), .B1(new_n620), .B2(new_n626), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n409), .A2(new_n337), .A3(new_n421), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n335), .B(new_n261), .C1(new_n628), .C2(new_n422), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n609), .A2(new_n611), .A3(new_n600), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n633), .A2(KEYINPUT76), .A3(new_n606), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n634), .A2(new_n613), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n459), .A2(new_n460), .B1(new_n466), .B2(new_n467), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n476), .B1(new_n636), .B2(new_n475), .ZN(new_n637));
  INV_X1    g451(.A(new_n477), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n484), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AOI211_X1 g453(.A(G469), .B(G902), .C1(new_n639), .C2(new_n486), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n497), .A2(new_n493), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n426), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n635), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(G472), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n554), .B2(new_n187), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n557), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n632), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  AOI21_X1  g466(.A(KEYINPUT90), .B1(new_n324), .B2(new_n325), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n328), .A2(new_n325), .A3(new_n322), .A4(new_n329), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT90), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n326), .B(new_n331), .C1(new_n653), .C2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n250), .A2(new_n251), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n657), .A2(new_n630), .A3(new_n310), .A4(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n649), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT35), .B(G107), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT91), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n661), .B(new_n663), .ZN(G9));
  NAND2_X1  g478(.A1(new_n591), .A2(KEYINPUT92), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n591), .A2(KEYINPUT92), .ZN(new_n667));
  OAI22_X1  g481(.A1(new_n666), .A2(new_n667), .B1(KEYINPUT36), .B2(new_n595), .ZN(new_n668));
  INV_X1    g482(.A(new_n667), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n595), .A2(KEYINPUT36), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n669), .A2(new_n670), .A3(new_n665), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n668), .A2(new_n671), .A3(new_n601), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n612), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NOR4_X1   g488(.A1(new_n334), .A2(new_n499), .A3(new_n648), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT37), .B(G110), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G12));
  NOR3_X1   g491(.A1(new_n561), .A2(new_n642), .A3(new_n674), .ZN(new_n678));
  INV_X1    g492(.A(G900), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n256), .B1(new_n258), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n309), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n657), .A2(new_n425), .A3(new_n681), .A4(new_n658), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(KEYINPUT93), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT93), .ZN(new_n684));
  INV_X1    g498(.A(new_n680), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n310), .A2(new_n685), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n330), .A2(KEYINPUT85), .A3(KEYINPUT20), .ZN(new_n687));
  AOI21_X1  g501(.A(KEYINPUT85), .B1(new_n330), .B2(KEYINPUT20), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n654), .B(new_n655), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n686), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n335), .B1(new_n628), .B2(new_n422), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n251), .B2(new_n250), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n684), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n678), .B1(new_n683), .B2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT94), .B(G128), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G30));
  XOR2_X1   g511(.A(new_n680), .B(KEYINPUT39), .Z(new_n698));
  NAND3_X1  g512(.A1(new_n498), .A2(new_n426), .A3(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(KEYINPUT96), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT40), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n699), .A2(KEYINPUT96), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n703), .ZN(new_n705));
  OAI21_X1  g519(.A(KEYINPUT40), .B1(new_n705), .B2(new_n700), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n673), .A2(new_n336), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n423), .A2(KEYINPUT38), .A3(new_n424), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT38), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n709), .B1(new_n628), .B2(new_n422), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n707), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n333), .A2(new_n310), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n711), .A2(new_n712), .A3(new_n658), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n522), .B1(new_n515), .B2(new_n516), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n542), .A2(new_n516), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n187), .B1(new_n715), .B2(new_n521), .ZN(new_n716));
  OAI21_X1  g530(.A(G472), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n560), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n559), .B1(new_n554), .B2(new_n556), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT95), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OAI211_X1 g536(.A(KEYINPUT95), .B(new_n717), .C1(new_n718), .C2(new_n719), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n704), .A2(new_n706), .A3(new_n713), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G143), .ZN(G45));
  NOR3_X1   g540(.A1(new_n561), .A2(new_n499), .A3(new_n674), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n626), .A2(new_n620), .ZN(new_n728));
  INV_X1    g542(.A(new_n332), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n687), .A2(new_n688), .A3(new_n729), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n728), .B(new_n685), .C1(new_n730), .C2(new_n309), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G146), .ZN(G48));
  OAI21_X1  g548(.A(new_n187), .B1(new_n487), .B2(new_n490), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(G469), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(new_n426), .A3(new_n491), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n544), .A2(new_n545), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n187), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n534), .B1(new_n523), .B2(new_n531), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n645), .B1(new_n742), .B2(new_n535), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n718), .A2(new_n719), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n635), .B(new_n738), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n631), .ZN(new_n746));
  XOR2_X1   g560(.A(KEYINPUT41), .B(G113), .Z(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G15));
  NOR2_X1   g562(.A1(new_n745), .A2(new_n659), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n195), .ZN(G18));
  OAI21_X1  g564(.A(new_n673), .B1(new_n743), .B2(new_n744), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n737), .A2(new_n692), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n752), .A2(new_n310), .A3(new_n262), .A4(new_n333), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n344), .ZN(G21));
  NAND3_X1  g569(.A1(new_n712), .A2(new_n425), .A3(new_n658), .ZN(new_n756));
  AND4_X1   g570(.A1(new_n426), .A2(new_n736), .A3(new_n491), .A4(new_n261), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n540), .B(new_n522), .C1(new_n541), .C2(new_n543), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n549), .A3(new_n553), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT97), .B1(new_n759), .B2(new_n556), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n646), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT98), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n762), .B1(new_n633), .B2(new_n606), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n607), .A2(KEYINPUT98), .A3(new_n612), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n759), .A2(KEYINPUT97), .A3(new_n556), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n757), .A2(new_n761), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n756), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g582(.A(KEYINPUT99), .B(G122), .Z(new_n769));
  XNOR2_X1  g583(.A(new_n768), .B(new_n769), .ZN(G24));
  INV_X1    g584(.A(KEYINPUT100), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n731), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n761), .A2(new_n766), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n674), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n712), .A2(KEYINPUT100), .A3(new_n728), .A4(new_n685), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n772), .A2(new_n752), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G125), .ZN(G27));
  NOR3_X1   g591(.A1(new_n628), .A2(new_n422), .A3(new_n336), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n426), .A3(new_n498), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n561), .A2(new_n616), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n772), .A2(new_n780), .A3(new_n775), .ZN(new_n781));
  XOR2_X1   g595(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n765), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n561), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n423), .A2(new_n335), .A3(new_n424), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n642), .A2(new_n786), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n787), .A2(KEYINPUT42), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n772), .A2(new_n775), .A3(new_n785), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n783), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g604(.A(KEYINPUT102), .B(G131), .Z(new_n791));
  XNOR2_X1  g605(.A(new_n790), .B(new_n791), .ZN(G33));
  OAI211_X1 g606(.A(new_n787), .B(new_n635), .C1(new_n743), .C2(new_n744), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n691), .A2(new_n658), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XOR2_X1   g609(.A(KEYINPUT103), .B(G134), .Z(new_n796));
  XNOR2_X1  g610(.A(new_n795), .B(new_n796), .ZN(G36));
  AOI21_X1  g611(.A(KEYINPUT45), .B1(new_n495), .B2(new_n496), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n798), .A2(new_n427), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n495), .A2(KEYINPUT45), .A3(new_n496), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n492), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n801), .A2(KEYINPUT46), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n491), .B1(new_n801), .B2(KEYINPUT46), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n804), .A2(new_n426), .A3(new_n698), .A4(new_n778), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n554), .A2(new_n556), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n646), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(new_n674), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT106), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n333), .A2(new_n728), .A3(new_n310), .ZN(new_n810));
  XOR2_X1   g624(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(KEYINPUT105), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT43), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n812), .B1(new_n813), .B2(new_n810), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT105), .B1(new_n810), .B2(new_n811), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n809), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT44), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n805), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n809), .B(KEYINPUT44), .C1(new_n814), .C2(new_n815), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G137), .ZN(G39));
  NAND4_X1  g635(.A1(new_n732), .A2(new_n561), .A3(new_n616), .A4(new_n778), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n804), .A2(KEYINPUT47), .A3(new_n426), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n426), .B1(new_n802), .B2(new_n803), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT47), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n822), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(KEYINPUT107), .B(G140), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n827), .B(new_n828), .ZN(G42));
  OR2_X1    g643(.A1(new_n814), .A2(new_n815), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n830), .A2(new_n256), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n737), .A2(new_n786), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(new_n774), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n724), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n832), .A2(new_n635), .A3(new_n256), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OR3_X1    g650(.A1(new_n836), .A2(new_n712), .A3(new_n728), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n773), .A2(new_n784), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n831), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n736), .A2(new_n491), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n823), .B(new_n826), .C1(new_n426), .C2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n778), .ZN(new_n843));
  OR2_X1    g657(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n838), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n738), .A2(new_n336), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n846), .A2(KEYINPUT113), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n846), .A2(KEYINPUT113), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n708), .A2(new_n710), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n847), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n831), .A2(new_n839), .A3(new_n851), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT50), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT51), .ZN(new_n854));
  OR3_X1    g668(.A1(new_n845), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n854), .B1(new_n845), .B2(new_n853), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n834), .A2(new_n627), .A3(new_n835), .ZN(new_n857));
  INV_X1    g671(.A(new_n752), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n253), .B(new_n857), .C1(new_n840), .C2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n831), .A2(new_n832), .ZN(new_n860));
  INV_X1    g674(.A(new_n785), .ZN(new_n861));
  OR3_X1    g675(.A1(new_n860), .A2(KEYINPUT48), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT48), .B1(new_n860), .B2(new_n861), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n859), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n855), .A2(new_n856), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT110), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n745), .B1(new_n631), .B2(new_n659), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n658), .A2(new_n674), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n868), .B1(new_n743), .B2(new_n744), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n643), .A2(new_n657), .A3(new_n681), .A4(new_n778), .ZN(new_n870));
  OAI22_X1  g684(.A1(new_n793), .A2(new_n794), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI22_X1  g685(.A1(new_n751), .A2(new_n753), .B1(new_n756), .B2(new_n767), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n867), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n772), .A2(new_n774), .A3(new_n775), .A4(new_n787), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n790), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT108), .ZN(new_n876));
  INV_X1    g690(.A(new_n658), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n876), .B1(new_n712), .B2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n333), .A2(new_n658), .A3(KEYINPUT108), .A4(new_n310), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n635), .A2(new_n643), .A3(new_n630), .A4(new_n807), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n500), .A2(new_n807), .A3(new_n673), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT109), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n881), .B1(new_n878), .B2(new_n879), .ZN(new_n887));
  OAI21_X1  g701(.A(KEYINPUT109), .B1(new_n887), .B2(new_n675), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n632), .A2(new_n649), .B1(new_n500), .B2(new_n617), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n886), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n866), .B1(new_n875), .B2(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n886), .A2(new_n888), .A3(new_n889), .ZN(new_n892));
  INV_X1    g706(.A(new_n871), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n617), .B(new_n738), .C1(new_n632), .C2(new_n660), .ZN(new_n894));
  INV_X1    g708(.A(new_n872), .ZN(new_n895));
  AND4_X1   g709(.A1(new_n874), .A2(new_n893), .A3(new_n894), .A4(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n892), .A2(new_n896), .A3(KEYINPUT110), .A4(new_n790), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n891), .A2(new_n897), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n712), .A2(new_n425), .A3(new_n658), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n642), .A2(new_n673), .A3(new_n680), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n724), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n695), .A2(new_n776), .A3(new_n733), .A4(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT52), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT111), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n682), .A2(KEYINPUT93), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n691), .A2(new_n684), .A3(new_n693), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI22_X1  g722(.A1(new_n908), .A2(new_n678), .B1(new_n732), .B2(new_n727), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n909), .A2(KEYINPUT52), .A3(new_n776), .A4(new_n901), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n904), .A2(new_n905), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n902), .A2(KEYINPUT111), .A3(new_n903), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT53), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n898), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n904), .A2(new_n910), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT112), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n904), .A2(KEYINPUT112), .A3(new_n910), .ZN(new_n919));
  AOI22_X1  g733(.A1(new_n918), .A2(new_n919), .B1(new_n891), .B2(new_n897), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n915), .B(KEYINPUT54), .C1(new_n920), .C2(new_n914), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT54), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n875), .A2(new_n890), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n923), .A2(new_n911), .A3(KEYINPUT53), .A4(new_n912), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n922), .B(new_n924), .C1(new_n920), .C2(KEYINPUT53), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n921), .A2(new_n925), .ZN(new_n926));
  OAI22_X1  g740(.A1(new_n865), .A2(new_n926), .B1(G952), .B2(G953), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n841), .B(KEYINPUT49), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n765), .A2(new_n335), .A3(new_n426), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n928), .A2(new_n929), .A3(new_n850), .ZN(new_n930));
  INV_X1    g744(.A(new_n810), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n834), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n927), .A2(new_n932), .ZN(G75));
  NAND2_X1  g747(.A1(new_n384), .A2(new_n408), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(new_n407), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT55), .Z(new_n936));
  NOR2_X1   g750(.A1(new_n936), .A2(KEYINPUT56), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n918), .A2(new_n919), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT53), .B1(new_n938), .B2(new_n898), .ZN(new_n939));
  INV_X1    g753(.A(new_n924), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(G210), .A2(G902), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n937), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n252), .A2(G952), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT114), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n947), .B1(new_n941), .B2(new_n942), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT56), .ZN(new_n949));
  INV_X1    g763(.A(new_n942), .ZN(new_n950));
  OAI211_X1 g764(.A(KEYINPUT114), .B(new_n950), .C1(new_n939), .C2(new_n940), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n946), .B1(new_n952), .B2(new_n936), .ZN(G51));
  XNOR2_X1  g767(.A(new_n492), .B(KEYINPUT57), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n938), .A2(new_n898), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n914), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n922), .B1(new_n956), .B2(new_n924), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n939), .A2(KEYINPUT54), .A3(new_n940), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n954), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n487), .A2(new_n490), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n941), .A2(new_n187), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n963), .A2(new_n800), .A3(new_n799), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n944), .B1(new_n962), .B2(new_n964), .ZN(G54));
  AND2_X1   g779(.A1(KEYINPUT58), .A2(G475), .ZN(new_n966));
  OAI211_X1 g780(.A(G902), .B(new_n966), .C1(new_n939), .C2(new_n940), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT115), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n328), .A2(new_n329), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n945), .B1(new_n967), .B2(new_n969), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n968), .B1(new_n967), .B2(new_n969), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(G60));
  NAND2_X1  g787(.A1(G478), .A2(G902), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT59), .Z(new_n975));
  AOI21_X1  g789(.A(new_n975), .B1(new_n921), .B2(new_n925), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n624), .A2(new_n625), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n945), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n977), .A2(new_n975), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n957), .B2(new_n958), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(KEYINPUT116), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT116), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n983), .B(new_n980), .C1(new_n957), .C2(new_n958), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n979), .B1(new_n982), .B2(new_n984), .ZN(G63));
  NAND2_X1  g799(.A1(new_n596), .A2(new_n599), .ZN(new_n986));
  NAND2_X1  g800(.A1(G217), .A2(G902), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT119), .ZN(new_n988));
  XOR2_X1   g802(.A(KEYINPUT118), .B(KEYINPUT60), .Z(new_n989));
  XOR2_X1   g803(.A(new_n988), .B(new_n989), .Z(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n986), .B1(new_n941), .B2(new_n991), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n668), .A2(new_n671), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n993), .B(new_n990), .C1(new_n939), .C2(new_n940), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n992), .A2(KEYINPUT61), .A3(new_n945), .A4(new_n994), .ZN(new_n995));
  AND3_X1   g809(.A1(new_n992), .A2(new_n945), .A3(new_n994), .ZN(new_n996));
  XOR2_X1   g810(.A(KEYINPUT117), .B(KEYINPUT61), .Z(new_n997));
  OAI21_X1  g811(.A(new_n995), .B1(new_n996), .B2(new_n997), .ZN(G66));
  NOR2_X1   g812(.A1(new_n867), .A2(new_n872), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n886), .A2(new_n888), .A3(new_n999), .A4(new_n889), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT120), .Z(new_n1001));
  NOR2_X1   g815(.A1(new_n1001), .A2(G953), .ZN(new_n1002));
  OAI21_X1  g816(.A(G953), .B1(new_n259), .B2(new_n401), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT121), .Z(new_n1004));
  NOR2_X1   g818(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT122), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n934), .B1(G898), .B2(new_n252), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT122), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1005), .B(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(new_n1007), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1009), .A2(new_n1012), .ZN(G69));
  NOR2_X1   g827(.A1(new_n880), .A2(new_n627), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n617), .A2(new_n701), .A3(new_n703), .A4(new_n778), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI211_X1 g830(.A(new_n1016), .B(new_n827), .C1(new_n818), .C2(new_n819), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n725), .A2(new_n695), .A3(new_n776), .A4(new_n733), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT62), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1018), .B(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT123), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1017), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1021), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n252), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AND2_X1   g839(.A1(new_n510), .A2(new_n514), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1026), .B(new_n316), .Z(new_n1027));
  INV_X1    g841(.A(new_n1027), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1025), .A2(KEYINPUT124), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT124), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n827), .B1(new_n818), .B2(new_n819), .ZN(new_n1031));
  INV_X1    g845(.A(new_n1016), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g847(.A(new_n1018), .B(KEYINPUT62), .ZN(new_n1034));
  OAI21_X1  g848(.A(KEYINPUT123), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g849(.A(G953), .B1(new_n1035), .B2(new_n1022), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1030), .B1(new_n1036), .B2(new_n1027), .ZN(new_n1037));
  AND2_X1   g851(.A1(new_n909), .A2(new_n776), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n804), .A2(new_n426), .A3(new_n698), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n899), .A2(new_n785), .ZN(new_n1040));
  OAI22_X1  g854(.A1(new_n1039), .A2(new_n1040), .B1(new_n793), .B2(new_n794), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n1041), .B1(new_n783), .B2(new_n789), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n1031), .A2(new_n1038), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1043), .A2(KEYINPUT126), .ZN(new_n1044));
  INV_X1    g858(.A(KEYINPUT126), .ZN(new_n1045));
  NAND4_X1  g859(.A1(new_n1031), .A2(new_n1045), .A3(new_n1038), .A4(new_n1042), .ZN(new_n1046));
  AOI21_X1  g860(.A(G953), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g861(.A1(new_n252), .A2(G900), .ZN(new_n1048));
  OAI21_X1  g862(.A(new_n1027), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n1029), .A2(new_n1037), .A3(new_n1049), .ZN(new_n1050));
  OAI21_X1  g864(.A(G953), .B1(new_n482), .B2(new_n679), .ZN(new_n1051));
  XNOR2_X1  g865(.A(new_n1051), .B(KEYINPUT125), .ZN(new_n1052));
  XNOR2_X1  g866(.A(new_n1050), .B(new_n1052), .ZN(G72));
  NAND3_X1  g867(.A1(new_n1044), .A2(new_n1001), .A3(new_n1046), .ZN(new_n1054));
  NAND2_X1  g868(.A1(G472), .A2(G902), .ZN(new_n1055));
  XOR2_X1   g869(.A(new_n1055), .B(KEYINPUT63), .Z(new_n1056));
  NAND2_X1  g870(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g871(.A1(new_n517), .A2(new_n521), .ZN(new_n1058));
  AOI21_X1  g872(.A(new_n944), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AND3_X1   g873(.A1(new_n1035), .A2(new_n1001), .A3(new_n1022), .ZN(new_n1060));
  INV_X1    g874(.A(new_n1056), .ZN(new_n1061));
  OAI21_X1  g875(.A(new_n714), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NOR3_X1   g876(.A1(new_n1058), .A2(new_n714), .A3(new_n1061), .ZN(new_n1063));
  OAI211_X1 g877(.A(new_n915), .B(new_n1063), .C1(new_n920), .C2(new_n914), .ZN(new_n1064));
  NAND3_X1  g878(.A1(new_n1059), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g879(.A1(new_n1065), .A2(KEYINPUT127), .ZN(new_n1066));
  INV_X1    g880(.A(KEYINPUT127), .ZN(new_n1067));
  NAND4_X1  g881(.A1(new_n1059), .A2(new_n1062), .A3(new_n1067), .A4(new_n1064), .ZN(new_n1068));
  NAND2_X1  g882(.A1(new_n1066), .A2(new_n1068), .ZN(G57));
endmodule


