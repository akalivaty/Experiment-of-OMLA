//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n787, new_n788, new_n789, new_n790, new_n791, new_n793,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n988, new_n989, new_n990, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1028, new_n1029, new_n1030;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT3), .ZN(new_n203));
  XNOR2_X1  g002(.A(G155gat), .B(G162gat), .ZN(new_n204));
  INV_X1    g003(.A(G141gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G148gat), .ZN(new_n206));
  INV_X1    g005(.A(G148gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G141gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  AOI22_X1  g008(.A1(new_n206), .A2(new_n208), .B1(KEYINPUT2), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT77), .ZN(new_n211));
  OAI211_X1 g010(.A(KEYINPUT78), .B(new_n204), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT78), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n209), .A2(KEYINPUT2), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n207), .A2(G141gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n205), .A2(G148gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n213), .B1(new_n217), .B2(KEYINPUT77), .ZN(new_n218));
  XOR2_X1   g017(.A(G155gat), .B(G162gat), .Z(new_n219));
  AOI21_X1  g018(.A(new_n219), .B1(new_n217), .B2(new_n213), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n203), .B(new_n212), .C1(new_n218), .C2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT29), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT73), .ZN(new_n224));
  NAND2_X1  g023(.A1(G211gat), .A2(G218gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT22), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(G197gat), .A2(G204gat), .ZN(new_n228));
  AND2_X1   g027(.A1(G197gat), .A2(G204gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT72), .ZN(new_n231));
  XNOR2_X1  g030(.A(G211gat), .B(G218gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n232), .B1(new_n230), .B2(new_n231), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n224), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(G211gat), .A2(G218gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(G211gat), .A2(G218gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n228), .ZN(new_n241));
  NAND2_X1  g040(.A1(G197gat), .A2(G204gat), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n239), .B1(new_n243), .B2(KEYINPUT72), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n244), .A2(new_n233), .A3(KEYINPUT73), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n236), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n223), .A2(new_n246), .ZN(new_n247));
  AND2_X1   g046(.A1(G228gat), .A2(G233gat), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n244), .A2(new_n233), .A3(new_n222), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n203), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT78), .B1(new_n210), .B2(new_n211), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n204), .B1(new_n210), .B2(KEYINPUT78), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(new_n212), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n249), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n247), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n229), .A2(new_n228), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n232), .B1(new_n259), .B2(new_n240), .ZN(new_n260));
  XNOR2_X1  g059(.A(G197gat), .B(G204gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n239), .A2(new_n261), .A3(new_n227), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n260), .A2(new_n262), .A3(new_n222), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n254), .A2(new_n212), .B1(new_n263), .B2(new_n203), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(KEYINPUT79), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n247), .A2(KEYINPUT80), .ZN(new_n266));
  AOI22_X1  g065(.A1(new_n221), .A2(new_n222), .B1(new_n236), .B2(new_n245), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT80), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n265), .A2(new_n266), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n258), .B1(new_n270), .B2(new_n249), .ZN(new_n271));
  XOR2_X1   g070(.A(KEYINPUT81), .B(G22gat), .Z(new_n272));
  OAI21_X1  g071(.A(new_n202), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G141gat), .B(G148gat), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n209), .A2(KEYINPUT2), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT77), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n213), .B1(new_n274), .B2(new_n275), .ZN(new_n277));
  AOI22_X1  g076(.A1(KEYINPUT78), .A2(new_n276), .B1(new_n277), .B2(new_n204), .ZN(new_n278));
  INV_X1    g077(.A(new_n212), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n260), .A2(new_n262), .A3(new_n222), .ZN(new_n280));
  OAI22_X1  g079(.A1(new_n278), .A2(new_n279), .B1(new_n280), .B2(KEYINPUT3), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT79), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT79), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n264), .A2(new_n283), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n282), .B(new_n284), .C1(new_n267), .C2(new_n268), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n247), .A2(KEYINPUT80), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n249), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(new_n257), .ZN(new_n288));
  INV_X1    g087(.A(new_n272), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(KEYINPUT82), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n287), .A2(new_n272), .A3(new_n257), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n273), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G78gat), .B(G106gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(KEYINPUT31), .B(G50gat), .ZN(new_n294));
  XOR2_X1   g093(.A(new_n293), .B(new_n294), .Z(new_n295));
  NAND2_X1  g094(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n295), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G22gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n271), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT83), .ZN(new_n304));
  AND3_X1   g103(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G190gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT64), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT64), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G190gat), .ZN(new_n311));
  INV_X1    g110(.A(G183gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n309), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT23), .ZN(new_n315));
  NOR3_X1   g114(.A1(new_n315), .A2(G169gat), .A3(G176gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(G169gat), .A2(G176gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT23), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n316), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n314), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT25), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n317), .B1(KEYINPUT23), .B2(new_n319), .ZN(new_n324));
  NOR3_X1   g123(.A1(new_n324), .A2(KEYINPUT25), .A3(new_n316), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n307), .B1(G183gat), .B2(G190gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n309), .A2(new_n311), .A3(KEYINPUT28), .ZN(new_n328));
  AND2_X1   g127(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT65), .B1(new_n312), .B2(KEYINPUT66), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT27), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI211_X1 g134(.A(KEYINPUT65), .B(KEYINPUT27), .C1(new_n312), .C2(KEYINPUT66), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT64), .B(G190gat), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT65), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n329), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n335), .A2(new_n336), .A3(new_n337), .A4(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT28), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n332), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT26), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n318), .A2(new_n343), .A3(new_n319), .ZN(new_n344));
  NAND2_X1  g143(.A1(G183gat), .A2(G190gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n317), .A2(KEYINPUT26), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n323), .B(new_n327), .C1(new_n342), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(new_n222), .ZN(new_n349));
  NAND2_X1  g148(.A1(G226gat), .A2(G233gat), .ZN(new_n350));
  XOR2_X1   g149(.A(new_n350), .B(KEYINPUT74), .Z(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n348), .A2(new_n351), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n353), .A2(new_n246), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n246), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n351), .B1(new_n348), .B2(new_n222), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n341), .ZN(new_n358));
  INV_X1    g157(.A(new_n332), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n347), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n322), .A2(KEYINPUT25), .B1(new_n325), .B2(new_n326), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n352), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n356), .B1(new_n357), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n355), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G8gat), .B(G36gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(G64gat), .B(G92gat), .ZN(new_n368));
  XOR2_X1   g167(.A(new_n367), .B(new_n368), .Z(new_n369));
  NOR2_X1   g168(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n246), .B1(new_n353), .B2(new_n354), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n357), .A2(new_n364), .A3(new_n356), .ZN(new_n372));
  OAI211_X1 g171(.A(KEYINPUT30), .B(new_n369), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT75), .ZN(new_n374));
  INV_X1    g173(.A(new_n369), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n375), .B1(new_n355), .B2(new_n365), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT75), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT30), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n370), .B1(new_n374), .B2(new_n378), .ZN(new_n379));
  OR2_X1    g178(.A1(new_n376), .A2(KEYINPUT76), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT30), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n376), .A2(KEYINPUT76), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT3), .B1(new_n278), .B2(new_n279), .ZN(new_n384));
  INV_X1    g183(.A(G113gat), .ZN(new_n385));
  INV_X1    g184(.A(G120gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT1), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n389), .B1(G113gat), .B2(G120gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G127gat), .B(G134gat), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n388), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(G134gat), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n394), .A2(G127gat), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(G127gat), .ZN(new_n396));
  OAI22_X1  g195(.A1(new_n387), .A2(new_n390), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n384), .A2(new_n221), .A3(new_n399), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n254), .A2(new_n212), .A3(new_n398), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT4), .ZN(new_n402));
  NAND2_X1  g201(.A1(G225gat), .A2(G233gat), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n254), .A2(new_n212), .A3(new_n398), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT4), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n400), .A2(new_n402), .A3(new_n403), .A4(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n403), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n398), .B1(new_n254), .B2(new_n212), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n408), .B1(new_n401), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT5), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n404), .B(KEYINPUT4), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n413), .A2(KEYINPUT5), .A3(new_n403), .A4(new_n400), .ZN(new_n414));
  XNOR2_X1  g213(.A(G1gat), .B(G29gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(KEYINPUT0), .ZN(new_n416));
  XNOR2_X1  g215(.A(G57gat), .B(G85gat), .ZN(new_n417));
  XOR2_X1   g216(.A(new_n416), .B(new_n417), .Z(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n412), .A2(new_n414), .A3(KEYINPUT6), .A4(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n412), .A2(new_n414), .A3(new_n419), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT6), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n419), .B1(new_n412), .B2(new_n414), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n420), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n379), .A2(new_n383), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n301), .B1(new_n292), .B2(new_n295), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT83), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n304), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT37), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n369), .B1(new_n366), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n355), .A2(new_n365), .A3(KEYINPUT37), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT86), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(KEYINPUT87), .B(KEYINPUT38), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n355), .A2(new_n365), .A3(KEYINPUT86), .A4(KEYINPUT37), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n432), .A2(new_n435), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n376), .A2(KEYINPUT76), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT76), .ZN(new_n440));
  AOI211_X1 g239(.A(new_n440), .B(new_n375), .C1(new_n355), .C2(new_n365), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n436), .B1(new_n432), .B2(new_n433), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT85), .B1(new_n423), .B2(new_n424), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n412), .A2(new_n414), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n418), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT85), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n448), .A2(new_n449), .A3(new_n422), .A4(new_n421), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n446), .A2(new_n420), .A3(new_n450), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n445), .A2(new_n451), .B1(new_n296), .B2(new_n302), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n413), .A2(new_n400), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT39), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n453), .A2(new_n454), .A3(new_n408), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n418), .ZN(new_n456));
  OR2_X1    g255(.A1(new_n401), .A2(new_n409), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT39), .B1(new_n457), .B2(new_n408), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n458), .B1(new_n408), .B2(new_n453), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT40), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT84), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT40), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n462), .B(new_n463), .C1(new_n456), .C2(new_n459), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n461), .A2(new_n421), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT84), .B1(new_n460), .B2(KEYINPUT40), .ZN(new_n466));
  NOR3_X1   g265(.A1(new_n439), .A2(new_n441), .A3(KEYINPUT30), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n373), .A2(KEYINPUT75), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n377), .B1(new_n376), .B2(KEYINPUT30), .ZN(new_n469));
  OAI22_X1  g268(.A1(new_n468), .A2(new_n469), .B1(new_n369), .B2(new_n366), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n465), .B(new_n466), .C1(new_n467), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n452), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT69), .ZN(new_n473));
  XOR2_X1   g272(.A(G15gat), .B(G43gat), .Z(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(KEYINPUT67), .ZN(new_n475));
  XOR2_X1   g274(.A(G71gat), .B(G99gat), .Z(new_n476));
  XNOR2_X1  g275(.A(new_n475), .B(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(G227gat), .ZN(new_n478));
  INV_X1    g277(.A(G233gat), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n323), .A2(new_n327), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n347), .B1(new_n358), .B2(new_n359), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n399), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n363), .B(new_n398), .C1(new_n342), .C2(new_n347), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n481), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n477), .B1(new_n486), .B2(KEYINPUT33), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT32), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n484), .A2(new_n485), .ZN(new_n491));
  AOI221_X4 g290(.A(new_n488), .B1(KEYINPUT33), .B2(new_n477), .C1(new_n491), .C2(new_n480), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n473), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n484), .A2(new_n481), .A3(new_n485), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT68), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT34), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT34), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n495), .B(new_n498), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n499), .B(new_n473), .C1(new_n490), .C2(new_n492), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(new_n500), .A3(KEYINPUT36), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT70), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n497), .A2(new_n500), .A3(KEYINPUT70), .A4(KEYINPUT36), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n490), .A2(new_n492), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(new_n496), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n499), .B1(new_n490), .B2(new_n492), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XOR2_X1   g308(.A(KEYINPUT71), .B(KEYINPUT36), .Z(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n430), .A2(new_n472), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n426), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n500), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n303), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT35), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n379), .A2(new_n383), .A3(new_n507), .A4(new_n508), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT35), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n446), .A2(new_n420), .A3(new_n450), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n520), .A2(new_n303), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n513), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(G50gat), .ZN(new_n526));
  AND2_X1   g325(.A1(KEYINPUT90), .A2(G43gat), .ZN(new_n527));
  NOR2_X1   g326(.A1(KEYINPUT90), .A2(G43gat), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(G43gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(G50gat), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT15), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT14), .ZN(new_n533));
  INV_X1    g332(.A(G36gat), .ZN(new_n534));
  NOR3_X1   g333(.A1(new_n533), .A2(new_n534), .A3(G29gat), .ZN(new_n535));
  INV_X1    g334(.A(G29gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT14), .ZN(new_n537));
  AOI21_X1  g336(.A(G36gat), .B1(new_n533), .B2(G29gat), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G43gat), .B(G50gat), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT15), .B1(new_n540), .B2(KEYINPUT89), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n526), .A2(G43gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n531), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT89), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI22_X1  g344(.A1(new_n532), .A2(new_n539), .B1(new_n541), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT17), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n538), .A2(new_n537), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n548), .B1(new_n534), .B2(new_n537), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n540), .A2(KEYINPUT89), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n543), .A2(new_n544), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n549), .A2(KEYINPUT15), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n546), .A2(new_n547), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT91), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n546), .A2(KEYINPUT91), .A3(new_n552), .A4(new_n547), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G15gat), .B(G22gat), .ZN(new_n558));
  INV_X1    g357(.A(G1gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT16), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n561), .B1(G1gat), .B2(new_n558), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(G8gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n552), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n563), .B1(KEYINPUT17), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n564), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n557), .A2(new_n565), .B1(new_n566), .B2(new_n563), .ZN(new_n567));
  NAND2_X1  g366(.A1(G229gat), .A2(G233gat), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n567), .A2(KEYINPUT92), .A3(KEYINPUT18), .A4(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n563), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(new_n564), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n566), .A2(new_n563), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n568), .B(KEYINPUT13), .Z(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n569), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G113gat), .B(G141gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(G197gat), .ZN(new_n578));
  XOR2_X1   g377(.A(KEYINPUT11), .B(G169gat), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(KEYINPUT88), .B(KEYINPUT12), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT18), .B1(new_n567), .B2(new_n568), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT93), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n557), .A2(new_n565), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n586), .A2(new_n572), .A3(KEYINPUT18), .A4(new_n568), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT92), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n586), .A2(new_n568), .A3(new_n572), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT18), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT93), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n576), .A2(new_n585), .A3(new_n589), .A4(new_n593), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n589), .A2(new_n592), .A3(new_n569), .A4(new_n575), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(new_n582), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT100), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT9), .ZN(new_n599));
  INV_X1    g398(.A(G71gat), .ZN(new_n600));
  INV_X1    g399(.A(G78gat), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT94), .ZN(new_n603));
  XOR2_X1   g402(.A(G57gat), .B(G64gat), .Z(new_n604));
  XNOR2_X1  g403(.A(G71gat), .B(G78gat), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT94), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n606), .B(new_n599), .C1(new_n600), .C2(new_n601), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n603), .A2(new_n604), .A3(new_n605), .A4(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(G71gat), .B(G78gat), .Z(new_n609));
  XNOR2_X1  g408(.A(G57gat), .B(G64gat), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n609), .B1(new_n599), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT95), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n608), .A2(KEYINPUT95), .A3(new_n611), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT21), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n570), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G127gat), .B(G155gat), .Z(new_n620));
  NAND2_X1  g419(.A1(G231gat), .A2(G233gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n619), .B(new_n622), .Z(new_n623));
  XOR2_X1   g422(.A(G183gat), .B(G211gat), .Z(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(KEYINPUT96), .B(KEYINPUT21), .Z(new_n628));
  AOI21_X1  g427(.A(new_n627), .B1(new_n617), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n617), .A2(new_n628), .A3(new_n627), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n625), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n630), .A2(new_n625), .A3(new_n631), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n623), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n619), .B(new_n622), .ZN(new_n636));
  INV_X1    g435(.A(new_n634), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n636), .B1(new_n637), .B2(new_n632), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  AND2_X1   g438(.A1(G232gat), .A2(G233gat), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n640), .A2(KEYINPUT41), .ZN(new_n641));
  XNOR2_X1  g440(.A(G134gat), .B(G162gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(G85gat), .ZN(new_n645));
  INV_X1    g444(.A(G92gat), .ZN(new_n646));
  OAI22_X1  g445(.A1(new_n645), .A2(new_n646), .B1(KEYINPUT97), .B2(KEYINPUT7), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT97), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT7), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n648), .A2(new_n649), .A3(G85gat), .A4(G92gat), .ZN(new_n650));
  NAND2_X1  g449(.A1(KEYINPUT97), .A2(KEYINPUT7), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n647), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  OR2_X1    g451(.A1(G99gat), .A2(G106gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(G99gat), .A2(G106gat), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n653), .A2(KEYINPUT98), .A3(new_n654), .ZN(new_n655));
  AOI22_X1  g454(.A1(KEYINPUT8), .A2(new_n654), .B1(new_n645), .B2(new_n646), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n652), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT98), .B1(new_n653), .B2(new_n654), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n658), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n660), .A2(new_n652), .A3(new_n655), .A4(new_n656), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n662), .B1(new_n564), .B2(KEYINPUT17), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n557), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g463(.A(G190gat), .B(G218gat), .Z(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  AOI22_X1  g465(.A1(new_n566), .A2(new_n662), .B1(KEYINPUT41), .B2(new_n640), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n664), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n666), .B1(new_n664), .B2(new_n667), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n644), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n670), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n672), .A2(new_n643), .A3(new_n668), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n639), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(G120gat), .B(G148gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(G176gat), .B(G204gat), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n676), .B(new_n677), .Z(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(G230gat), .A2(G233gat), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT99), .ZN(new_n682));
  AOI22_X1  g481(.A1(new_n659), .A2(new_n661), .B1(new_n611), .B2(new_n608), .ZN(new_n683));
  INV_X1    g482(.A(new_n662), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n683), .B1(new_n616), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n682), .B1(new_n685), .B2(KEYINPUT10), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n608), .A2(KEYINPUT95), .A3(new_n611), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT95), .B1(new_n608), .B2(new_n611), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n659), .B(new_n661), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n662), .A2(new_n612), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT10), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(KEYINPUT99), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n686), .A2(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n617), .A2(new_n684), .A3(new_n692), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n681), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n691), .A2(new_n680), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n679), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT99), .B1(new_n691), .B2(new_n692), .ZN(new_n700));
  AOI211_X1 g499(.A(new_n682), .B(KEYINPUT10), .C1(new_n689), .C2(new_n690), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n696), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n680), .ZN(new_n703));
  INV_X1    g502(.A(new_n698), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(new_n704), .A3(new_n678), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n699), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n598), .B1(new_n675), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n678), .B1(new_n703), .B2(new_n704), .ZN(new_n708));
  AOI211_X1 g507(.A(new_n698), .B(new_n679), .C1(new_n702), .C2(new_n680), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI22_X1  g509(.A1(new_n635), .A2(new_n638), .B1(new_n671), .B2(new_n673), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(new_n711), .A3(KEYINPUT100), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n525), .A2(new_n597), .A3(new_n707), .A4(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(new_n425), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(new_n559), .ZN(G1324gat));
  INV_X1    g514(.A(KEYINPUT42), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n470), .A2(new_n467), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n716), .B1(new_n719), .B2(G8gat), .ZN(new_n720));
  XOR2_X1   g519(.A(KEYINPUT16), .B(G8gat), .Z(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT101), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(KEYINPUT102), .A2(KEYINPUT42), .ZN(new_n724));
  MUX2_X1   g523(.A(KEYINPUT102), .B(new_n724), .S(new_n722), .Z(new_n725));
  AOI22_X1  g524(.A1(new_n720), .A2(new_n723), .B1(new_n718), .B2(new_n725), .ZN(G1325gat));
  OAI21_X1  g525(.A(G15gat), .B1(new_n713), .B2(new_n512), .ZN(new_n727));
  OR2_X1    g526(.A1(new_n509), .A2(G15gat), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(new_n713), .B2(new_n728), .ZN(G1326gat));
  NAND2_X1  g528(.A1(new_n304), .A2(new_n429), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n713), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g530(.A(KEYINPUT43), .B(G22gat), .Z(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(G1327gat));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n515), .B1(new_n296), .B2(new_n302), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n521), .B1(new_n735), .B2(new_n514), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n522), .A2(new_n521), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n737), .A2(new_n427), .A3(new_n519), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT104), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT104), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n427), .A2(new_n426), .A3(new_n515), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n523), .B(new_n740), .C1(new_n521), .C2(new_n741), .ZN(new_n742));
  AOI22_X1  g541(.A1(new_n471), .A2(new_n452), .B1(new_n505), .B2(new_n511), .ZN(new_n743));
  AOI22_X1  g542(.A1(new_n739), .A2(new_n742), .B1(new_n743), .B2(new_n430), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n734), .B1(new_n744), .B2(new_n674), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n674), .B1(new_n513), .B2(new_n524), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT44), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n597), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n749), .A2(new_n639), .A3(new_n706), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT103), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G29gat), .B1(new_n752), .B2(new_n425), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n746), .A2(new_n750), .ZN(new_n754));
  INV_X1    g553(.A(new_n425), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n754), .A2(new_n536), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT45), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n753), .A2(new_n757), .ZN(G1328gat));
  INV_X1    g557(.A(new_n717), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n754), .A2(new_n534), .A3(new_n759), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(KEYINPUT46), .Z(new_n761));
  OAI21_X1  g560(.A(G36gat), .B1(new_n752), .B2(new_n717), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(G1329gat));
  INV_X1    g562(.A(new_n752), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n527), .A2(new_n528), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n512), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n509), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n754), .A2(new_n767), .ZN(new_n768));
  AOI22_X1  g567(.A1(new_n764), .A2(new_n766), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n769), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g569(.A(G50gat), .B1(new_n752), .B2(new_n303), .ZN(new_n771));
  INV_X1    g570(.A(new_n730), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n754), .A2(new_n526), .A3(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n771), .A2(KEYINPUT48), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(G50gat), .B1(new_n752), .B2(new_n730), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n775), .A2(KEYINPUT105), .A3(new_n773), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT48), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n777), .B1(new_n775), .B2(KEYINPUT105), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n774), .B1(new_n776), .B2(new_n778), .ZN(G1331gat));
  NOR4_X1   g578(.A1(new_n744), .A2(new_n597), .A3(new_n675), .A4(new_n710), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n755), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n759), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n783), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n784));
  XOR2_X1   g583(.A(KEYINPUT49), .B(G64gat), .Z(new_n785));
  OAI21_X1  g584(.A(new_n784), .B1(new_n783), .B2(new_n785), .ZN(G1333gat));
  NAND3_X1  g585(.A1(new_n780), .A2(new_n600), .A3(new_n767), .ZN(new_n787));
  INV_X1    g586(.A(new_n512), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n780), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n787), .B1(new_n789), .B2(new_n600), .ZN(new_n790));
  XOR2_X1   g589(.A(KEYINPUT106), .B(KEYINPUT50), .Z(new_n791));
  XNOR2_X1  g590(.A(new_n790), .B(new_n791), .ZN(G1334gat));
  NAND2_X1  g591(.A1(new_n780), .A2(new_n772), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g593(.A(new_n740), .B1(new_n518), .B2(new_n523), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n736), .A2(new_n738), .A3(KEYINPUT104), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n513), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n671), .A2(new_n673), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n597), .A2(new_n639), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n797), .A2(KEYINPUT51), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT109), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT110), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n739), .A2(new_n742), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n674), .B1(new_n804), .B2(new_n513), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n805), .A2(KEYINPUT109), .A3(KEYINPUT51), .A4(new_n799), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n802), .A2(new_n803), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n799), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n803), .B1(new_n802), .B2(new_n806), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(new_n710), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n814), .A2(new_n645), .A3(new_n755), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n706), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(KEYINPUT107), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n747), .B(new_n817), .C1(new_n805), .C2(KEYINPUT44), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT108), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT108), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n745), .A2(new_n820), .A3(new_n747), .A4(new_n817), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(G85gat), .B1(new_n822), .B2(new_n425), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n815), .A2(new_n823), .ZN(G1336gat));
  NOR2_X1   g623(.A1(new_n717), .A2(G92gat), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n706), .B(new_n825), .C1(new_n811), .C2(new_n812), .ZN(new_n826));
  OAI21_X1  g625(.A(G92gat), .B1(new_n818), .B2(new_n717), .ZN(new_n827));
  XOR2_X1   g626(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n819), .A2(new_n759), .A3(new_n821), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(G92gat), .ZN(new_n831));
  INV_X1    g630(.A(new_n799), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n744), .A2(new_n674), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT109), .B1(new_n833), .B2(KEYINPUT51), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n800), .A2(new_n801), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n810), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n717), .A2(G92gat), .A3(new_n710), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n831), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(KEYINPUT111), .B1(new_n839), .B2(KEYINPUT52), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT111), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n842));
  AOI211_X1 g641(.A(new_n841), .B(new_n842), .C1(new_n831), .C2(new_n838), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n829), .B1(new_n840), .B2(new_n843), .ZN(G1337gat));
  INV_X1    g643(.A(G99gat), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n814), .A2(new_n845), .A3(new_n767), .ZN(new_n846));
  OAI21_X1  g645(.A(G99gat), .B1(new_n822), .B2(new_n512), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(G1338gat));
  NOR3_X1   g647(.A1(new_n303), .A2(G106gat), .A3(new_n710), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n849), .B1(new_n811), .B2(new_n812), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(KEYINPUT113), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT113), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n852), .B(new_n849), .C1(new_n811), .C2(new_n812), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n748), .A2(new_n427), .A3(new_n817), .ZN(new_n854));
  AOI21_X1  g653(.A(KEYINPUT53), .B1(new_n854), .B2(G106gat), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n851), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(G106gat), .B1(new_n822), .B2(new_n730), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n836), .A2(new_n849), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT53), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n856), .A2(new_n860), .ZN(G1339gat));
  NAND3_X1  g660(.A1(new_n749), .A2(new_n711), .A3(new_n710), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n678), .B1(new_n697), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n694), .A2(new_n681), .A3(new_n696), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n703), .A2(KEYINPUT54), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n866), .A3(KEYINPUT55), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n705), .ZN(new_n868));
  OAI22_X1  g667(.A1(new_n567), .A2(new_n568), .B1(new_n573), .B2(new_n574), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n580), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n594), .A2(new_n798), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(KEYINPUT55), .B1(new_n864), .B2(new_n866), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n868), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT55), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n695), .B1(new_n686), .B2(new_n693), .ZN(new_n875));
  OAI21_X1  g674(.A(KEYINPUT54), .B1(new_n875), .B2(new_n681), .ZN(new_n876));
  AOI211_X1 g675(.A(new_n680), .B(new_n695), .C1(new_n686), .C2(new_n693), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n702), .A2(new_n863), .A3(new_n680), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n679), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n874), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n597), .A2(new_n881), .A3(new_n705), .A4(new_n867), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT114), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n585), .A2(new_n593), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n589), .A2(new_n569), .A3(new_n575), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n870), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n883), .B1(new_n886), .B2(new_n710), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n706), .A2(new_n594), .A3(KEYINPUT114), .A4(new_n870), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n882), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n873), .B1(new_n889), .B2(new_n674), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n862), .B1(new_n890), .B2(new_n639), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(new_n425), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n759), .A2(new_n427), .A3(new_n515), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(G113gat), .B1(new_n896), .B2(new_n597), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n893), .A2(new_n520), .A3(new_n730), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT115), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n749), .A2(new_n385), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(G1340gat));
  INV_X1    g700(.A(new_n899), .ZN(new_n902));
  OAI21_X1  g701(.A(G120gat), .B1(new_n902), .B2(new_n710), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n706), .A2(new_n386), .ZN(new_n904));
  XOR2_X1   g703(.A(new_n904), .B(KEYINPUT116), .Z(new_n905));
  OAI21_X1  g704(.A(new_n903), .B1(new_n895), .B2(new_n905), .ZN(G1341gat));
  INV_X1    g705(.A(new_n639), .ZN(new_n907));
  OAI21_X1  g706(.A(G127gat), .B1(new_n902), .B2(new_n907), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n907), .A2(G127gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n895), .B2(new_n909), .ZN(G1342gat));
  OAI21_X1  g709(.A(G134gat), .B1(new_n902), .B2(new_n674), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n798), .A2(new_n394), .ZN(new_n912));
  OAI22_X1  g711(.A1(new_n895), .A2(new_n912), .B1(KEYINPUT117), .B2(KEYINPUT56), .ZN(new_n913));
  NAND2_X1  g712(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n914));
  XOR2_X1   g713(.A(new_n913), .B(new_n914), .Z(new_n915));
  NAND2_X1  g714(.A1(new_n911), .A2(new_n915), .ZN(G1343gat));
  NOR3_X1   g715(.A1(new_n788), .A2(new_n425), .A3(new_n759), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT57), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT118), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n919), .B1(new_n878), .B2(new_n880), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n864), .A2(new_n866), .A3(KEYINPUT118), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n920), .A2(new_n874), .A3(new_n921), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n867), .A2(new_n705), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n922), .A2(new_n923), .A3(new_n597), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n706), .A2(new_n594), .A3(new_n870), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n798), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n907), .B1(new_n926), .B2(new_n873), .ZN(new_n927));
  AOI211_X1 g726(.A(new_n918), .B(new_n730), .C1(new_n927), .C2(new_n862), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT57), .B1(new_n891), .B2(new_n427), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n917), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(G141gat), .B1(new_n930), .B2(new_n749), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n788), .A2(new_n759), .A3(new_n303), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n893), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n205), .A3(new_n597), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g735(.A1(new_n933), .A2(new_n207), .A3(new_n706), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n930), .A2(new_n710), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n939), .A2(KEYINPUT59), .A3(new_n207), .ZN(new_n940));
  XOR2_X1   g739(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n941));
  AOI21_X1  g740(.A(new_n918), .B1(new_n891), .B2(new_n427), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n730), .A2(KEYINPUT57), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n707), .A2(new_n712), .A3(new_n749), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT120), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n945), .B(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n944), .B1(new_n927), .B2(new_n947), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n942), .A2(new_n948), .A3(new_n710), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(new_n917), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n941), .B1(new_n950), .B2(G148gat), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n937), .B1(new_n940), .B2(new_n951), .ZN(G1345gat));
  NAND2_X1  g751(.A1(new_n933), .A2(new_n639), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n953), .A2(KEYINPUT121), .ZN(new_n954));
  INV_X1    g753(.A(G155gat), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n955), .B1(new_n953), .B2(KEYINPUT121), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n639), .A2(G155gat), .ZN(new_n957));
  OAI22_X1  g756(.A1(new_n954), .A2(new_n956), .B1(new_n930), .B2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(G1346gat));
  INV_X1    g758(.A(G162gat), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n933), .A2(new_n960), .A3(new_n798), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT122), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n961), .B(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(G162gat), .B1(new_n930), .B2(new_n674), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(KEYINPUT123), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT123), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n963), .A2(new_n967), .A3(new_n964), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n968), .ZN(G1347gat));
  NOR2_X1   g768(.A1(new_n717), .A2(new_n755), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n891), .A2(new_n767), .A3(new_n730), .A4(new_n970), .ZN(new_n971));
  INV_X1    g770(.A(G169gat), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n971), .A2(new_n972), .A3(new_n749), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n892), .A2(new_n755), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n735), .A2(new_n759), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n975), .B(KEYINPUT124), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  INV_X1    g776(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n978), .A2(new_n597), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n973), .B1(new_n979), .B2(new_n972), .ZN(G1348gat));
  OAI21_X1  g779(.A(G176gat), .B1(new_n971), .B2(new_n710), .ZN(new_n981));
  OR2_X1    g780(.A1(new_n710), .A2(G176gat), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n981), .B1(new_n977), .B2(new_n982), .ZN(G1349gat));
  OAI21_X1  g782(.A(G183gat), .B1(new_n971), .B2(new_n907), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n639), .B1(new_n329), .B2(new_n330), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n984), .B1(new_n977), .B2(new_n985), .ZN(new_n986));
  XNOR2_X1  g785(.A(new_n986), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g786(.A(G190gat), .B1(new_n971), .B2(new_n674), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n988), .B(KEYINPUT61), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n978), .A2(new_n337), .A3(new_n798), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(G1351gat));
  NAND4_X1  g790(.A1(new_n974), .A2(new_n759), .A3(new_n427), .A4(new_n512), .ZN(new_n992));
  INV_X1    g791(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g792(.A(G197gat), .B1(new_n993), .B2(new_n597), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n512), .A2(new_n970), .ZN(new_n995));
  NOR3_X1   g794(.A1(new_n942), .A2(new_n948), .A3(new_n995), .ZN(new_n996));
  AND3_X1   g795(.A1(new_n996), .A2(G197gat), .A3(new_n597), .ZN(new_n997));
  NOR2_X1   g796(.A1(new_n994), .A2(new_n997), .ZN(G1352gat));
  NOR2_X1   g797(.A1(new_n710), .A2(G204gat), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n993), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g799(.A1(new_n1000), .A2(KEYINPUT62), .ZN(new_n1001));
  XNOR2_X1  g800(.A(new_n1001), .B(KEYINPUT125), .ZN(new_n1002));
  INV_X1    g801(.A(new_n949), .ZN(new_n1003));
  OAI21_X1  g802(.A(G204gat), .B1(new_n1003), .B2(new_n995), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1000), .A2(KEYINPUT62), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .ZN(G1353gat));
  INV_X1    g805(.A(G211gat), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n993), .A2(new_n1007), .A3(new_n639), .ZN(new_n1008));
  NOR4_X1   g807(.A1(new_n942), .A2(new_n948), .A3(new_n995), .A4(new_n907), .ZN(new_n1009));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n1010));
  AOI21_X1  g809(.A(new_n1007), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n891), .A2(new_n427), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1012), .A2(KEYINPUT57), .ZN(new_n1013));
  INV_X1    g812(.A(new_n948), .ZN(new_n1014));
  INV_X1    g813(.A(new_n995), .ZN(new_n1015));
  NAND4_X1  g814(.A1(new_n1013), .A2(new_n1014), .A3(new_n639), .A4(new_n1015), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1016), .A2(KEYINPUT126), .ZN(new_n1017));
  AOI21_X1  g816(.A(KEYINPUT63), .B1(new_n1011), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g817(.A(G211gat), .B1(new_n1016), .B2(KEYINPUT126), .ZN(new_n1019));
  AOI21_X1  g818(.A(new_n1010), .B1(new_n996), .B2(new_n639), .ZN(new_n1020));
  INV_X1    g819(.A(KEYINPUT63), .ZN(new_n1021));
  NOR3_X1   g820(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  OAI21_X1  g821(.A(new_n1008), .B1(new_n1018), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g822(.A(KEYINPUT127), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OAI211_X1 g824(.A(new_n1008), .B(KEYINPUT127), .C1(new_n1018), .C2(new_n1022), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n1025), .A2(new_n1026), .ZN(G1354gat));
  NOR3_X1   g826(.A1(new_n992), .A2(G218gat), .A3(new_n674), .ZN(new_n1028));
  INV_X1    g827(.A(G218gat), .ZN(new_n1029));
  AOI21_X1  g828(.A(new_n1029), .B1(new_n996), .B2(new_n798), .ZN(new_n1030));
  OR2_X1    g829(.A1(new_n1028), .A2(new_n1030), .ZN(G1355gat));
endmodule


