

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592;

  XNOR2_X1 U324 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U325 ( .A(n350), .B(n349), .ZN(n386) );
  XNOR2_X1 U326 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U327 ( .A(n340), .B(n339), .ZN(n342) );
  XNOR2_X1 U328 ( .A(KEYINPUT48), .B(KEYINPUT112), .ZN(n395) );
  XNOR2_X1 U329 ( .A(n396), .B(n395), .ZN(n547) );
  INV_X1 U330 ( .A(G169GAT), .ZN(n456) );
  XNOR2_X1 U331 ( .A(n456), .B(KEYINPUT122), .ZN(n457) );
  XNOR2_X1 U332 ( .A(n458), .B(n457), .ZN(G1348GAT) );
  XOR2_X1 U333 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n293) );
  NAND2_X1 U334 ( .A1(G229GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U335 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U336 ( .A(n294), .B(KEYINPUT69), .Z(n304) );
  XOR2_X1 U337 ( .A(G43GAT), .B(G29GAT), .Z(n296) );
  XNOR2_X1 U338 ( .A(KEYINPUT68), .B(G50GAT), .ZN(n295) );
  XNOR2_X1 U339 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U340 ( .A(n297), .B(KEYINPUT8), .Z(n299) );
  XNOR2_X1 U341 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n298) );
  XNOR2_X1 U342 ( .A(n299), .B(n298), .ZN(n382) );
  XOR2_X1 U343 ( .A(KEYINPUT67), .B(KEYINPUT70), .Z(n301) );
  XNOR2_X1 U344 ( .A(G197GAT), .B(KEYINPUT29), .ZN(n300) );
  XNOR2_X1 U345 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U346 ( .A(n382), .B(n302), .ZN(n303) );
  XNOR2_X1 U347 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U348 ( .A(G1GAT), .B(G8GAT), .Z(n365) );
  XNOR2_X1 U349 ( .A(n305), .B(n365), .ZN(n308) );
  XNOR2_X1 U350 ( .A(G169GAT), .B(G15GAT), .ZN(n306) );
  XNOR2_X1 U351 ( .A(n306), .B(G113GAT), .ZN(n326) );
  XOR2_X1 U352 ( .A(G141GAT), .B(G22GAT), .Z(n428) );
  XOR2_X1 U353 ( .A(n326), .B(n428), .Z(n307) );
  XNOR2_X1 U354 ( .A(n308), .B(n307), .ZN(n578) );
  INV_X1 U355 ( .A(n578), .ZN(n502) );
  XOR2_X1 U356 ( .A(n502), .B(KEYINPUT71), .Z(n530) );
  INV_X1 U357 ( .A(n530), .ZN(n455) );
  XOR2_X1 U358 ( .A(KEYINPUT87), .B(KEYINPUT64), .Z(n310) );
  XNOR2_X1 U359 ( .A(KEYINPUT86), .B(KEYINPUT90), .ZN(n309) );
  XNOR2_X1 U360 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U361 ( .A(KEYINPUT88), .B(n311), .Z(n313) );
  NAND2_X1 U362 ( .A1(G227GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U364 ( .A(n314), .B(KEYINPUT20), .Z(n319) );
  XOR2_X1 U365 ( .A(KEYINPUT89), .B(KEYINPUT17), .Z(n316) );
  XNOR2_X1 U366 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n315) );
  XNOR2_X1 U367 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U368 ( .A(KEYINPUT19), .B(n317), .Z(n413) );
  XNOR2_X1 U369 ( .A(n413), .B(KEYINPUT85), .ZN(n318) );
  XNOR2_X1 U370 ( .A(n319), .B(n318), .ZN(n324) );
  XNOR2_X1 U371 ( .A(G71GAT), .B(G176GAT), .ZN(n320) );
  XNOR2_X1 U372 ( .A(n320), .B(G120GAT), .ZN(n344) );
  XOR2_X1 U373 ( .A(G190GAT), .B(G134GAT), .Z(n375) );
  XOR2_X1 U374 ( .A(n344), .B(n375), .Z(n322) );
  XNOR2_X1 U375 ( .A(G43GAT), .B(G99GAT), .ZN(n321) );
  XNOR2_X1 U376 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U377 ( .A(n324), .B(n323), .Z(n328) );
  XNOR2_X1 U378 ( .A(G127GAT), .B(KEYINPUT0), .ZN(n325) );
  XNOR2_X1 U379 ( .A(n325), .B(KEYINPUT84), .ZN(n446) );
  XNOR2_X1 U380 ( .A(n326), .B(n446), .ZN(n327) );
  XOR2_X2 U381 ( .A(n328), .B(n327), .Z(n519) );
  INV_X1 U382 ( .A(n519), .ZN(n528) );
  XOR2_X1 U383 ( .A(G92GAT), .B(G85GAT), .Z(n330) );
  XNOR2_X1 U384 ( .A(G99GAT), .B(G106GAT), .ZN(n329) );
  XNOR2_X1 U385 ( .A(n330), .B(n329), .ZN(n373) );
  XNOR2_X1 U386 ( .A(n373), .B(KEYINPUT33), .ZN(n334) );
  INV_X1 U387 ( .A(n334), .ZN(n332) );
  AND2_X1 U388 ( .A1(G230GAT), .A2(G233GAT), .ZN(n333) );
  INV_X1 U389 ( .A(n333), .ZN(n331) );
  NAND2_X1 U390 ( .A1(n332), .A2(n331), .ZN(n336) );
  NAND2_X1 U391 ( .A1(n334), .A2(n333), .ZN(n335) );
  NAND2_X1 U392 ( .A1(n336), .A2(n335), .ZN(n340) );
  XOR2_X1 U393 ( .A(G148GAT), .B(G78GAT), .Z(n422) );
  XOR2_X1 U394 ( .A(n422), .B(KEYINPUT32), .Z(n338) );
  INV_X1 U395 ( .A(KEYINPUT31), .ZN(n337) );
  XNOR2_X1 U396 ( .A(G204GAT), .B(G64GAT), .ZN(n341) );
  XNOR2_X1 U397 ( .A(n341), .B(KEYINPUT73), .ZN(n406) );
  XNOR2_X1 U398 ( .A(n342), .B(n406), .ZN(n346) );
  XNOR2_X1 U399 ( .A(G57GAT), .B(KEYINPUT72), .ZN(n343) );
  XNOR2_X1 U400 ( .A(n343), .B(KEYINPUT13), .ZN(n366) );
  XOR2_X1 U401 ( .A(n344), .B(n366), .Z(n345) );
  XNOR2_X1 U402 ( .A(n346), .B(n345), .ZN(n390) );
  XOR2_X1 U403 ( .A(n390), .B(KEYINPUT41), .Z(n552) );
  OR2_X1 U404 ( .A1(n578), .A2(n552), .ZN(n350) );
  INV_X1 U405 ( .A(KEYINPUT111), .ZN(n348) );
  INV_X1 U406 ( .A(KEYINPUT46), .ZN(n347) );
  XOR2_X1 U407 ( .A(KEYINPUT81), .B(KEYINPUT12), .Z(n352) );
  XNOR2_X1 U408 ( .A(G64GAT), .B(KEYINPUT14), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n352), .B(n351), .ZN(n364) );
  XOR2_X1 U410 ( .A(G71GAT), .B(G127GAT), .Z(n354) );
  XNOR2_X1 U411 ( .A(G15GAT), .B(G183GAT), .ZN(n353) );
  XNOR2_X1 U412 ( .A(n354), .B(n353), .ZN(n362) );
  XOR2_X1 U413 ( .A(KEYINPUT15), .B(KEYINPUT79), .Z(n356) );
  XNOR2_X1 U414 ( .A(KEYINPUT78), .B(KEYINPUT80), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U416 ( .A(G78GAT), .B(G155GAT), .Z(n358) );
  XNOR2_X1 U417 ( .A(G22GAT), .B(G211GAT), .ZN(n357) );
  XNOR2_X1 U418 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U419 ( .A(n360), .B(n359), .Z(n361) );
  XNOR2_X1 U420 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n370) );
  XOR2_X1 U422 ( .A(n366), .B(n365), .Z(n368) );
  NAND2_X1 U423 ( .A1(G231GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U424 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U425 ( .A(n370), .B(n369), .Z(n585) );
  XOR2_X1 U426 ( .A(KEYINPUT75), .B(KEYINPUT10), .Z(n372) );
  XNOR2_X1 U427 ( .A(KEYINPUT9), .B(KEYINPUT11), .ZN(n371) );
  XNOR2_X1 U428 ( .A(n372), .B(n371), .ZN(n374) );
  XOR2_X1 U429 ( .A(n374), .B(n373), .Z(n377) );
  XOR2_X1 U430 ( .A(G218GAT), .B(G162GAT), .Z(n421) );
  XNOR2_X1 U431 ( .A(n375), .B(n421), .ZN(n376) );
  XNOR2_X1 U432 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U433 ( .A(KEYINPUT76), .B(KEYINPUT65), .Z(n379) );
  NAND2_X1 U434 ( .A1(G232GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U436 ( .A(n381), .B(n380), .Z(n384) );
  XNOR2_X1 U437 ( .A(n382), .B(KEYINPUT74), .ZN(n383) );
  XNOR2_X1 U438 ( .A(n384), .B(n383), .ZN(n559) );
  NAND2_X1 U439 ( .A1(n585), .A2(n559), .ZN(n385) );
  OR2_X1 U440 ( .A1(n386), .A2(n385), .ZN(n387) );
  XNOR2_X1 U441 ( .A(n387), .B(KEYINPUT47), .ZN(n394) );
  XOR2_X1 U442 ( .A(KEYINPUT77), .B(n559), .Z(n570) );
  XNOR2_X1 U443 ( .A(KEYINPUT36), .B(KEYINPUT100), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n570), .B(n388), .ZN(n589) );
  NOR2_X1 U445 ( .A1(n589), .A2(n585), .ZN(n389) );
  XNOR2_X1 U446 ( .A(KEYINPUT45), .B(n389), .ZN(n391) );
  NAND2_X1 U447 ( .A1(n391), .A2(n390), .ZN(n392) );
  NOR2_X1 U448 ( .A1(n530), .A2(n392), .ZN(n393) );
  NOR2_X1 U449 ( .A1(n394), .A2(n393), .ZN(n396) );
  XOR2_X1 U450 ( .A(KEYINPUT76), .B(G92GAT), .Z(n398) );
  XNOR2_X1 U451 ( .A(G36GAT), .B(G218GAT), .ZN(n397) );
  XNOR2_X1 U452 ( .A(n398), .B(n397), .ZN(n402) );
  XOR2_X1 U453 ( .A(G176GAT), .B(G190GAT), .Z(n400) );
  XNOR2_X1 U454 ( .A(G169GAT), .B(G8GAT), .ZN(n399) );
  XNOR2_X1 U455 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U456 ( .A(n402), .B(n401), .Z(n411) );
  XOR2_X1 U457 ( .A(KEYINPUT21), .B(KEYINPUT93), .Z(n404) );
  XNOR2_X1 U458 ( .A(KEYINPUT92), .B(G211GAT), .ZN(n403) );
  XNOR2_X1 U459 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U460 ( .A(G197GAT), .B(n405), .Z(n427) );
  XOR2_X1 U461 ( .A(n406), .B(KEYINPUT96), .Z(n408) );
  NAND2_X1 U462 ( .A1(G226GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U463 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U464 ( .A(n427), .B(n409), .ZN(n410) );
  XNOR2_X1 U465 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U466 ( .A(n413), .B(n412), .ZN(n517) );
  NOR2_X1 U467 ( .A1(n547), .A2(n517), .ZN(n414) );
  XNOR2_X1 U468 ( .A(n414), .B(KEYINPUT54), .ZN(n575) );
  XNOR2_X1 U469 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n415) );
  XNOR2_X1 U470 ( .A(n415), .B(KEYINPUT2), .ZN(n439) );
  XOR2_X1 U471 ( .A(n439), .B(KEYINPUT23), .Z(n420) );
  XOR2_X1 U472 ( .A(KEYINPUT24), .B(G204GAT), .Z(n417) );
  XNOR2_X1 U473 ( .A(G50GAT), .B(G106GAT), .ZN(n416) );
  XNOR2_X1 U474 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n418), .B(KEYINPUT22), .ZN(n419) );
  XNOR2_X1 U476 ( .A(n420), .B(n419), .ZN(n426) );
  XOR2_X1 U477 ( .A(n422), .B(n421), .Z(n424) );
  NAND2_X1 U478 ( .A1(G228GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U480 ( .A(n426), .B(n425), .Z(n430) );
  XNOR2_X1 U481 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U482 ( .A(n430), .B(n429), .ZN(n464) );
  XOR2_X1 U483 ( .A(KEYINPUT4), .B(G57GAT), .Z(n432) );
  XNOR2_X1 U484 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n431) );
  XNOR2_X1 U485 ( .A(n432), .B(n431), .ZN(n450) );
  XOR2_X1 U486 ( .A(G85GAT), .B(G120GAT), .Z(n434) );
  XNOR2_X1 U487 ( .A(G113GAT), .B(G134GAT), .ZN(n433) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U489 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n436) );
  XNOR2_X1 U490 ( .A(G141GAT), .B(G148GAT), .ZN(n435) );
  XNOR2_X1 U491 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U492 ( .A(n438), .B(n437), .Z(n444) );
  XOR2_X1 U493 ( .A(G162GAT), .B(n439), .Z(n441) );
  NAND2_X1 U494 ( .A1(G225GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U496 ( .A(G29GAT), .B(n442), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U498 ( .A(n445), .B(KEYINPUT6), .Z(n448) );
  XNOR2_X1 U499 ( .A(n446), .B(KEYINPUT1), .ZN(n447) );
  XNOR2_X1 U500 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U501 ( .A(n450), .B(n449), .Z(n459) );
  NOR2_X1 U502 ( .A1(n464), .A2(n459), .ZN(n451) );
  AND2_X1 U503 ( .A1(n575), .A2(n451), .ZN(n453) );
  XNOR2_X1 U504 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n452) );
  XNOR2_X1 U505 ( .A(n453), .B(n452), .ZN(n454) );
  NAND2_X1 U506 ( .A1(n528), .A2(n454), .ZN(n569) );
  NOR2_X1 U507 ( .A1(n455), .A2(n569), .ZN(n458) );
  INV_X1 U508 ( .A(n459), .ZN(n574) );
  AND2_X1 U509 ( .A1(n530), .A2(n390), .ZN(n490) );
  XOR2_X1 U510 ( .A(KEYINPUT91), .B(n519), .Z(n461) );
  XOR2_X1 U511 ( .A(KEYINPUT27), .B(n517), .Z(n467) );
  NAND2_X1 U512 ( .A1(n459), .A2(n467), .ZN(n546) );
  XOR2_X1 U513 ( .A(n464), .B(KEYINPUT28), .Z(n523) );
  INV_X1 U514 ( .A(n523), .ZN(n460) );
  NOR2_X1 U515 ( .A1(n546), .A2(n460), .ZN(n527) );
  NAND2_X1 U516 ( .A1(n461), .A2(n527), .ZN(n473) );
  NOR2_X1 U517 ( .A1(n519), .A2(n517), .ZN(n462) );
  NOR2_X1 U518 ( .A1(n464), .A2(n462), .ZN(n463) );
  XNOR2_X1 U519 ( .A(n463), .B(KEYINPUT25), .ZN(n469) );
  NAND2_X1 U520 ( .A1(n464), .A2(n519), .ZN(n466) );
  XNOR2_X1 U521 ( .A(KEYINPUT97), .B(KEYINPUT26), .ZN(n465) );
  XNOR2_X1 U522 ( .A(n466), .B(n465), .ZN(n576) );
  NAND2_X1 U523 ( .A1(n576), .A2(n467), .ZN(n468) );
  NAND2_X1 U524 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U525 ( .A(n470), .B(KEYINPUT98), .ZN(n471) );
  NAND2_X1 U526 ( .A1(n471), .A2(n574), .ZN(n472) );
  NAND2_X1 U527 ( .A1(n473), .A2(n472), .ZN(n486) );
  XOR2_X1 U528 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n475) );
  INV_X1 U529 ( .A(n585), .ZN(n537) );
  NAND2_X1 U530 ( .A1(n570), .A2(n537), .ZN(n474) );
  XNOR2_X1 U531 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U532 ( .A(KEYINPUT16), .B(n476), .Z(n477) );
  AND2_X1 U533 ( .A1(n486), .A2(n477), .ZN(n503) );
  NAND2_X1 U534 ( .A1(n490), .A2(n503), .ZN(n484) );
  NOR2_X1 U535 ( .A1(n574), .A2(n484), .ZN(n478) );
  XOR2_X1 U536 ( .A(KEYINPUT34), .B(n478), .Z(n479) );
  XNOR2_X1 U537 ( .A(G1GAT), .B(n479), .ZN(G1324GAT) );
  NOR2_X1 U538 ( .A1(n517), .A2(n484), .ZN(n480) );
  XOR2_X1 U539 ( .A(G8GAT), .B(n480), .Z(G1325GAT) );
  NOR2_X1 U540 ( .A1(n519), .A2(n484), .ZN(n482) );
  XNOR2_X1 U541 ( .A(KEYINPUT99), .B(KEYINPUT35), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U543 ( .A(G15GAT), .B(n483), .Z(G1326GAT) );
  NOR2_X1 U544 ( .A1(n523), .A2(n484), .ZN(n485) );
  XOR2_X1 U545 ( .A(G22GAT), .B(n485), .Z(G1327GAT) );
  NAND2_X1 U546 ( .A1(n585), .A2(n486), .ZN(n487) );
  NOR2_X1 U547 ( .A1(n589), .A2(n487), .ZN(n489) );
  XNOR2_X1 U548 ( .A(KEYINPUT37), .B(KEYINPUT101), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(n514) );
  NAND2_X1 U550 ( .A1(n490), .A2(n514), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n491), .B(KEYINPUT38), .ZN(n500) );
  NOR2_X1 U552 ( .A1(n500), .A2(n574), .ZN(n493) );
  XNOR2_X1 U553 ( .A(KEYINPUT102), .B(KEYINPUT39), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U555 ( .A(G29GAT), .B(n494), .ZN(G1328GAT) );
  NOR2_X1 U556 ( .A1(n500), .A2(n517), .ZN(n496) );
  XNOR2_X1 U557 ( .A(G36GAT), .B(KEYINPUT103), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(G1329GAT) );
  NOR2_X1 U559 ( .A1(n500), .A2(n519), .ZN(n498) );
  XNOR2_X1 U560 ( .A(KEYINPUT40), .B(KEYINPUT104), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U562 ( .A(G43GAT), .B(n499), .Z(G1330GAT) );
  NOR2_X1 U563 ( .A1(n523), .A2(n500), .ZN(n501) );
  XOR2_X1 U564 ( .A(G50GAT), .B(n501), .Z(G1331GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT105), .B(n552), .Z(n561) );
  NOR2_X1 U566 ( .A1(n502), .A2(n561), .ZN(n513) );
  NAND2_X1 U567 ( .A1(n513), .A2(n503), .ZN(n509) );
  NOR2_X1 U568 ( .A1(n574), .A2(n509), .ZN(n504) );
  XOR2_X1 U569 ( .A(G57GAT), .B(n504), .Z(n505) );
  XNOR2_X1 U570 ( .A(KEYINPUT42), .B(n505), .ZN(G1332GAT) );
  NOR2_X1 U571 ( .A1(n517), .A2(n509), .ZN(n506) );
  XOR2_X1 U572 ( .A(KEYINPUT106), .B(n506), .Z(n507) );
  XNOR2_X1 U573 ( .A(G64GAT), .B(n507), .ZN(G1333GAT) );
  NOR2_X1 U574 ( .A1(n519), .A2(n509), .ZN(n508) );
  XOR2_X1 U575 ( .A(G71GAT), .B(n508), .Z(G1334GAT) );
  NOR2_X1 U576 ( .A1(n523), .A2(n509), .ZN(n511) );
  XNOR2_X1 U577 ( .A(KEYINPUT43), .B(KEYINPUT107), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n511), .B(n510), .ZN(n512) );
  XOR2_X1 U579 ( .A(G78GAT), .B(n512), .Z(G1335GAT) );
  NAND2_X1 U580 ( .A1(n514), .A2(n513), .ZN(n522) );
  NOR2_X1 U581 ( .A1(n574), .A2(n522), .ZN(n515) );
  XOR2_X1 U582 ( .A(G85GAT), .B(n515), .Z(n516) );
  XNOR2_X1 U583 ( .A(KEYINPUT108), .B(n516), .ZN(G1336GAT) );
  NOR2_X1 U584 ( .A1(n517), .A2(n522), .ZN(n518) );
  XOR2_X1 U585 ( .A(G92GAT), .B(n518), .Z(G1337GAT) );
  NOR2_X1 U586 ( .A1(n519), .A2(n522), .ZN(n521) );
  XNOR2_X1 U587 ( .A(G99GAT), .B(KEYINPUT109), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(G1338GAT) );
  NOR2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n525) );
  XNOR2_X1 U590 ( .A(KEYINPUT110), .B(KEYINPUT44), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U592 ( .A(G106GAT), .B(n526), .Z(G1339GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n532) );
  NAND2_X1 U594 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U595 ( .A1(n547), .A2(n529), .ZN(n538) );
  NAND2_X1 U596 ( .A1(n538), .A2(n530), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U598 ( .A(G113GAT), .B(n533), .ZN(G1340GAT) );
  INV_X1 U599 ( .A(n538), .ZN(n542) );
  NOR2_X1 U600 ( .A1(n561), .A2(n542), .ZN(n535) );
  XNOR2_X1 U601 ( .A(KEYINPUT115), .B(KEYINPUT49), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U603 ( .A(G120GAT), .B(n536), .Z(G1341GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n540) );
  NAND2_X1 U605 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U607 ( .A(G127GAT), .B(n541), .Z(G1342GAT) );
  NOR2_X1 U608 ( .A1(n570), .A2(n542), .ZN(n544) );
  XNOR2_X1 U609 ( .A(KEYINPUT117), .B(KEYINPUT51), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U611 ( .A(G134GAT), .B(n545), .Z(G1343GAT) );
  NOR2_X1 U612 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U613 ( .A1(n548), .A2(n576), .ZN(n558) );
  NOR2_X1 U614 ( .A1(n578), .A2(n558), .ZN(n550) );
  XNOR2_X1 U615 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G141GAT), .B(n551), .ZN(G1344GAT) );
  NOR2_X1 U618 ( .A1(n552), .A2(n558), .ZN(n554) );
  XNOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(n555), .ZN(G1345GAT) );
  NOR2_X1 U622 ( .A1(n585), .A2(n558), .ZN(n556) );
  XOR2_X1 U623 ( .A(KEYINPUT120), .B(n556), .Z(n557) );
  XNOR2_X1 U624 ( .A(G155GAT), .B(n557), .ZN(G1346GAT) );
  NOR2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U626 ( .A(G162GAT), .B(n560), .Z(G1347GAT) );
  NOR2_X1 U627 ( .A1(n569), .A2(n561), .ZN(n563) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n565) );
  XOR2_X1 U630 ( .A(KEYINPUT56), .B(KEYINPUT123), .Z(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  INV_X1 U632 ( .A(KEYINPUT124), .ZN(n567) );
  NOR2_X1 U633 ( .A1(n585), .A2(n569), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(G183GAT), .B(n568), .ZN(G1350GAT) );
  INV_X1 U636 ( .A(KEYINPUT58), .ZN(n572) );
  NOR2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(G190GAT), .B(n573), .ZN(G1351GAT) );
  AND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n588) );
  NOR2_X1 U642 ( .A1(n588), .A2(n578), .ZN(n582) );
  XOR2_X1 U643 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n580) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  NOR2_X1 U647 ( .A1(n390), .A2(n588), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NOR2_X1 U650 ( .A1(n585), .A2(n588), .ZN(n586) );
  XOR2_X1 U651 ( .A(KEYINPUT126), .B(n586), .Z(n587) );
  XNOR2_X1 U652 ( .A(G211GAT), .B(n587), .ZN(G1354GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n591) );
  XNOR2_X1 U654 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

