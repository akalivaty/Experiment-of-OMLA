//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(KEYINPUT1), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n188), .A2(new_n190), .A3(new_n192), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n187), .A2(new_n189), .A3(G143), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n191), .B(G146), .C1(new_n187), .C2(KEYINPUT1), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n193), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT11), .ZN(new_n197));
  INV_X1    g011(.A(G134), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(G137), .ZN(new_n199));
  INV_X1    g013(.A(G137), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(KEYINPUT11), .A3(G134), .ZN(new_n201));
  INV_X1    g015(.A(G131), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(G137), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n199), .A2(new_n201), .A3(new_n202), .A4(new_n203), .ZN(new_n204));
  AND3_X1   g018(.A1(new_n200), .A2(KEYINPUT66), .A3(G134), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n200), .A2(G134), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT66), .B1(new_n200), .B2(G134), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n196), .B(new_n204), .C1(new_n208), .C2(new_n202), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT67), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(new_n206), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n200), .A2(KEYINPUT66), .A3(G134), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n202), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT67), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n214), .A2(new_n215), .A3(new_n196), .A4(new_n204), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n199), .A2(new_n203), .A3(new_n201), .ZN(new_n217));
  NAND2_X1  g031(.A1(KEYINPUT65), .A2(G131), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n199), .A2(new_n201), .A3(new_n218), .A4(new_n203), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(G143), .B(G146), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT0), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n223), .B1(new_n224), .B2(new_n187), .ZN(new_n225));
  XOR2_X1   g039(.A(KEYINPUT0), .B(G128), .Z(new_n226));
  OAI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(new_n223), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n222), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n210), .A2(new_n216), .A3(new_n228), .ZN(new_n229));
  XOR2_X1   g043(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  XOR2_X1   g045(.A(G116), .B(G119), .Z(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT2), .B(G113), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n232), .B(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n222), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n220), .A2(KEYINPUT68), .A3(new_n221), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(new_n227), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n239));
  INV_X1    g053(.A(new_n204), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n239), .B1(new_n213), .B2(new_n240), .ZN(new_n241));
  OAI211_X1 g055(.A(KEYINPUT69), .B(new_n204), .C1(new_n208), .C2(new_n202), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(new_n242), .A3(new_n196), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n238), .A2(KEYINPUT30), .A3(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n231), .A2(new_n234), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n234), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n238), .A2(new_n246), .A3(new_n243), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n238), .A2(new_n243), .A3(KEYINPUT70), .A4(new_n246), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n251), .B(G101), .ZN(new_n252));
  NOR2_X1   g066(.A1(G237), .A2(G953), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G210), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n252), .B(new_n254), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n245), .A2(new_n249), .A3(new_n250), .A4(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT31), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n249), .A2(new_n250), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT31), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n258), .A2(new_n259), .A3(new_n255), .A4(new_n245), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT28), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n247), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n229), .A2(new_n234), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n249), .A2(new_n250), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n263), .B1(new_n265), .B2(KEYINPUT28), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n257), .B(new_n260), .C1(new_n255), .C2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(G472), .A2(G902), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT32), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT32), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n267), .A2(new_n271), .A3(new_n268), .ZN(new_n272));
  INV_X1    g086(.A(new_n255), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT29), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n249), .A2(KEYINPUT71), .A3(new_n250), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT71), .B1(new_n249), .B2(new_n250), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n246), .B1(new_n238), .B2(new_n243), .ZN(new_n278));
  NOR3_X1   g092(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n262), .B(new_n275), .C1(new_n279), .C2(new_n261), .ZN(new_n280));
  XOR2_X1   g094(.A(KEYINPUT72), .B(G902), .Z(new_n281));
  NAND2_X1  g095(.A1(new_n266), .A2(new_n255), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n245), .A2(new_n249), .A3(new_n250), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT29), .B1(new_n283), .B2(new_n273), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n280), .A2(new_n285), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n270), .A2(new_n272), .B1(new_n286), .B2(G472), .ZN(new_n287));
  INV_X1    g101(.A(G217), .ZN(new_n288));
  INV_X1    g102(.A(new_n281), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n288), .B1(new_n289), .B2(G234), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(G902), .ZN(new_n291));
  XOR2_X1   g105(.A(G119), .B(G128), .Z(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT24), .B(G110), .ZN(new_n293));
  OR2_X1    g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G119), .ZN(new_n295));
  OR3_X1    g109(.A1(new_n295), .A2(KEYINPUT23), .A3(G128), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT23), .B1(new_n295), .B2(G128), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n296), .A2(new_n297), .B1(new_n295), .B2(G128), .ZN(new_n298));
  INV_X1    g112(.A(G110), .ZN(new_n299));
  OR2_X1    g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G140), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G125), .ZN(new_n302));
  INV_X1    g116(.A(G125), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G140), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n302), .A2(new_n304), .A3(KEYINPUT74), .A4(KEYINPUT16), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n302), .A2(new_n304), .A3(KEYINPUT16), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT16), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(new_n301), .A3(G125), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT74), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n189), .B(new_n305), .C1(new_n306), .C2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n302), .A2(new_n304), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n309), .B(new_n308), .C1(new_n313), .C2(new_n307), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n189), .B1(new_n314), .B2(new_n305), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n294), .B(new_n300), .C1(new_n312), .C2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n305), .B1(new_n306), .B2(new_n310), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G146), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n302), .A2(new_n304), .A3(new_n189), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n298), .A2(new_n299), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n292), .A2(new_n293), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n318), .B(new_n319), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT22), .B(G137), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n323), .B(KEYINPUT75), .ZN(new_n324));
  INV_X1    g138(.A(G953), .ZN(new_n325));
  AND3_X1   g139(.A1(new_n325), .A2(G221), .A3(G234), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n324), .B(new_n326), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n316), .A2(new_n322), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n327), .B1(new_n316), .B2(new_n322), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n330), .A2(KEYINPUT78), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n330), .A2(KEYINPUT78), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n291), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n316), .A2(new_n322), .ZN(new_n335));
  INV_X1    g149(.A(new_n327), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n316), .A2(new_n327), .A3(new_n322), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n289), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT76), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n334), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(KEYINPUT77), .B1(new_n330), .B2(new_n289), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT25), .ZN(new_n343));
  NOR3_X1   g157(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NOR3_X1   g158(.A1(new_n328), .A2(new_n329), .A3(new_n281), .ZN(new_n345));
  OAI211_X1 g159(.A(KEYINPUT77), .B(new_n343), .C1(new_n345), .C2(KEYINPUT76), .ZN(new_n346));
  XOR2_X1   g160(.A(new_n290), .B(KEYINPUT73), .Z(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n333), .B1(new_n344), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n287), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(G110), .B(G140), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n325), .A2(G227), .ZN(new_n353));
  XOR2_X1   g167(.A(new_n352), .B(new_n353), .Z(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G104), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT3), .B1(new_n356), .B2(G107), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT3), .ZN(new_n358));
  INV_X1    g172(.A(G107), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n359), .A3(G104), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n356), .A2(G107), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n357), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G101), .ZN(new_n363));
  INV_X1    g177(.A(G101), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n357), .A2(new_n360), .A3(new_n364), .A4(new_n361), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n363), .A2(KEYINPUT4), .A3(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT4), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n362), .A2(new_n367), .A3(G101), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n366), .A2(new_n368), .A3(new_n227), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n359), .A2(G104), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n356), .A2(G107), .ZN(new_n372));
  OAI21_X1  g186(.A(G101), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n365), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n370), .B1(new_n375), .B2(new_n196), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n193), .A2(new_n194), .A3(new_n195), .ZN(new_n377));
  NOR3_X1   g191(.A1(new_n377), .A2(new_n374), .A3(KEYINPUT10), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n369), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n236), .A2(new_n237), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n375), .A2(new_n370), .A3(new_n196), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n196), .A2(new_n373), .A3(new_n365), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT10), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n380), .B1(new_n386), .B2(new_n369), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n355), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n380), .A3(new_n369), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n377), .A2(new_n374), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n384), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n222), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT12), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT12), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n391), .A2(new_n394), .A3(new_n237), .A4(new_n236), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n389), .A2(new_n393), .A3(new_n395), .A4(new_n354), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n388), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G469), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n398), .A3(new_n289), .ZN(new_n399));
  INV_X1    g213(.A(G902), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n389), .A2(new_n393), .A3(new_n395), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n355), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n379), .A2(new_n381), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(new_n389), .A3(new_n354), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n399), .B(new_n402), .C1(new_n407), .C2(new_n398), .ZN(new_n408));
  INV_X1    g222(.A(G221), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT9), .B(G234), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n409), .B1(new_n411), .B2(new_n400), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(G116), .B(G119), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT5), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT5), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(new_n295), .A3(G116), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT79), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n417), .A2(new_n295), .A3(KEYINPUT79), .A4(G116), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n416), .A2(G113), .A3(new_n420), .A4(new_n421), .ZN(new_n422));
  OR2_X1    g236(.A1(new_n232), .A2(new_n233), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n374), .A2(KEYINPUT81), .ZN(new_n425));
  OR2_X1    g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(G110), .B(G122), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(KEYINPUT8), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n424), .A2(new_n425), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n234), .A2(new_n366), .A3(new_n368), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n375), .A2(new_n422), .A3(new_n423), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n432), .A3(new_n427), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n227), .A2(G125), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(G125), .B2(new_n377), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n325), .A2(G224), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT7), .ZN(new_n437));
  NAND2_X1  g251(.A1(KEYINPUT82), .A2(KEYINPUT7), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n435), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n437), .B1(new_n435), .B2(new_n438), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n430), .B(new_n433), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(KEYINPUT80), .A2(KEYINPUT6), .ZN(new_n442));
  AOI211_X1 g256(.A(new_n427), .B(new_n442), .C1(new_n431), .C2(new_n432), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n427), .B1(new_n431), .B2(new_n432), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n442), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n433), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n443), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  XOR2_X1   g262(.A(new_n435), .B(new_n436), .Z(new_n449));
  OAI211_X1 g263(.A(new_n400), .B(new_n441), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G210), .B1(G237), .B2(G902), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n435), .B(new_n436), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n444), .B1(new_n433), .B2(new_n446), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n454), .B1(new_n455), .B2(new_n443), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n456), .A2(new_n400), .A3(new_n451), .A4(new_n441), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(G214), .B1(G237), .B2(G902), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n414), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G237), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(new_n325), .A3(G214), .ZN(new_n463));
  NAND2_X1  g277(.A1(KEYINPUT83), .A2(G143), .ZN(new_n464));
  OR2_X1    g278(.A1(KEYINPUT83), .A2(G143), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(KEYINPUT83), .A2(G143), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n253), .A2(new_n467), .A3(G214), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n466), .A2(KEYINPUT17), .A3(G131), .A4(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n318), .A2(new_n311), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT88), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n466), .A2(G131), .A3(new_n468), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(G131), .B1(new_n466), .B2(new_n468), .ZN(new_n475));
  OR3_X1    g289(.A1(new_n474), .A2(KEYINPUT17), .A3(new_n475), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n318), .A2(KEYINPUT88), .A3(new_n311), .A4(new_n469), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n472), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT18), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT84), .B1(new_n479), .B2(new_n202), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT83), .B(G143), .ZN(new_n481));
  INV_X1    g295(.A(G214), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n482), .A2(G237), .A3(G953), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n480), .B(new_n468), .C1(new_n481), .C2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n479), .A2(new_n202), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT84), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n313), .A2(G146), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n319), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n466), .A2(new_n486), .A3(new_n485), .A4(new_n468), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n488), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT85), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT85), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n488), .A2(new_n494), .A3(new_n490), .A4(new_n491), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  XOR2_X1   g310(.A(G113), .B(G122), .Z(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(KEYINPUT87), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n498), .B(new_n356), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n478), .A2(new_n496), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(KEYINPUT86), .B1(new_n474), .B2(new_n475), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n466), .A2(new_n468), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n202), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT86), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(new_n505), .A3(new_n473), .ZN(new_n506));
  OR2_X1    g320(.A1(new_n313), .A2(KEYINPUT19), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n313), .A2(KEYINPUT19), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n189), .A3(new_n508), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n502), .A2(new_n506), .A3(new_n318), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n496), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n499), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n501), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(G475), .A2(G902), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT20), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT20), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n513), .A2(new_n517), .A3(new_n514), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n513), .A2(KEYINPUT89), .A3(new_n517), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n516), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(G128), .B(G143), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n198), .ZN(new_n522));
  INV_X1    g336(.A(G122), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G116), .ZN(new_n524));
  INV_X1    g338(.A(G116), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G122), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n524), .A2(new_n526), .A3(new_n359), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n359), .B1(new_n524), .B2(new_n526), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n522), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n191), .A2(G128), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n187), .A2(G143), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n531), .A3(KEYINPUT13), .ZN(new_n532));
  OR3_X1    g346(.A1(new_n187), .A2(KEYINPUT13), .A3(G143), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n532), .A2(G134), .A3(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT90), .B1(new_n529), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n528), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n524), .A2(new_n526), .A3(new_n359), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n532), .A2(new_n533), .A3(G134), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT90), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n538), .A2(new_n539), .A3(new_n540), .A4(new_n522), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n521), .B(new_n198), .ZN(new_n543));
  OR2_X1    g357(.A1(new_n526), .A2(KEYINPUT14), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT14), .B1(new_n523), .B2(G116), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT91), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT91), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n526), .A2(new_n547), .A3(KEYINPUT14), .ZN(new_n548));
  AND4_X1   g362(.A1(new_n524), .A2(new_n544), .A3(new_n546), .A4(new_n548), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n537), .B(new_n543), .C1(new_n549), .C2(new_n359), .ZN(new_n550));
  NOR3_X1   g364(.A1(new_n410), .A2(new_n288), .A3(G953), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n542), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n551), .B1(new_n542), .B2(new_n550), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n289), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT92), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(G478), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n557), .A2(KEYINPUT15), .ZN(new_n558));
  OAI211_X1 g372(.A(KEYINPUT92), .B(new_n289), .C1(new_n552), .C2(new_n553), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n556), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  OR2_X1    g374(.A1(new_n554), .A2(new_n558), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n478), .A2(new_n496), .A3(new_n500), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n500), .B1(new_n478), .B2(new_n496), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n400), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G475), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n513), .A2(KEYINPUT89), .A3(new_n517), .A4(new_n514), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n520), .A2(new_n562), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n325), .A2(G952), .ZN(new_n570));
  NAND2_X1  g384(.A1(G234), .A2(G237), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n281), .A2(G953), .A3(new_n571), .ZN(new_n574));
  XOR2_X1   g388(.A(new_n574), .B(KEYINPUT93), .Z(new_n575));
  XNOR2_X1  g389(.A(KEYINPUT21), .B(G898), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n573), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n461), .A2(new_n569), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n351), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(G101), .ZN(G3));
  INV_X1    g396(.A(G472), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n267), .B2(new_n289), .ZN(new_n584));
  INV_X1    g398(.A(new_n268), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n257), .A2(new_n260), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n265), .A2(KEYINPUT28), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n255), .B1(new_n587), .B2(new_n262), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n585), .B1(new_n586), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n414), .ZN(new_n592));
  INV_X1    g406(.A(new_n350), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT94), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT94), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n591), .A2(new_n596), .A3(new_n592), .A4(new_n593), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g412(.A(new_n598), .B(KEYINPUT95), .Z(new_n599));
  NAND3_X1  g413(.A1(new_n520), .A2(new_n566), .A3(new_n567), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n601));
  OAI21_X1  g415(.A(KEYINPUT33), .B1(new_n551), .B2(KEYINPUT96), .ZN(new_n602));
  OR3_X1    g416(.A1(new_n552), .A2(new_n553), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n602), .B1(new_n552), .B2(new_n553), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n603), .A2(G478), .A3(new_n289), .A4(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n600), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n459), .ZN(new_n609));
  AOI211_X1 g423(.A(new_n609), .B(new_n577), .C1(new_n453), .C2(new_n457), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n599), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT34), .B(G104), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  AOI21_X1  g427(.A(new_n517), .B1(new_n513), .B2(new_n514), .ZN(new_n614));
  INV_X1    g428(.A(new_n514), .ZN(new_n615));
  AOI211_X1 g429(.A(KEYINPUT20), .B(new_n615), .C1(new_n501), .C2(new_n512), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n566), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(new_n562), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n599), .A2(new_n610), .A3(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT35), .B(G107), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT97), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n619), .B(new_n621), .ZN(G9));
  NAND2_X1  g436(.A1(new_n257), .A2(new_n260), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n289), .B1(new_n623), .B2(new_n588), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(G472), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n269), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n579), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n336), .A2(KEYINPUT36), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(new_n335), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n291), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n630), .B1(new_n344), .B2(new_n349), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G110), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT98), .B(KEYINPUT37), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G12));
  AOI21_X1  g449(.A(new_n609), .B1(new_n453), .B2(new_n457), .ZN(new_n636));
  INV_X1    g450(.A(G900), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n575), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n572), .B(KEYINPUT99), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n618), .A2(KEYINPUT100), .A3(new_n636), .A4(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT100), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n516), .A2(new_n518), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n560), .A2(new_n561), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n644), .A2(new_n645), .A3(new_n566), .A4(new_n641), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n643), .B1(new_n646), .B2(new_n460), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n414), .B1(new_n642), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g462(.A(KEYINPUT77), .B1(new_n345), .B2(KEYINPUT76), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n339), .A2(new_n334), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n649), .A2(KEYINPUT25), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n347), .B1(new_n341), .B2(new_n343), .ZN(new_n652));
  AOI22_X1  g466(.A1(new_n651), .A2(new_n652), .B1(new_n291), .B2(new_n629), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n270), .A2(new_n272), .ZN(new_n654));
  INV_X1    g468(.A(new_n275), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n249), .A2(new_n250), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT71), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n278), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n249), .A2(KEYINPUT71), .A3(new_n250), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  AOI211_X1 g475(.A(new_n263), .B(new_n655), .C1(new_n661), .C2(KEYINPUT28), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n283), .A2(new_n273), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n274), .ZN(new_n664));
  AOI211_X1 g478(.A(new_n273), .B(new_n263), .C1(new_n265), .C2(KEYINPUT28), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n289), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(G472), .B1(new_n662), .B2(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n653), .B1(new_n654), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n648), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G128), .ZN(G30));
  AOI21_X1  g484(.A(new_n271), .B1(new_n267), .B2(new_n268), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n267), .A2(new_n271), .A3(new_n268), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n283), .A2(new_n255), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  AOI211_X1 g488(.A(G902), .B(new_n674), .C1(new_n279), .C2(new_n273), .ZN(new_n675));
  OAI22_X1  g489(.A1(new_n671), .A2(new_n672), .B1(new_n675), .B2(new_n583), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT101), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n562), .A2(new_n609), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n678), .A2(new_n600), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n640), .B(KEYINPUT39), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n414), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT40), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n631), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n458), .B(KEYINPUT38), .ZN(new_n685));
  OAI21_X1  g499(.A(KEYINPUT40), .B1(new_n414), .B2(new_n681), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n680), .A2(new_n684), .A3(new_n685), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G143), .ZN(G45));
  OAI21_X1  g502(.A(new_n667), .B1(new_n671), .B2(new_n672), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n600), .A2(new_n606), .A3(new_n641), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n689), .A2(new_n690), .A3(new_n461), .A4(new_n631), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  AND4_X1   g506(.A1(new_n389), .A2(new_n393), .A3(new_n395), .A4(new_n354), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n354), .B1(new_n405), .B2(new_n389), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n289), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(G469), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n696), .A2(new_n697), .A3(new_n399), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n695), .A2(KEYINPUT102), .A3(G469), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n412), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AND4_X1   g514(.A1(new_n600), .A2(new_n700), .A3(new_n610), .A4(new_n606), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(new_n593), .A3(new_n689), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT103), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT41), .B(G113), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G15));
  OAI211_X1 g519(.A(new_n645), .B(new_n566), .C1(new_n614), .C2(new_n616), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n350), .A2(new_n706), .A3(new_n577), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n698), .A2(new_n699), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n708), .A2(new_n636), .A3(new_n413), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n672), .A2(new_n671), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n583), .B1(new_n280), .B2(new_n285), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n707), .B(new_n709), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G116), .ZN(G18));
  NOR3_X1   g527(.A1(new_n568), .A2(new_n577), .A3(new_n653), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n689), .A2(new_n714), .A3(new_n709), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G119), .ZN(G21));
  AND3_X1   g530(.A1(new_n600), .A2(new_n458), .A3(new_n679), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n263), .B1(new_n661), .B2(KEYINPUT28), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n586), .B1(new_n718), .B2(new_n255), .ZN(new_n719));
  XOR2_X1   g533(.A(new_n268), .B(KEYINPUT104), .Z(new_n720));
  AOI22_X1  g534(.A1(new_n719), .A2(new_n720), .B1(new_n624), .B2(G472), .ZN(new_n721));
  AOI211_X1 g535(.A(new_n412), .B(new_n577), .C1(new_n698), .C2(new_n699), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n717), .A2(new_n593), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G122), .ZN(G24));
  INV_X1    g538(.A(KEYINPUT105), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n690), .A2(new_n709), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n262), .B1(new_n279), .B2(new_n261), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n623), .B1(new_n727), .B2(new_n273), .ZN(new_n728));
  INV_X1    g542(.A(new_n720), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n625), .B(new_n631), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n725), .B1(new_n726), .B2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n730), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n600), .A2(new_n606), .A3(new_n641), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n708), .A2(new_n636), .A3(new_n413), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n732), .A2(new_n735), .A3(KEYINPUT105), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G125), .ZN(G27));
  INV_X1    g552(.A(KEYINPUT42), .ZN(new_n739));
  INV_X1    g553(.A(new_n399), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n401), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n404), .A2(KEYINPUT106), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT106), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n403), .A2(new_n743), .A3(new_n355), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n742), .A2(new_n406), .A3(new_n744), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n745), .A2(new_n398), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n412), .B1(new_n741), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n689), .A2(new_n593), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n453), .A2(new_n459), .A3(new_n457), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n690), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n739), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n733), .A2(new_n749), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n351), .A2(new_n753), .A3(KEYINPUT42), .A4(new_n747), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G131), .ZN(G33));
  OR3_X1    g570(.A1(new_n748), .A2(new_n646), .A3(new_n749), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G134), .ZN(G36));
  NAND4_X1  g572(.A1(new_n520), .A2(new_n606), .A3(new_n566), .A4(new_n567), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT43), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n759), .B(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT107), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n762), .B1(new_n626), .B2(new_n631), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n762), .B(new_n631), .C1(new_n584), .C2(new_n590), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n761), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT44), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n407), .A2(new_n769), .ZN(new_n770));
  OAI211_X1 g584(.A(G469), .B(new_n770), .C1(new_n745), .C2(new_n769), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT46), .B1(new_n771), .B2(new_n402), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n740), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n771), .A2(KEYINPUT46), .A3(new_n402), .ZN(new_n774));
  AOI211_X1 g588(.A(new_n412), .B(new_n681), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n761), .B(KEYINPUT44), .C1(new_n763), .C2(new_n765), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n768), .A2(new_n750), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G137), .ZN(G39));
  NOR2_X1   g592(.A1(new_n689), .A2(new_n593), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n412), .B1(new_n773), .B2(new_n774), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n780), .A2(KEYINPUT47), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n780), .A2(KEYINPUT47), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n753), .B(new_n779), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G140), .ZN(G42));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n785));
  INV_X1    g599(.A(new_n617), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n689), .A2(new_n592), .A3(new_n562), .A4(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n608), .A2(new_n721), .A3(new_n747), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n653), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n749), .A2(new_n640), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT110), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n734), .B1(new_n654), .B2(new_n667), .ZN(new_n793));
  AOI22_X1  g607(.A1(new_n351), .A2(new_n701), .B1(new_n793), .B2(new_n714), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n723), .A2(new_n712), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n792), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n702), .A2(new_n715), .A3(new_n723), .A4(new_n712), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(KEYINPUT110), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n791), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  AOI22_X1  g613(.A1(new_n627), .A2(new_n631), .B1(new_n351), .B2(new_n580), .ZN(new_n800));
  OR3_X1    g614(.A1(new_n600), .A2(KEYINPUT111), .A3(new_n562), .ZN(new_n801));
  OAI21_X1  g615(.A(KEYINPUT111), .B1(new_n600), .B2(new_n562), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(new_n607), .A3(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(new_n595), .A3(new_n610), .A4(new_n597), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n755), .A2(new_n757), .A3(new_n800), .A4(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n785), .B1(new_n799), .B2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT105), .B1(new_n732), .B2(new_n735), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n730), .A2(new_n733), .A3(new_n725), .A4(new_n734), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n669), .B(new_n691), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n676), .A2(new_n717), .A3(new_n653), .A4(new_n641), .ZN(new_n811));
  INV_X1    g625(.A(new_n747), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n807), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n813), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n592), .A2(new_n636), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n287), .A2(new_n816), .A3(new_n653), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n817), .A2(new_n690), .B1(new_n648), .B2(new_n668), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n815), .A2(new_n737), .A3(new_n818), .A4(KEYINPUT52), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n794), .A2(new_n795), .A3(new_n792), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n797), .A2(KEYINPUT110), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n821), .A2(new_n822), .B1(new_n789), .B2(new_n790), .ZN(new_n823));
  AND4_X1   g637(.A1(new_n755), .A2(new_n757), .A3(new_n800), .A4(new_n804), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n824), .A3(KEYINPUT112), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n806), .A2(new_n820), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n806), .A2(new_n825), .A3(KEYINPUT53), .A4(new_n820), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT54), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n678), .A2(new_n350), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n700), .A2(new_n750), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT115), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n832), .A2(new_n573), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n608), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n761), .A2(new_n639), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n351), .A3(new_n834), .ZN(new_n838));
  NAND2_X1  g652(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n570), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OR2_X1    g654(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n838), .A2(new_n839), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n600), .ZN(new_n844));
  INV_X1    g658(.A(new_n606), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n835), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n781), .A2(new_n782), .ZN(new_n847));
  INV_X1    g661(.A(new_n708), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n847), .B1(new_n413), .B2(new_n848), .ZN(new_n849));
  AND4_X1   g663(.A1(new_n593), .A2(new_n761), .A3(new_n639), .A4(new_n721), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n849), .A2(new_n750), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n837), .A2(new_n732), .A3(new_n834), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n846), .A2(new_n851), .A3(KEYINPUT51), .A4(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT113), .ZN(new_n854));
  INV_X1    g668(.A(new_n685), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n850), .A2(new_n855), .A3(new_n700), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n854), .B1(new_n856), .B2(new_n459), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT50), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n854), .B(KEYINPUT50), .C1(new_n856), .C2(new_n459), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n836), .B(new_n843), .C1(new_n853), .C2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT51), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n846), .A2(new_n851), .A3(new_n852), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n861), .A2(KEYINPUT114), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT114), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n859), .A2(new_n866), .A3(new_n860), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n864), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n862), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n797), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n827), .B1(new_n789), .B2(new_n790), .ZN(new_n871));
  AND4_X1   g685(.A1(new_n820), .A2(new_n870), .A3(new_n824), .A4(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n826), .B2(new_n827), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n850), .A2(new_n709), .ZN(new_n876));
  AND4_X1   g690(.A1(new_n831), .A2(new_n869), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(G952), .A2(G953), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n350), .A2(new_n609), .A3(new_n412), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT108), .ZN(new_n880));
  OR4_X1    g694(.A1(new_n685), .A2(new_n678), .A3(new_n759), .A4(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n848), .B1(KEYINPUT109), .B2(KEYINPUT49), .ZN(new_n882));
  NOR2_X1   g696(.A1(KEYINPUT109), .A2(KEYINPUT49), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n882), .B(new_n883), .ZN(new_n884));
  OAI22_X1  g698(.A1(new_n877), .A2(new_n878), .B1(new_n881), .B2(new_n884), .ZN(G75));
  NOR2_X1   g699(.A1(new_n325), .A2(G952), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT117), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT56), .ZN(new_n888));
  INV_X1    g702(.A(new_n872), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n828), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n281), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n888), .B1(new_n891), .B2(new_n451), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n448), .B(new_n454), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT55), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n894), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n888), .B(new_n896), .C1(new_n891), .C2(new_n451), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n887), .B1(new_n895), .B2(new_n897), .ZN(G51));
  XNOR2_X1  g712(.A(new_n401), .B(KEYINPUT57), .ZN(new_n899));
  AOI211_X1 g713(.A(KEYINPUT54), .B(new_n872), .C1(new_n827), .C2(new_n826), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n874), .B1(new_n828), .B2(new_n889), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n397), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n891), .A2(new_n771), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n886), .B1(new_n903), .B2(new_n904), .ZN(G54));
  NOR2_X1   g719(.A1(new_n873), .A2(new_n289), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(KEYINPUT58), .A3(G475), .ZN(new_n907));
  INV_X1    g721(.A(new_n513), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n886), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n906), .A2(KEYINPUT58), .A3(G475), .A4(new_n513), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(G60));
  INV_X1    g726(.A(new_n887), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n603), .A2(new_n604), .ZN(new_n914));
  NAND2_X1  g728(.A1(G478), .A2(G902), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT59), .Z(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n914), .B(new_n917), .C1(new_n900), .C2(new_n901), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n916), .B1(new_n831), .B2(new_n875), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n913), .B(new_n918), .C1(new_n919), .C2(new_n914), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(G63));
  XNOR2_X1  g735(.A(KEYINPUT118), .B(KEYINPUT60), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n288), .A2(new_n400), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n922), .B(new_n923), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n629), .B(KEYINPUT119), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n890), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n331), .A2(new_n332), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n924), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n928), .B1(new_n873), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n926), .A2(new_n930), .A3(new_n913), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n926), .A2(new_n930), .A3(KEYINPUT61), .A4(new_n913), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(G66));
  NAND2_X1  g749(.A1(new_n821), .A2(new_n822), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n800), .A2(new_n804), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n939), .A2(KEYINPUT120), .A3(G953), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n939), .A2(G953), .ZN(new_n942));
  INV_X1    g756(.A(G224), .ZN(new_n943));
  OAI21_X1  g757(.A(G953), .B1(new_n576), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT120), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n941), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n448), .B1(G898), .B2(new_n325), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n946), .B(new_n947), .Z(G69));
  AOI21_X1  g762(.A(new_n325), .B1(G227), .B2(G900), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(KEYINPUT126), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n949), .A2(KEYINPUT126), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n231), .A2(new_n244), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT121), .Z(new_n953));
  NAND2_X1  g767(.A1(new_n507), .A2(new_n508), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n955), .B1(G900), .B2(G953), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n808), .A2(new_n809), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n669), .A2(new_n691), .ZN(new_n959));
  OAI21_X1  g773(.A(KEYINPUT122), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT122), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n737), .A2(new_n818), .A3(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n960), .A2(new_n777), .A3(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT124), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n960), .A2(new_n777), .A3(new_n962), .A4(KEYINPUT124), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n775), .A2(new_n351), .A3(new_n717), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n783), .A2(new_n755), .A3(new_n968), .A4(new_n757), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(KEYINPUT125), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT125), .ZN(new_n972));
  AOI211_X1 g786(.A(new_n972), .B(new_n969), .C1(new_n965), .C2(new_n966), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n957), .B1(new_n974), .B2(new_n325), .ZN(new_n975));
  INV_X1    g789(.A(new_n955), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n687), .A2(new_n960), .A3(new_n962), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n977), .B1(KEYINPUT123), .B2(KEYINPUT62), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n803), .A2(new_n351), .A3(new_n682), .A4(new_n750), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n777), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g794(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n687), .A2(new_n960), .A3(new_n962), .A4(new_n981), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n978), .A2(new_n783), .A3(new_n980), .A4(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n976), .B1(new_n983), .B2(new_n325), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n950), .B(new_n951), .C1(new_n975), .C2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n967), .A2(new_n970), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(new_n972), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n967), .A2(KEYINPUT125), .A3(new_n970), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n987), .A2(new_n325), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n956), .ZN(new_n990));
  INV_X1    g804(.A(new_n984), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n990), .A2(new_n991), .A3(KEYINPUT126), .A4(new_n949), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n985), .A2(new_n992), .ZN(G72));
  NOR2_X1   g807(.A1(new_n283), .A2(new_n255), .ZN(new_n994));
  NOR3_X1   g808(.A1(new_n971), .A2(new_n973), .A3(new_n938), .ZN(new_n995));
  NAND2_X1  g809(.A1(G472), .A2(G902), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n996), .B(KEYINPUT63), .Z(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n994), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n997), .B1(new_n983), .B2(new_n938), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n886), .B1(new_n1000), .B2(new_n674), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n674), .B1(new_n828), .B2(new_n829), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT127), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n994), .A2(new_n998), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1003), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n999), .B(new_n1001), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(G57));
endmodule


