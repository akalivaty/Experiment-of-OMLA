//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n769, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n988,
    new_n989;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n202));
  INV_X1    g001(.A(G226gat), .ZN(new_n203));
  INV_X1    g002(.A(G233gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G183gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT27), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT27), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G183gat), .ZN(new_n209));
  INV_X1    g008(.A(G190gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n207), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT28), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT27), .B(G183gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(KEYINPUT28), .A3(new_n210), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  INV_X1    g016(.A(G169gat), .ZN(new_n218));
  INV_X1    g017(.A(G176gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT69), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT26), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n220), .B1(KEYINPUT67), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT26), .B1(new_n224), .B2(new_n221), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n217), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n216), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n206), .A2(new_n210), .ZN(new_n229));
  NAND3_X1  g028(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT68), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT24), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n232), .B1(new_n227), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n227), .A2(new_n232), .A3(new_n233), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n231), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT23), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n220), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT23), .ZN(new_n240));
  NOR3_X1   g039(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n239), .B(new_n217), .C1(new_n240), .C2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT25), .B1(new_n237), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT25), .ZN(new_n244));
  NOR2_X1   g043(.A1(G169gat), .A2(G176gat), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n244), .B(new_n217), .C1(new_n245), .C2(KEYINPUT23), .ZN(new_n246));
  XOR2_X1   g045(.A(KEYINPUT66), .B(G176gat), .Z(new_n247));
  NOR2_X1   g046(.A1(new_n238), .A2(G169gat), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(G183gat), .A2(G190gat), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n250), .B1(new_n233), .B2(new_n227), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n230), .A2(KEYINPUT65), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n230), .A2(KEYINPUT65), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n228), .A2(new_n243), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT29), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n205), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n205), .ZN(new_n259));
  AND2_X1   g058(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n250), .B1(new_n260), .B2(G190gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n236), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n261), .B1(new_n262), .B2(new_n234), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n239), .A2(new_n217), .ZN(new_n264));
  INV_X1    g063(.A(new_n241), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n265), .A2(KEYINPUT23), .A3(new_n224), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n263), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n267), .A2(KEYINPUT25), .B1(new_n254), .B2(new_n249), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n259), .B1(new_n268), .B2(new_n228), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n258), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G211gat), .B(G218gat), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(G218gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT75), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT75), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(G218gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT22), .B1(new_n277), .B2(G211gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(G197gat), .B(G204gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n272), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G211gat), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n282), .B1(new_n274), .B2(new_n276), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n271), .B(new_n279), .C1(new_n283), .C2(KEYINPUT22), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n281), .A2(KEYINPUT76), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT22), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT75), .B(G218gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n286), .B1(new_n287), .B2(new_n282), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n271), .B1(new_n288), .B2(new_n279), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT76), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT77), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n285), .A2(KEYINPUT77), .A3(new_n291), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n270), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT78), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n295), .B(new_n294), .C1(new_n258), .C2(new_n269), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n295), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT77), .B1(new_n285), .B2(new_n291), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n303), .B(KEYINPUT78), .C1(new_n258), .C2(new_n269), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G8gat), .B(G36gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n306), .B(G64gat), .ZN(new_n307));
  INV_X1    g106(.A(G92gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT30), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n305), .A2(KEYINPUT30), .A3(new_n309), .ZN(new_n313));
  OR2_X1    g112(.A1(new_n305), .A2(new_n309), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT5), .ZN(new_n316));
  OR2_X1    g115(.A1(G141gat), .A2(G148gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(G141gat), .A2(G148gat), .ZN(new_n318));
  AND2_X1   g117(.A1(G155gat), .A2(G162gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT2), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n317), .B(new_n318), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT80), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT79), .ZN(new_n323));
  INV_X1    g122(.A(G155gat), .ZN(new_n324));
  INV_X1    g123(.A(G162gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT79), .B1(G155gat), .B2(G162gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n319), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n322), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AOI211_X1 g129(.A(KEYINPUT80), .B(new_n319), .C1(new_n326), .C2(new_n327), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n321), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n318), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT81), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT81), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n317), .A2(new_n335), .A3(new_n318), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n324), .A3(new_n325), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n329), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n334), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n332), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(G113gat), .ZN(new_n341));
  INV_X1    g140(.A(G120gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT1), .ZN(new_n344));
  NAND2_X1  g143(.A1(G113gat), .A2(G120gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(G134gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(G127gat), .ZN(new_n348));
  INV_X1    g147(.A(G127gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G134gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT1), .B1(new_n341), .B2(new_n342), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n353), .A2(new_n345), .B1(new_n348), .B2(new_n350), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n340), .B(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(G225gat), .A2(G233gat), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n316), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n340), .A2(KEYINPUT3), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT3), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n332), .A2(new_n362), .A3(new_n339), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n361), .A2(new_n363), .A3(new_n356), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n365));
  OAI22_X1  g164(.A1(new_n340), .A2(new_n356), .B1(new_n365), .B2(new_n359), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT70), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n367), .B1(new_n352), .B2(new_n354), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n346), .A2(new_n351), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n353), .A2(new_n345), .A3(new_n348), .A4(new_n350), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT70), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n332), .A2(new_n339), .A3(new_n368), .A4(new_n371), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n364), .B(new_n366), .C1(new_n365), .C2(new_n372), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n360), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n359), .A2(KEYINPUT5), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n372), .A2(new_n365), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n332), .A2(KEYINPUT4), .A3(new_n339), .A4(new_n355), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n376), .A2(KEYINPUT83), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT83), .B1(new_n376), .B2(new_n377), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n364), .B(new_n375), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT84), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT83), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n334), .A2(new_n336), .A3(new_n338), .ZN(new_n383));
  INV_X1    g182(.A(new_n327), .ZN(new_n384));
  NOR3_X1   g183(.A1(KEYINPUT79), .A2(G155gat), .A3(G162gat), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n329), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT80), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n328), .A2(new_n322), .A3(new_n329), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n383), .B1(new_n389), .B2(new_n321), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n352), .A2(new_n354), .A3(new_n367), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT70), .B1(new_n369), .B2(new_n370), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT4), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n377), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n382), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n376), .A2(KEYINPUT83), .A3(new_n377), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT84), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n398), .A2(new_n399), .A3(new_n364), .A4(new_n375), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n374), .B1(new_n381), .B2(new_n400), .ZN(new_n401));
  XOR2_X1   g200(.A(G57gat), .B(G85gat), .Z(new_n402));
  XNOR2_X1  g201(.A(G1gat), .B(G29gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n404), .B(new_n405), .Z(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT6), .B1(new_n401), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n374), .ZN(new_n409));
  INV_X1    g208(.A(new_n400), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n361), .A2(new_n363), .A3(new_n356), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n411), .B1(new_n396), .B2(new_n397), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n399), .B1(new_n412), .B2(new_n375), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n409), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n406), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n408), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n414), .A2(KEYINPUT6), .A3(new_n406), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n315), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT89), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n256), .A2(new_n393), .ZN(new_n420));
  NAND2_X1  g219(.A1(G227gat), .A2(G233gat), .ZN(new_n421));
  XOR2_X1   g220(.A(new_n421), .B(KEYINPUT64), .Z(new_n422));
  NAND2_X1  g221(.A1(new_n368), .A2(new_n371), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n423), .A2(new_n228), .A3(new_n243), .A4(new_n255), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n420), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT33), .ZN(new_n426));
  INV_X1    g225(.A(G99gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(G15gat), .B(G43gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n428), .B(KEYINPUT71), .ZN(new_n429));
  INV_X1    g228(.A(G71gat), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT71), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n428), .B(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n433), .A2(G71gat), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n427), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(G71gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n429), .A2(new_n430), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(new_n437), .A3(G99gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n425), .B(KEYINPUT32), .C1(new_n426), .C2(new_n439), .ZN(new_n440));
  OR2_X1    g239(.A1(new_n426), .A2(KEYINPUT32), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n439), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT72), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT72), .ZN(new_n445));
  AOI211_X1 g244(.A(new_n445), .B(new_n439), .C1(new_n425), .C2(new_n441), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n440), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n422), .ZN(new_n448));
  INV_X1    g247(.A(new_n424), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n423), .B1(new_n268), .B2(new_n228), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n452), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n448), .B(new_n454), .C1(new_n449), .C2(new_n450), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n447), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT74), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT74), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n447), .A2(new_n460), .A3(new_n457), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(G22gat), .B(G50gat), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n363), .A2(new_n257), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n294), .A2(new_n295), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n284), .ZN(new_n467));
  OAI211_X1 g266(.A(KEYINPUT85), .B(new_n257), .C1(new_n467), .C2(new_n289), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n362), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n281), .A2(new_n284), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT85), .B1(new_n470), .B2(new_n257), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n340), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(G228gat), .A2(G233gat), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n466), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n285), .A2(new_n257), .A3(new_n291), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n362), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n340), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n473), .B1(new_n466), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(G78gat), .B(G106gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n479), .B(KEYINPUT31), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n474), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n480), .ZN(new_n482));
  INV_X1    g281(.A(new_n473), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n294), .A2(new_n295), .A3(new_n465), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n390), .B1(new_n475), .B2(new_n362), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n466), .A2(new_n472), .A3(new_n473), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n482), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n464), .B1(new_n481), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n480), .B1(new_n474), .B2(new_n478), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n485), .B1(new_n303), .B2(new_n465), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n487), .B(new_n482), .C1(new_n491), .C2(new_n473), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(new_n492), .A3(new_n463), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n456), .B(new_n440), .C1(new_n444), .C2(new_n446), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n489), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n419), .B1(new_n462), .B2(new_n495), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n490), .A2(new_n492), .A3(new_n463), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n463), .B1(new_n490), .B2(new_n492), .ZN(new_n498));
  INV_X1    g297(.A(new_n494), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n447), .A2(new_n460), .A3(new_n457), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n460), .B1(new_n447), .B2(new_n457), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n500), .A2(new_n503), .A3(KEYINPUT89), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n418), .A2(new_n496), .A3(new_n504), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n505), .A2(KEYINPUT90), .A3(KEYINPUT35), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT90), .B1(new_n505), .B2(KEYINPUT35), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n416), .A2(new_n417), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n458), .A2(new_n494), .ZN(new_n510));
  OR3_X1    g309(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT35), .ZN(new_n511));
  NOR4_X1   g310(.A1(new_n509), .A2(new_n315), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  NOR3_X1   g311(.A1(new_n506), .A2(new_n507), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n503), .A2(KEYINPUT36), .A3(new_n494), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT36), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n497), .A2(new_n498), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n517), .B1(new_n418), .B2(new_n518), .ZN(new_n519));
  OR3_X1    g318(.A1(new_n412), .A2(KEYINPUT39), .A3(new_n358), .ZN(new_n520));
  OR2_X1    g319(.A1(new_n357), .A2(new_n359), .ZN(new_n521));
  OAI211_X1 g320(.A(KEYINPUT39), .B(new_n521), .C1(new_n412), .C2(new_n358), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(new_n407), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT40), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n520), .A2(KEYINPUT40), .A3(new_n407), .A4(new_n522), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(new_n415), .A3(new_n526), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT86), .ZN(new_n529));
  OR3_X1    g328(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n529), .B1(new_n527), .B2(new_n528), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n518), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT37), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n309), .B1(new_n305), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n535), .B1(new_n534), .B2(new_n305), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT38), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT87), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n297), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n270), .A2(KEYINPUT87), .A3(new_n296), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT88), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n299), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n299), .A2(new_n541), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n539), .B(new_n540), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT38), .B1(new_n544), .B2(KEYINPUT37), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n535), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n537), .A2(new_n310), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n533), .B1(new_n547), .B2(new_n509), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n519), .B1(new_n532), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n202), .B1(new_n513), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n505), .A2(KEYINPUT35), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT90), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n505), .A2(KEYINPUT90), .A3(KEYINPUT35), .ZN(new_n554));
  OR4_X1    g353(.A1(new_n509), .A2(new_n315), .A3(new_n510), .A4(new_n511), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n532), .A2(new_n548), .ZN(new_n557));
  INV_X1    g356(.A(new_n519), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n556), .A2(new_n559), .A3(KEYINPUT91), .ZN(new_n560));
  XNOR2_X1  g359(.A(G43gat), .B(G50gat), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n561), .A2(KEYINPUT15), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(KEYINPUT15), .ZN(new_n563));
  INV_X1    g362(.A(G29gat), .ZN(new_n564));
  INV_X1    g363(.A(G36gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n564), .A2(new_n565), .A3(KEYINPUT14), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT14), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n567), .B1(G29gat), .B2(G36gat), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n566), .B(new_n568), .C1(new_n564), .C2(new_n565), .ZN(new_n569));
  OR3_X1    g368(.A1(new_n562), .A2(new_n563), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT92), .ZN(new_n571));
  OR2_X1    g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n570), .A2(new_n571), .B1(new_n569), .B2(new_n562), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT17), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G15gat), .B(G22gat), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT16), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n575), .B1(new_n576), .B2(G1gat), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n577), .B1(G1gat), .B2(new_n575), .ZN(new_n578));
  INV_X1    g377(.A(G8gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n574), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n572), .A2(new_n573), .A3(KEYINPUT17), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n572), .A2(new_n573), .ZN(new_n584));
  AOI22_X1  g383(.A1(new_n582), .A2(new_n583), .B1(new_n584), .B2(new_n581), .ZN(new_n585));
  NAND2_X1  g384(.A1(G229gat), .A2(G233gat), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n585), .A2(KEYINPUT18), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT93), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n585), .A2(KEYINPUT93), .A3(KEYINPUT18), .A4(new_n586), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT18), .B1(new_n585), .B2(new_n586), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n584), .B(new_n580), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n586), .B(KEYINPUT13), .Z(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n591), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G113gat), .B(G141gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT11), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(new_n218), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(G197gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT12), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n598), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n591), .A2(new_n603), .A3(new_n597), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AND3_X1   g406(.A1(new_n550), .A2(new_n560), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G57gat), .B(G64gat), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G71gat), .B(G78gat), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n613), .B(KEYINPUT94), .Z(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n581), .B1(new_n615), .B2(KEYINPUT21), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(G183gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT95), .ZN(new_n619));
  NAND2_X1  g418(.A1(G231gat), .A2(G233gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n617), .B(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n615), .A2(KEYINPUT21), .ZN(new_n623));
  XNOR2_X1  g422(.A(G127gat), .B(G155gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(new_n282), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n622), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n574), .ZN(new_n630));
  INV_X1    g429(.A(G85gat), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT96), .B1(new_n631), .B2(new_n308), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT96), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n633), .A2(G85gat), .A3(G92gat), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n634), .A3(KEYINPUT7), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT7), .ZN(new_n636));
  OAI211_X1 g435(.A(KEYINPUT96), .B(new_n636), .C1(new_n631), .C2(new_n308), .ZN(new_n637));
  NAND2_X1  g436(.A1(G99gat), .A2(G106gat), .ZN(new_n638));
  AOI22_X1  g437(.A1(KEYINPUT8), .A2(new_n638), .B1(new_n631), .B2(new_n308), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n635), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT97), .ZN(new_n641));
  XOR2_X1   g440(.A(G99gat), .B(G106gat), .Z(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n641), .B(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n630), .A2(new_n583), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n641), .B(new_n642), .ZN(new_n646));
  AND2_X1   g445(.A1(G232gat), .A2(G233gat), .ZN(new_n647));
  AOI22_X1  g446(.A1(new_n646), .A2(new_n584), .B1(KEYINPUT41), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G190gat), .B(G218gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n650), .B(new_n651), .Z(new_n652));
  AND2_X1   g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n649), .A2(new_n652), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n647), .A2(KEYINPUT41), .ZN(new_n655));
  XNOR2_X1  g454(.A(G134gat), .B(G162gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  OR3_X1    g457(.A1(new_n653), .A2(new_n654), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n658), .B1(new_n653), .B2(new_n654), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n629), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(G230gat), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n664), .A2(new_n204), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n644), .A2(new_n614), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n646), .A2(new_n613), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT10), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n615), .A2(KEYINPUT10), .A3(new_n646), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n665), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n666), .A2(new_n667), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n665), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(G120gat), .B(G148gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(G176gat), .ZN(new_n677));
  INV_X1    g476(.A(G204gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n672), .A2(new_n674), .A3(new_n679), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n663), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n608), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n685), .A2(new_n508), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT100), .B(G1gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1324gat));
  NOR2_X1   g487(.A1(new_n685), .A2(new_n528), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n689), .A2(new_n579), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT42), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT16), .B(G8gat), .Z(new_n692));
  NAND2_X1  g491(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n690), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(new_n691), .B2(new_n693), .ZN(G1325gat));
  OAI21_X1  g494(.A(G15gat), .B1(new_n685), .B2(new_n517), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n510), .A2(G15gat), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n696), .B1(new_n685), .B2(new_n697), .ZN(G1326gat));
  NOR2_X1   g497(.A1(new_n685), .A2(new_n518), .ZN(new_n699));
  XOR2_X1   g498(.A(KEYINPUT43), .B(G22gat), .Z(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  INV_X1    g500(.A(new_n629), .ZN(new_n702));
  INV_X1    g501(.A(new_n683), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n702), .A2(new_n661), .A3(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n608), .A2(new_n564), .A3(new_n509), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT45), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n662), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n550), .A2(new_n560), .A3(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n507), .A2(new_n512), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n549), .B1(new_n711), .B2(new_n554), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n708), .B1(new_n712), .B2(new_n662), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n683), .B(KEYINPUT101), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n606), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n603), .B1(new_n591), .B2(new_n597), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n716), .A2(new_n719), .A3(new_n629), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n714), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(G29gat), .B1(new_n721), .B2(new_n508), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n722), .ZN(G1328gat));
  NAND4_X1  g522(.A1(new_n608), .A2(new_n565), .A3(new_n315), .A4(new_n705), .ZN(new_n724));
  XOR2_X1   g523(.A(new_n724), .B(KEYINPUT46), .Z(new_n725));
  OAI21_X1  g524(.A(G36gat), .B1(new_n721), .B2(new_n528), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(G1329gat));
  INV_X1    g526(.A(new_n517), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n710), .A2(new_n728), .A3(new_n713), .A4(new_n720), .ZN(new_n729));
  OR3_X1    g528(.A1(new_n704), .A2(G43gat), .A3(new_n510), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  AOI22_X1  g530(.A1(new_n729), .A2(G43gat), .B1(new_n608), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n732), .A2(KEYINPUT47), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n733), .A2(KEYINPUT102), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT102), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n732), .A2(new_n735), .A3(KEYINPUT47), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT103), .B1(new_n732), .B2(KEYINPUT47), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n732), .A2(KEYINPUT103), .A3(KEYINPUT47), .ZN(new_n738));
  OAI22_X1  g537(.A1(new_n734), .A2(new_n736), .B1(new_n737), .B2(new_n738), .ZN(G1330gat));
  NAND3_X1  g538(.A1(new_n714), .A2(new_n533), .A3(new_n720), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(G50gat), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT104), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT48), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n704), .A2(G50gat), .A3(new_n518), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n608), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n741), .B(new_n745), .C1(new_n742), .C2(KEYINPUT48), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(G1331gat));
  INV_X1    g548(.A(KEYINPUT105), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n716), .A2(new_n719), .A3(new_n629), .A4(new_n662), .ZN(new_n751));
  OR3_X1    g550(.A1(new_n712), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n712), .B2(new_n751), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n509), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g556(.A(new_n528), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  OR3_X1    g558(.A1(new_n754), .A2(KEYINPUT106), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT106), .B1(new_n754), .B2(new_n759), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n762), .B(new_n763), .ZN(G1333gat));
  OAI21_X1  g563(.A(G71gat), .B1(new_n754), .B2(new_n517), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n458), .A2(new_n430), .A3(new_n494), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n765), .B1(new_n754), .B2(new_n766), .ZN(new_n767));
  XOR2_X1   g566(.A(new_n767), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g567(.A1(new_n754), .A2(new_n518), .ZN(new_n769));
  XNOR2_X1  g568(.A(KEYINPUT107), .B(G78gat), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n769), .B(new_n770), .ZN(G1335gat));
  NOR2_X1   g570(.A1(new_n629), .A2(new_n607), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n683), .ZN(new_n773));
  XOR2_X1   g572(.A(new_n773), .B(KEYINPUT108), .Z(new_n774));
  NAND2_X1  g573(.A1(new_n714), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(G85gat), .B1(new_n775), .B2(new_n508), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n712), .A2(new_n662), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT51), .B1(new_n777), .B2(new_n772), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n556), .A2(new_n559), .ZN(new_n779));
  AND4_X1   g578(.A1(KEYINPUT51), .A2(new_n779), .A3(new_n661), .A4(new_n772), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n683), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n509), .A2(new_n631), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n776), .B1(new_n782), .B2(new_n783), .ZN(G1336gat));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n710), .A2(new_n315), .A3(new_n713), .A4(new_n774), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G92gat), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT109), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n715), .A2(G92gat), .A3(new_n528), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(new_n778), .B2(new_n780), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n788), .B1(new_n787), .B2(new_n790), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n785), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n787), .A2(new_n790), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT109), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n795), .A2(KEYINPUT52), .A3(new_n796), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n793), .A2(new_n797), .ZN(G1337gat));
  OAI21_X1  g597(.A(G99gat), .B1(new_n775), .B2(new_n517), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n458), .A2(new_n427), .A3(new_n494), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n799), .B1(new_n782), .B2(new_n800), .ZN(G1338gat));
  NAND3_X1  g600(.A1(new_n714), .A2(new_n533), .A3(new_n774), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(G106gat), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n715), .A2(G106gat), .A3(new_n518), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n781), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n803), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  XOR2_X1   g606(.A(new_n805), .B(KEYINPUT110), .Z(new_n808));
  NAND3_X1  g607(.A1(new_n781), .A2(KEYINPUT111), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n808), .B1(new_n778), .B2(new_n780), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT111), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n803), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n807), .B1(new_n813), .B2(new_n804), .ZN(G1339gat));
  NAND3_X1  g613(.A1(new_n669), .A2(new_n665), .A3(new_n670), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n672), .A2(KEYINPUT54), .A3(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n679), .B1(new_n671), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT55), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n816), .A2(KEYINPUT55), .A3(new_n818), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n607), .A2(new_n820), .A3(new_n682), .A4(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(KEYINPUT112), .B1(new_n585), .B2(new_n586), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n593), .A2(new_n595), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n585), .A2(KEYINPUT112), .A3(new_n586), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n602), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT113), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT113), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n829), .B(new_n602), .C1(new_n825), .C2(new_n826), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n683), .A2(new_n828), .A3(new_n606), .A4(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n661), .B1(new_n822), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n820), .A2(new_n661), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n828), .A2(new_n606), .A3(new_n830), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n821), .A2(new_n682), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n702), .B1(new_n832), .B2(new_n836), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n663), .A2(new_n607), .A3(new_n683), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n533), .A2(new_n510), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n508), .A2(new_n315), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(G113gat), .B1(new_n844), .B2(new_n719), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n508), .B1(new_n837), .B2(new_n839), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n496), .A2(new_n504), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(new_n315), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n607), .A2(new_n341), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(KEYINPUT114), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n845), .A2(new_n852), .ZN(G1340gat));
  OAI21_X1  g652(.A(G120gat), .B1(new_n844), .B2(new_n715), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT115), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n849), .A2(new_n342), .A3(new_n683), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1341gat));
  OAI21_X1  g656(.A(G127gat), .B1(new_n844), .B2(new_n702), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n849), .A2(new_n349), .A3(new_n629), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1342gat));
  NAND2_X1  g659(.A1(new_n661), .A2(new_n528), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n861), .B(KEYINPUT116), .ZN(new_n862));
  OR3_X1    g661(.A1(new_n848), .A2(G134gat), .A3(new_n862), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n864));
  OAI21_X1  g663(.A(G134gat), .B1(new_n844), .B2(new_n662), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(G1343gat));
  OR2_X1    g666(.A1(new_n846), .A2(KEYINPUT121), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n728), .A2(new_n518), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n870), .B1(new_n846), .B2(KEYINPUT121), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n719), .A2(G141gat), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n868), .A2(new_n871), .A3(new_n528), .A4(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n821), .B(new_n682), .C1(new_n717), .C2(new_n718), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n831), .B1(new_n876), .B2(new_n819), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n662), .ZN(new_n878));
  INV_X1    g677(.A(new_n836), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n629), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI211_X1 g679(.A(KEYINPUT121), .B(new_n509), .C1(new_n880), .C2(new_n838), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n869), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n846), .A2(KEYINPUT121), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n884), .A2(KEYINPUT122), .A3(new_n528), .A4(new_n872), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n875), .A2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n843), .A2(new_n517), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT117), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n518), .B1(new_n837), .B2(new_n839), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT57), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(new_n876), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n819), .B(KEYINPUT119), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT118), .ZN(new_n895));
  AOI22_X1  g694(.A1(new_n893), .A2(new_n894), .B1(new_n895), .B2(new_n831), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n831), .A2(new_n895), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n661), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n702), .B1(new_n898), .B2(new_n836), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n518), .B1(new_n899), .B2(new_n839), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n607), .B(new_n892), .C1(new_n900), .C2(new_n891), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT58), .B1(new_n901), .B2(G141gat), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n886), .A2(new_n887), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n887), .B1(new_n886), .B2(new_n902), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n893), .A2(new_n894), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n831), .A2(new_n895), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n905), .A2(new_n897), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n836), .B1(new_n907), .B2(new_n662), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n839), .B1(new_n908), .B2(new_n629), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n891), .B1(new_n909), .B2(new_n533), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n890), .A2(new_n891), .ZN(new_n911));
  INV_X1    g710(.A(new_n889), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT120), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n915), .B(new_n892), .C1(new_n900), .C2(new_n891), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n914), .A2(new_n916), .A3(new_n607), .ZN(new_n917));
  INV_X1    g716(.A(new_n884), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n918), .A2(new_n315), .ZN(new_n919));
  AOI22_X1  g718(.A1(new_n917), .A2(G141gat), .B1(new_n919), .B2(new_n872), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT58), .ZN(new_n921));
  OAI22_X1  g720(.A1(new_n903), .A2(new_n904), .B1(new_n920), .B2(new_n921), .ZN(G1344gat));
  INV_X1    g721(.A(G148gat), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n923), .A2(KEYINPUT59), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n914), .A2(new_n916), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n924), .B1(new_n925), .B2(new_n703), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n900), .A2(new_n891), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n890), .A2(new_n891), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n683), .ZN(new_n930));
  OAI21_X1  g729(.A(G148gat), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT59), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n926), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n919), .A2(new_n923), .A3(new_n683), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1345gat));
  OAI21_X1  g734(.A(G155gat), .B1(new_n925), .B2(new_n702), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n919), .A2(new_n324), .A3(new_n629), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1346gat));
  OAI21_X1  g737(.A(G162gat), .B1(new_n925), .B2(new_n662), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n862), .A2(G162gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n918), .B2(new_n940), .ZN(G1347gat));
  AOI21_X1  g740(.A(new_n509), .B1(new_n837), .B2(new_n839), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n942), .A2(new_n315), .A3(new_n847), .ZN(new_n943));
  AOI21_X1  g742(.A(G169gat), .B1(new_n943), .B2(new_n607), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n509), .A2(new_n528), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n840), .A2(new_n841), .A3(new_n945), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n719), .A2(new_n218), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(G1348gat));
  AOI21_X1  g747(.A(G176gat), .B1(new_n943), .B2(new_n683), .ZN(new_n949));
  XOR2_X1   g748(.A(new_n949), .B(KEYINPUT124), .Z(new_n950));
  INV_X1    g749(.A(new_n946), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n951), .A2(new_n247), .A3(new_n715), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n950), .A2(new_n952), .ZN(G1349gat));
  OAI21_X1  g752(.A(G183gat), .B1(new_n951), .B2(new_n702), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n943), .A2(new_n214), .A3(new_n629), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g756(.A1(new_n943), .A2(new_n210), .A3(new_n661), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT125), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n946), .A2(new_n661), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n959), .B1(new_n960), .B2(G190gat), .ZN(new_n961));
  AOI211_X1 g760(.A(KEYINPUT125), .B(new_n210), .C1(new_n946), .C2(new_n661), .ZN(new_n962));
  OR2_X1    g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n963), .A2(KEYINPUT61), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n963), .A2(KEYINPUT61), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n958), .B1(new_n964), .B2(new_n965), .ZN(G1351gat));
  AND3_X1   g765(.A1(new_n942), .A2(new_n315), .A3(new_n869), .ZN(new_n967));
  AOI21_X1  g766(.A(G197gat), .B1(new_n967), .B2(new_n607), .ZN(new_n968));
  INV_X1    g767(.A(new_n929), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n728), .A2(new_n509), .A3(new_n528), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g770(.A(new_n971), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n607), .A2(G197gat), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n968), .B1(new_n972), .B2(new_n973), .ZN(G1352gat));
  OAI21_X1  g773(.A(G204gat), .B1(new_n971), .B2(new_n715), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n967), .A2(new_n678), .A3(new_n683), .ZN(new_n976));
  AND2_X1   g775(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n977));
  NOR2_X1   g776(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI211_X1 g778(.A(new_n975), .B(new_n979), .C1(new_n977), .C2(new_n976), .ZN(G1353gat));
  NAND4_X1  g779(.A1(new_n927), .A2(new_n629), .A3(new_n928), .A4(new_n970), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(G211gat), .ZN(new_n982));
  OR2_X1    g781(.A1(new_n982), .A2(KEYINPUT63), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(KEYINPUT63), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n967), .A2(new_n282), .A3(new_n629), .ZN(new_n985));
  XOR2_X1   g784(.A(new_n985), .B(KEYINPUT127), .Z(new_n986));
  NAND3_X1  g785(.A1(new_n983), .A2(new_n984), .A3(new_n986), .ZN(G1354gat));
  AOI21_X1  g786(.A(G218gat), .B1(new_n967), .B2(new_n661), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n662), .A2(new_n287), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n988), .B1(new_n972), .B2(new_n989), .ZN(G1355gat));
endmodule


