//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1247, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1302, new_n1303, new_n1304, new_n1305;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g0005(.A(G50), .B1(G58), .B2(G68), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT64), .Z(new_n207));
  AND2_X1   g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G20), .ZN(new_n209));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR3_X1   g0011(.A1(new_n210), .A2(new_n211), .A3(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT0), .ZN(new_n214));
  OAI22_X1  g0014(.A1(new_n207), .A2(new_n209), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G116), .A2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n222));
  INV_X1    g0022(.A(G226), .ZN(new_n223));
  INV_X1    g0023(.A(G68), .ZN(new_n224));
  INV_X1    g0024(.A(G238), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n222), .B1(new_n202), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI211_X1 g0026(.A(new_n221), .B(new_n226), .C1(G97), .C2(G257), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(G1), .B2(G20), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT1), .Z(new_n229));
  AOI211_X1 g0029(.A(new_n215), .B(new_n229), .C1(new_n214), .C2(new_n213), .ZN(G361));
  XOR2_X1   g0030(.A(G250), .B(G257), .Z(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT66), .Z(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G238), .B(G244), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n234), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT67), .ZN(new_n244));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XOR2_X1   g0045(.A(G50), .B(G58), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(KEYINPUT16), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n252), .A2(new_n211), .A3(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT7), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g0056(.A1(new_n252), .A2(KEYINPUT7), .A3(new_n211), .A4(new_n253), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n224), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G58), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(new_n224), .ZN(new_n260));
  OAI21_X1  g0060(.A(G20), .B1(new_n260), .B2(new_n201), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G159), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n249), .B1(new_n258), .B2(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(KEYINPUT7), .B1(new_n268), .B2(new_n211), .ZN(new_n269));
  INV_X1    g0069(.A(new_n257), .ZN(new_n270));
  OAI21_X1  g0070(.A(G68), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n264), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(KEYINPUT16), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G1), .A2(G13), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n265), .A2(new_n273), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n274), .A2(KEYINPUT70), .A3(new_n275), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(KEYINPUT70), .B1(new_n274), .B2(new_n275), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n210), .A2(G13), .A3(G20), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT8), .B(G58), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n285), .B1(new_n210), .B2(G20), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n284), .A2(new_n286), .B1(new_n285), .B2(new_n283), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n277), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT69), .ZN(new_n289));
  AND2_X1   g0089(.A1(G33), .A2(G41), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n289), .B1(new_n290), .B2(new_n275), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G41), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n208), .A2(KEYINPUT69), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G223), .ZN(new_n295));
  INV_X1    g0095(.A(G1698), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n223), .A2(G1698), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n297), .B(new_n298), .C1(new_n266), .C2(new_n267), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G33), .A2(G87), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT80), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n299), .A2(KEYINPUT80), .A3(new_n300), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n294), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n292), .A2(G1), .A3(G13), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n306), .A2(G232), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT81), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT81), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n306), .A2(new_n307), .A3(new_n310), .A4(G232), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G274), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n313), .B1(new_n208), .B2(new_n292), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT68), .ZN(new_n315));
  NOR2_X1   g0115(.A1(G41), .A2(G45), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n315), .B1(new_n316), .B2(G1), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n210), .B(KEYINPUT68), .C1(G41), .C2(G45), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n314), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n312), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(G169), .B1(new_n305), .B2(new_n320), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n291), .A2(new_n293), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n299), .A2(KEYINPUT80), .A3(new_n300), .ZN(new_n323));
  AOI21_X1  g0123(.A(KEYINPUT80), .B1(new_n299), .B2(new_n300), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n317), .A2(new_n318), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n309), .A2(new_n311), .B1(new_n326), .B2(new_n314), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n325), .A2(new_n327), .A3(G179), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n321), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n288), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT18), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n288), .A2(new_n329), .A3(KEYINPUT18), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NOR3_X1   g0134(.A1(new_n305), .A2(new_n320), .A3(G190), .ZN(new_n335));
  AOI21_X1  g0135(.A(G200), .B1(new_n325), .B2(new_n327), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n287), .B(new_n277), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT17), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n337), .B(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(G20), .A2(G77), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n211), .A2(G33), .ZN(new_n342));
  XOR2_X1   g0142(.A(KEYINPUT15), .B(G87), .Z(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT71), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n285), .B(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n262), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n341), .B1(new_n342), .B2(new_n344), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n348), .A2(new_n276), .B1(new_n217), .B2(new_n283), .ZN(new_n349));
  INV_X1    g0149(.A(new_n276), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n210), .A2(G20), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(G77), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT3), .B(G33), .ZN(new_n354));
  NAND2_X1  g0154(.A1(G238), .A2(G1698), .ZN(new_n355));
  INV_X1    g0155(.A(G232), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n354), .B(new_n355), .C1(new_n356), .C2(G1698), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n322), .B(new_n357), .C1(G107), .C2(new_n354), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n306), .A2(new_n307), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n358), .B(new_n319), .C1(new_n218), .C2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G169), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n360), .A2(G179), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n353), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G190), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n360), .A2(G200), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n366), .A2(new_n367), .A3(new_n349), .A4(new_n352), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  OR2_X1    g0169(.A1(new_n369), .A2(KEYINPUT72), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n296), .A2(G222), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n354), .B(new_n371), .C1(new_n295), .C2(new_n296), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n322), .B(new_n372), .C1(G77), .C2(new_n354), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n373), .B(new_n319), .C1(new_n223), .C2(new_n359), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n374), .A2(new_n365), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT73), .B1(new_n374), .B2(G200), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n203), .A2(G20), .ZN(new_n377));
  INV_X1    g0177(.A(G150), .ZN(new_n378));
  OAI221_X1 g0178(.A(new_n377), .B1(new_n378), .B2(new_n347), .C1(new_n342), .C2(new_n285), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n379), .A2(new_n281), .B1(new_n202), .B2(new_n283), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n284), .A2(G50), .A3(new_n351), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT9), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n381), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT9), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n375), .A2(new_n376), .A3(new_n382), .A4(new_n385), .ZN(new_n386));
  OR2_X1    g0186(.A1(new_n386), .A2(KEYINPUT10), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(KEYINPUT10), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OR2_X1    g0189(.A1(new_n374), .A2(G179), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n374), .A2(new_n361), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(new_n383), .A3(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n340), .A2(new_n370), .A3(new_n389), .A4(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n319), .A2(KEYINPUT74), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT74), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n314), .A2(new_n317), .A3(new_n395), .A4(new_n318), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n306), .A2(G238), .A3(new_n307), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n356), .A2(G1698), .ZN(new_n399));
  OAI221_X1 g0199(.A(new_n399), .B1(G226), .B2(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G33), .A2(G97), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n322), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n397), .A2(new_n398), .A3(new_n403), .ZN(new_n404));
  XNOR2_X1  g0204(.A(KEYINPUT75), .B(KEYINPUT13), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n405), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n394), .A2(new_n396), .B1(new_n402), .B2(new_n322), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n407), .B1(new_n408), .B2(new_n398), .ZN(new_n409));
  OAI21_X1  g0209(.A(G169), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT79), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n411), .A2(KEYINPUT14), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n404), .A2(KEYINPUT76), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT76), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n408), .A2(new_n416), .A3(new_n398), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(KEYINPUT13), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n408), .A2(new_n407), .A3(new_n398), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n418), .A2(G179), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n404), .A2(new_n405), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n419), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n422), .A2(G169), .A3(new_n412), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n411), .A2(KEYINPUT14), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n414), .A2(new_n420), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n262), .A2(G50), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT78), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n426), .A2(new_n427), .B1(G20), .B2(new_n224), .ZN(new_n428));
  OAI221_X1 g0228(.A(new_n428), .B1(new_n427), .B2(new_n426), .C1(new_n217), .C2(new_n342), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n281), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT11), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n210), .A2(new_n224), .A3(G13), .A4(G20), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n433), .B(KEYINPUT12), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n429), .A2(KEYINPUT11), .A3(new_n281), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n350), .A2(G68), .A3(new_n351), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n432), .A2(new_n434), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n425), .A2(new_n437), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n419), .A2(G190), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n418), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT77), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n437), .B1(new_n422), .B2(G200), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT77), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n418), .A2(new_n439), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n369), .A2(KEYINPUT72), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n438), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n393), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n225), .A2(new_n296), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n218), .A2(G1698), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n449), .B(new_n450), .C1(new_n266), .C2(new_n267), .ZN(new_n451));
  INV_X1    g0251(.A(G116), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n251), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n322), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(G45), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(G1), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n313), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n459), .B(new_n306), .C1(G250), .C2(new_n458), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G190), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n343), .A2(new_n282), .ZN(new_n463));
  INV_X1    g0263(.A(G97), .ZN(new_n464));
  INV_X1    g0264(.A(G107), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n219), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n401), .A2(new_n211), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n466), .A2(new_n467), .A3(KEYINPUT19), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n211), .B(G68), .C1(new_n266), .C2(new_n267), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT19), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n470), .B1(new_n342), .B2(new_n464), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n468), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n463), .B1(new_n472), .B2(new_n276), .ZN(new_n473));
  INV_X1    g0273(.A(new_n280), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n278), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n210), .A2(G33), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n475), .A2(G87), .A3(new_n282), .A4(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G200), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n479), .B1(new_n456), .B2(new_n460), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n451), .A2(new_n454), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n460), .B1(new_n482), .B2(new_n294), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n475), .A2(new_n343), .A3(new_n282), .A4(new_n476), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n361), .A2(new_n483), .B1(new_n473), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G179), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n461), .A2(new_n486), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n462), .A2(new_n481), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G41), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n210), .B(G45), .C1(new_n489), .C2(KEYINPUT5), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT83), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT83), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT5), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G41), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n458), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n493), .A2(G41), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n491), .A2(new_n495), .A3(new_n314), .A4(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(G244), .B(new_n296), .C1(new_n266), .C2(new_n267), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n354), .A2(KEYINPUT4), .A3(G244), .A4(new_n296), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n354), .A2(G250), .A3(G1698), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G283), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT82), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(KEYINPUT82), .A2(G33), .A3(G283), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n502), .A2(new_n503), .A3(new_n504), .A4(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n499), .B1(new_n510), .B2(new_n322), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n490), .A2(new_n496), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n512), .B1(new_n208), .B2(new_n292), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G257), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n511), .A2(G179), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n510), .A2(new_n322), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n516), .A2(new_n514), .A3(new_n498), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n515), .B1(new_n517), .B2(new_n361), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n283), .A2(new_n464), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n282), .B(new_n476), .C1(new_n279), .C2(new_n280), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n520), .A2(new_n464), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n465), .B1(new_n256), .B2(new_n257), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n347), .A2(new_n217), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT6), .ZN(new_n525));
  AND2_X1   g0325(.A1(G97), .A2(G107), .ZN(new_n526));
  NOR2_X1   g0326(.A1(G97), .A2(G107), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n465), .A2(KEYINPUT6), .A3(G97), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n211), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n523), .A2(new_n524), .A3(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n519), .B(new_n522), .C1(new_n531), .C2(new_n350), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n532), .A2(KEYINPUT84), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT84), .ZN(new_n534));
  OAI21_X1  g0334(.A(G107), .B1(new_n269), .B2(new_n270), .ZN(new_n535));
  INV_X1    g0335(.A(new_n524), .ZN(new_n536));
  INV_X1    g0336(.A(new_n530), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n521), .B1(new_n538), .B2(new_n276), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n534), .B1(new_n539), .B2(new_n519), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n518), .B1(new_n533), .B2(new_n540), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n511), .A2(G190), .A3(new_n514), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n479), .B1(new_n511), .B2(new_n514), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n532), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n520), .A2(new_n465), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n211), .B(G87), .C1(new_n266), .C2(new_n267), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT22), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT22), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n354), .A2(new_n550), .A3(new_n211), .A4(G87), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(KEYINPUT90), .A2(KEYINPUT23), .A3(G107), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT90), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(G20), .B2(new_n465), .ZN(new_n555));
  AOI22_X1  g0355(.A1(KEYINPUT90), .A2(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n556));
  OAI22_X1  g0356(.A1(new_n555), .A2(KEYINPUT23), .B1(new_n556), .B2(G20), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n552), .A2(new_n553), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT24), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n557), .B1(new_n549), .B2(new_n551), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT24), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(new_n562), .A3(new_n553), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n547), .B1(new_n564), .B2(new_n276), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n513), .A2(G264), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n268), .B1(new_n220), .B2(new_n296), .ZN(new_n567));
  OR2_X1    g0367(.A1(new_n296), .A2(G257), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n567), .A2(new_n568), .B1(G33), .B2(G294), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n566), .B(new_n498), .C1(new_n569), .C2(new_n294), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G190), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(G200), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n283), .A2(new_n465), .ZN(new_n574));
  XNOR2_X1  g0374(.A(new_n574), .B(KEYINPUT91), .ZN(new_n575));
  XNOR2_X1  g0375(.A(new_n575), .B(KEYINPUT25), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n565), .A2(new_n572), .A3(new_n573), .A4(new_n576), .ZN(new_n577));
  AND4_X1   g0377(.A1(new_n488), .A2(new_n541), .A3(new_n546), .A4(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT89), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n579), .A2(KEYINPUT21), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT21), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n581), .A2(KEYINPUT89), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n296), .A2(G257), .ZN(new_n583));
  NAND2_X1  g0383(.A1(G264), .A2(G1698), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n583), .B(new_n584), .C1(new_n266), .C2(new_n267), .ZN(new_n585));
  INV_X1    g0385(.A(G303), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n252), .A2(new_n586), .A3(new_n253), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n585), .A2(new_n291), .A3(new_n587), .A4(new_n293), .ZN(new_n588));
  OAI211_X1 g0388(.A(G270), .B(new_n306), .C1(new_n490), .C2(new_n496), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n498), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n590), .A2(G169), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT85), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n282), .A2(new_n275), .A3(new_n274), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n476), .A2(G116), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n452), .B1(new_n210), .B2(G33), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n350), .A2(KEYINPUT85), .A3(new_n282), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n211), .B1(new_n464), .B2(G33), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n507), .B2(new_n508), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n274), .A2(new_n275), .B1(G20), .B2(new_n452), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(KEYINPUT87), .B(KEYINPUT20), .C1(new_n600), .C2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n282), .A2(G116), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT86), .ZN(new_n605));
  XNOR2_X1  g0405(.A(new_n604), .B(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n599), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n509), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(KEYINPUT87), .A2(KEYINPUT20), .ZN(new_n609));
  OR2_X1    g0409(.A1(KEYINPUT87), .A2(KEYINPUT20), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n608), .A2(new_n609), .A3(new_n610), .A4(new_n601), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n598), .A2(new_n603), .A3(new_n606), .A4(new_n611), .ZN(new_n612));
  AOI211_X1 g0412(.A(new_n580), .B(new_n582), .C1(new_n591), .C2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n590), .A2(KEYINPUT21), .A3(G169), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n498), .A2(new_n588), .A3(G179), .A4(new_n589), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n612), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT88), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n616), .A2(KEYINPUT88), .A3(new_n612), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n613), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AND4_X1   g0421(.A1(new_n562), .A2(new_n552), .A3(new_n553), .A4(new_n558), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n562), .B1(new_n561), .B2(new_n553), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n276), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n547), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(new_n625), .A3(new_n576), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n570), .A2(new_n361), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n571), .A2(new_n486), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  AND4_X1   g0429(.A1(new_n598), .A2(new_n603), .A3(new_n606), .A4(new_n611), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n590), .A2(G200), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n630), .B(new_n631), .C1(new_n365), .C2(new_n590), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n621), .A2(new_n629), .A3(new_n632), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n448), .A2(new_n578), .A3(new_n633), .ZN(G372));
  INV_X1    g0434(.A(new_n364), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n445), .A2(new_n635), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n636), .A2(KEYINPUT92), .A3(new_n438), .ZN(new_n637));
  AOI21_X1  g0437(.A(KEYINPUT92), .B1(new_n636), .B2(new_n438), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n637), .A2(new_n638), .A3(new_n339), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n389), .B1(new_n639), .B2(new_n334), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT93), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(new_n641), .A3(new_n392), .ZN(new_n642));
  INV_X1    g0442(.A(new_n389), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n636), .A2(new_n438), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT92), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n337), .B(KEYINPUT17), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n636), .A2(KEYINPUT92), .A3(new_n438), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n332), .A2(new_n333), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n643), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n392), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT93), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n642), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n448), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n485), .A2(new_n487), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n488), .B(new_n518), .C1(new_n533), .C2(new_n540), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n657), .B1(new_n658), .B2(KEYINPUT26), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n518), .A2(new_n532), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT26), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(new_n662), .A3(new_n488), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n541), .A2(new_n577), .A3(new_n546), .A4(new_n488), .ZN(new_n664));
  INV_X1    g0464(.A(new_n580), .ZN(new_n665));
  INV_X1    g0465(.A(new_n582), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n590), .A2(G169), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n665), .B(new_n666), .C1(new_n630), .C2(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n668), .A2(new_n617), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n629), .A2(new_n669), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n659), .B(new_n663), .C1(new_n664), .C2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n654), .B1(new_n655), .B2(new_n672), .ZN(G369));
  NAND3_X1  g0473(.A1(new_n210), .A2(new_n211), .A3(G13), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G213), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(G343), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n626), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n577), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n629), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n629), .A2(new_n679), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n621), .A2(new_n679), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n686), .A2(new_n683), .ZN(new_n687));
  INV_X1    g0487(.A(new_n679), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n630), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n669), .A2(new_n689), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n690), .B(new_n632), .C1(new_n621), .C2(new_n689), .ZN(new_n691));
  INV_X1    g0491(.A(G330), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n684), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n687), .B1(new_n694), .B2(new_n695), .ZN(G399));
  NOR2_X1   g0496(.A1(new_n466), .A2(G116), .ZN(new_n697));
  XOR2_X1   g0497(.A(new_n697), .B(KEYINPUT94), .Z(new_n698));
  INV_X1    g0498(.A(new_n212), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(G41), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n698), .A2(G1), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n206), .B2(new_n701), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT28), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n671), .A2(new_n688), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n705), .A2(KEYINPUT29), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n619), .A2(new_n620), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n629), .A2(new_n707), .A3(new_n668), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n481), .A2(new_n462), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n532), .A2(KEYINPUT84), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n539), .A2(new_n534), .A3(new_n519), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI22_X1  g0512(.A1(new_n712), .A2(new_n518), .B1(new_n544), .B2(new_n545), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n708), .A2(new_n709), .A3(new_n713), .A4(new_n577), .ZN(new_n714));
  INV_X1    g0514(.A(new_n488), .ZN(new_n715));
  OAI21_X1  g0515(.A(KEYINPUT26), .B1(new_n660), .B2(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n712), .A2(new_n662), .A3(new_n488), .A4(new_n518), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n717), .A2(new_n656), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n714), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n688), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(KEYINPUT29), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n706), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n566), .B1(new_n569), .B2(new_n294), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(new_n483), .ZN(new_n724));
  INV_X1    g0524(.A(new_n615), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(new_n517), .A3(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n517), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n590), .A2(new_n486), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n729), .A2(new_n570), .A3(new_n730), .A4(new_n483), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n724), .A2(new_n517), .A3(KEYINPUT30), .A4(new_n725), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n728), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n679), .ZN(new_n734));
  XNOR2_X1  g0534(.A(KEYINPUT95), .B(KEYINPUT31), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n578), .A2(new_n633), .A3(new_n688), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n734), .A2(new_n735), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n739), .A2(G330), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n722), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n704), .B1(new_n741), .B2(G1), .ZN(G364));
  INV_X1    g0542(.A(G13), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n743), .A2(new_n251), .A3(KEYINPUT98), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT98), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(G13), .B2(G33), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT102), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n691), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n211), .A2(G13), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT97), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n210), .B1(new_n753), .B2(G45), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n700), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n211), .A2(new_n365), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n486), .A2(new_n479), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT100), .ZN(new_n760));
  INV_X1    g0560(.A(G326), .ZN(new_n761));
  INV_X1    g0561(.A(G294), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G179), .A2(G200), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n211), .B1(new_n763), .B2(G190), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n760), .A2(new_n761), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT101), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n211), .A2(G190), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n479), .A2(G179), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G283), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n757), .A2(new_n768), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n268), .B1(new_n769), .B2(new_n770), .C1(new_n586), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n758), .A2(new_n767), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G317), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(KEYINPUT33), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n775), .A2(KEYINPUT33), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n774), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G329), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n767), .A2(new_n763), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n486), .A2(G200), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n767), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n772), .B(new_n781), .C1(G311), .C2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G322), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n757), .A2(new_n782), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n766), .B(new_n785), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n783), .A2(new_n217), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n764), .A2(new_n464), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(G68), .B2(new_n774), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT99), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n769), .A2(new_n465), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n759), .A2(new_n202), .B1(new_n787), .B2(new_n259), .ZN(new_n794));
  INV_X1    g0594(.A(new_n771), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n793), .B(new_n794), .C1(G87), .C2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT32), .ZN(new_n797));
  INV_X1    g0597(.A(new_n780), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n797), .B1(new_n798), .B2(G159), .ZN(new_n799));
  INV_X1    g0599(.A(G159), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n780), .A2(KEYINPUT32), .A3(new_n800), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n799), .A2(new_n268), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n792), .A2(new_n796), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n788), .B1(new_n789), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n275), .B1(G20), .B2(new_n361), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n749), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n247), .A2(G45), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n699), .A2(new_n354), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n807), .B(new_n808), .C1(G45), .C2(new_n207), .ZN(new_n809));
  INV_X1    g0609(.A(G355), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n354), .A2(new_n212), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n809), .B1(G116), .B2(new_n212), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n804), .A2(new_n805), .B1(new_n806), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n751), .A2(new_n756), .A3(new_n813), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n691), .A2(new_n692), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n756), .B1(new_n815), .B2(KEYINPUT96), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n694), .B1(new_n815), .B2(KEYINPUT96), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n814), .B1(new_n817), .B2(new_n818), .ZN(G396));
  NOR2_X1   g0619(.A1(new_n364), .A2(new_n679), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n353), .A2(new_n679), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n368), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n364), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n705), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n820), .B1(new_n364), .B2(new_n823), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n671), .A2(new_n688), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n740), .B(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n756), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n773), .A2(new_n770), .B1(new_n783), .B2(new_n452), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT103), .Z(new_n834));
  INV_X1    g0634(.A(new_n787), .ZN(new_n835));
  AOI22_X1  g0635(.A1(G107), .A2(new_n795), .B1(new_n835), .B2(G294), .ZN(new_n836));
  INV_X1    g0636(.A(G311), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n836), .B1(new_n219), .B2(new_n769), .C1(new_n837), .C2(new_n780), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n268), .B1(new_n759), .B2(new_n586), .ZN(new_n839));
  OR4_X1    g0639(.A1(new_n790), .A2(new_n834), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G143), .A2(new_n835), .B1(new_n774), .B2(G150), .ZN(new_n841));
  INV_X1    g0641(.A(G137), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n841), .B1(new_n842), .B2(new_n759), .C1(new_n800), .C2(new_n783), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT34), .ZN(new_n844));
  INV_X1    g0644(.A(G132), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n354), .B1(new_n780), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(G50), .B2(new_n795), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n844), .B(new_n847), .C1(new_n259), .C2(new_n764), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n769), .A2(new_n224), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n840), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n831), .B1(new_n850), .B2(new_n805), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n747), .A2(new_n805), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n851), .B1(G77), .B2(new_n853), .C1(new_n827), .C2(new_n748), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n832), .A2(new_n854), .ZN(G384));
  NAND2_X1  g0655(.A1(new_n437), .A2(new_n679), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n438), .A2(new_n445), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n425), .A2(new_n437), .A3(new_n679), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n825), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n733), .B(new_n679), .C1(KEYINPUT106), .C2(KEYINPUT31), .ZN(new_n860));
  NOR2_X1   g0660(.A1(KEYINPUT106), .A2(KEYINPUT31), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n734), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n737), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n265), .A2(new_n273), .A3(new_n281), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n287), .ZN(new_n866));
  INV_X1    g0666(.A(new_n677), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n277), .A2(new_n287), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n479), .B1(new_n305), .B2(new_n320), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n325), .A2(new_n327), .A3(new_n365), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n869), .A2(new_n872), .B1(new_n866), .B2(new_n329), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n868), .B1(new_n873), .B2(KEYINPUT104), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n866), .A2(new_n329), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n337), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT104), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT37), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n288), .A2(new_n867), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n330), .A2(new_n880), .A3(new_n337), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT105), .B1(new_n881), .B2(KEYINPUT37), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT105), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n885), .B(KEYINPUT37), .C1(new_n874), .C2(new_n878), .ZN(new_n886));
  INV_X1    g0686(.A(new_n868), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n334), .B2(new_n339), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n884), .A2(KEYINPUT38), .A3(new_n886), .A4(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n868), .B1(new_n647), .B2(new_n650), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n879), .B2(new_n883), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT38), .B1(new_n892), .B2(new_n886), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n864), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT40), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n880), .B1(new_n647), .B2(new_n650), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT37), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n881), .B(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n897), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n887), .B1(new_n876), .B2(new_n877), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n873), .A2(KEYINPUT104), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n899), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n886), .B(new_n888), .C1(new_n904), .C2(new_n882), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n901), .B1(new_n905), .B2(new_n897), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n864), .A2(new_n906), .A3(KEYINPUT40), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n896), .A2(new_n907), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n448), .A2(new_n863), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n908), .B(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(G330), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n655), .B1(new_n706), .B2(new_n721), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n642), .B2(new_n653), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT39), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n906), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n438), .A2(new_n679), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n888), .B1(new_n904), .B2(new_n882), .ZN(new_n917));
  INV_X1    g0717(.A(new_n886), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n897), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(KEYINPUT39), .A3(new_n889), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n915), .A2(new_n916), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n334), .A2(new_n677), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n828), .A2(new_n821), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n857), .A2(new_n858), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n923), .B(new_n924), .C1(new_n890), .C2(new_n893), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n921), .A2(new_n922), .A3(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n913), .B(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n911), .B(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n210), .B2(new_n753), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n528), .A2(new_n529), .ZN(new_n930));
  OAI211_X1 g0730(.A(G20), .B(new_n208), .C1(new_n930), .C2(KEYINPUT35), .ZN(new_n931));
  AOI211_X1 g0731(.A(new_n452), .B(new_n931), .C1(KEYINPUT35), .C2(new_n930), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n932), .B(KEYINPUT36), .Z(new_n933));
  OAI21_X1  g0733(.A(G77), .B1(new_n259), .B2(new_n224), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n934), .A2(new_n206), .B1(G50), .B2(new_n224), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n935), .A2(G1), .A3(new_n743), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n929), .A2(new_n933), .A3(new_n936), .ZN(G367));
  OAI21_X1  g0737(.A(new_n713), .B1(new_n545), .B2(new_n688), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n661), .A2(new_n679), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n687), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT45), .ZN(new_n943));
  OR3_X1    g0743(.A1(new_n687), .A2(KEYINPUT44), .A3(new_n941), .ZN(new_n944));
  OAI21_X1  g0744(.A(KEYINPUT44), .B1(new_n687), .B2(new_n941), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n694), .A2(new_n695), .ZN(new_n947));
  OR3_X1    g0747(.A1(new_n943), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n947), .B1(new_n943), .B2(new_n946), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n684), .A2(new_n685), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n950), .A2(new_n686), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n951), .A2(KEYINPUT110), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n952), .A2(new_n694), .ZN(new_n953));
  INV_X1    g0753(.A(new_n952), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n951), .A2(KEYINPUT110), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n953), .B1(new_n956), .B2(new_n694), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n948), .A2(new_n741), .A3(new_n949), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n741), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n700), .B(KEYINPUT41), .ZN(new_n960));
  AOI21_X1  g0760(.A(KEYINPUT111), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT111), .ZN(new_n962));
  INV_X1    g0762(.A(new_n960), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n962), .B(new_n963), .C1(new_n958), .C2(new_n741), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n754), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT109), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n686), .A2(new_n940), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT42), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT107), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n541), .B1(new_n940), .B2(new_n629), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n688), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n968), .B2(new_n967), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n478), .A2(new_n679), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n488), .A2(new_n975), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n656), .A2(new_n975), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT43), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n978), .B(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n966), .B1(new_n974), .B2(new_n981), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n974), .A2(new_n979), .A3(new_n976), .A4(new_n977), .ZN(new_n983));
  OAI211_X1 g0783(.A(KEYINPUT109), .B(new_n980), .C1(new_n970), .C2(new_n973), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n947), .A2(new_n941), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT108), .Z(new_n987));
  XNOR2_X1  g0787(.A(new_n985), .B(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n965), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n764), .A2(new_n224), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n354), .B1(new_n780), .B2(new_n842), .C1(new_n259), .C2(new_n771), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n990), .B(new_n991), .C1(G150), .C2(new_n835), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n773), .A2(new_n800), .B1(new_n769), .B2(new_n217), .ZN(new_n993));
  INV_X1    g0793(.A(new_n760), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n993), .B1(new_n994), .B2(G143), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n992), .B(new_n995), .C1(new_n202), .C2(new_n783), .ZN(new_n996));
  AOI22_X1  g0796(.A1(G294), .A2(new_n774), .B1(new_n784), .B2(G283), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n464), .B2(new_n769), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(G311), .B2(new_n994), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n771), .A2(new_n452), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n1000), .A2(KEYINPUT46), .B1(new_n465), .B2(new_n764), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n354), .B(new_n1001), .C1(KEYINPUT46), .C2(new_n1000), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n999), .B(new_n1002), .C1(new_n586), .C2(new_n787), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n780), .A2(new_n775), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n996), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT47), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n831), .B1(new_n1006), .B2(new_n805), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n808), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n806), .B1(new_n212), .B2(new_n344), .C1(new_n233), .C2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n976), .A2(new_n750), .A3(new_n977), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1007), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n989), .A2(new_n1011), .ZN(G387));
  OR2_X1    g0812(.A1(new_n957), .A2(new_n741), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n957), .A2(new_n741), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1013), .A2(new_n1014), .A3(new_n700), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n808), .B1(new_n239), .B2(new_n457), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n698), .B2(new_n811), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n346), .A2(G50), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1019), .A2(KEYINPUT50), .ZN(new_n1020));
  AOI21_X1  g0820(.A(G45), .B1(new_n1019), .B2(KEYINPUT50), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(G68), .A2(G77), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .A4(new_n698), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1017), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n699), .A2(new_n465), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n749), .B(new_n805), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n769), .A2(new_n452), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G311), .A2(new_n774), .B1(new_n784), .B2(G303), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n775), .B2(new_n787), .C1(new_n760), .C2(new_n786), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT48), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n770), .B2(new_n764), .C1(new_n762), .C2(new_n771), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT49), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n268), .B1(new_n761), .B2(new_n780), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1027), .B(new_n1033), .C1(new_n1032), .C2(new_n1031), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n285), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1035), .A2(new_n774), .B1(new_n798), .B2(G150), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n224), .B2(new_n783), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n795), .A2(G77), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1038), .B(new_n354), .C1(new_n464), .C2(new_n769), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n759), .A2(new_n800), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n344), .A2(new_n764), .B1(new_n202), .B2(new_n787), .ZN(new_n1041));
  NOR4_X1   g0841(.A1(new_n1037), .A2(new_n1039), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n805), .B1(new_n1034), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n756), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1026), .B(new_n1044), .C1(new_n695), .C2(new_n750), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n755), .B2(new_n957), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1015), .A2(new_n1046), .ZN(G393));
  NAND2_X1  g0847(.A1(new_n948), .A2(new_n949), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1048), .A2(new_n754), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n940), .A2(new_n749), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n759), .A2(new_n775), .B1(new_n787), .B2(new_n837), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT52), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1052), .B(new_n268), .C1(new_n452), .C2(new_n764), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n773), .A2(new_n586), .B1(new_n783), .B2(new_n762), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n780), .A2(new_n786), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n771), .A2(new_n770), .ZN(new_n1056));
  OR4_X1    g0856(.A1(new_n793), .A2(new_n1054), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n346), .A2(new_n783), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n764), .A2(new_n217), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(G143), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n771), .A2(new_n224), .B1(new_n780), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(G50), .B2(new_n774), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n769), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n268), .B1(new_n1064), .B2(G87), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1058), .A2(new_n1060), .A3(new_n1063), .A4(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n759), .A2(new_n378), .B1(new_n787), .B2(new_n800), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT51), .Z(new_n1068));
  OAI22_X1  g0868(.A1(new_n1053), .A2(new_n1057), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n831), .B1(new_n1069), .B2(new_n805), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1050), .A2(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n243), .A2(new_n808), .B1(G97), .B2(new_n699), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1071), .B1(new_n806), .B2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1049), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1048), .A2(new_n1014), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1075), .A2(new_n700), .A3(new_n958), .ZN(new_n1076));
  AND3_X1   g0876(.A1(new_n1074), .A2(KEYINPUT112), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(KEYINPUT112), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(G390));
  NOR2_X1   g0880(.A1(new_n825), .A2(new_n692), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n863), .A2(new_n1081), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n857), .A2(new_n858), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n916), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n923), .A2(new_n924), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n915), .A2(new_n920), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n889), .A2(new_n901), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n719), .A2(new_n688), .A3(new_n824), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1083), .B1(new_n1090), .B2(new_n821), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1089), .A2(new_n1091), .A3(new_n916), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1085), .B1(new_n1088), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1087), .A2(new_n1086), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n919), .A2(KEYINPUT39), .A3(new_n889), .ZN(new_n1095));
  AOI21_X1  g0895(.A(KEYINPUT39), .B1(new_n889), .B2(new_n901), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n1090), .A2(new_n821), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1086), .B(new_n906), .C1(new_n1098), .C2(new_n1083), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n739), .A2(new_n924), .A3(new_n1081), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1097), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1093), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n924), .B1(new_n739), .B2(new_n1081), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n923), .B1(new_n1084), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1098), .A2(new_n1106), .A3(new_n1100), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n912), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n909), .A2(G330), .ZN(new_n1110));
  AND4_X1   g0910(.A1(new_n654), .A2(new_n1108), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1093), .A2(new_n1102), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n913), .A2(new_n1110), .A3(new_n1108), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT113), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(KEYINPUT113), .B1(new_n1111), .B2(new_n1103), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n700), .B1(new_n1103), .B2(new_n1111), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1103), .A2(new_n755), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n747), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(G107), .A2(new_n774), .B1(new_n835), .B2(G116), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1120), .B1(new_n464), .B2(new_n783), .C1(new_n770), .C2(new_n759), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n268), .B1(new_n780), .B2(new_n762), .C1(new_n219), .C2(new_n771), .ZN(new_n1122));
  OR4_X1    g0922(.A1(new_n849), .A2(new_n1121), .A3(new_n1059), .A4(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n764), .A2(new_n800), .ZN(new_n1124));
  INV_X1    g0924(.A(G128), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n354), .B1(new_n773), .B2(new_n842), .C1(new_n1125), .C2(new_n759), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1124), .B(new_n1126), .C1(G50), .C2(new_n1064), .ZN(new_n1127));
  XOR2_X1   g0927(.A(KEYINPUT54), .B(G143), .Z(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(G125), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n1129), .A2(new_n783), .B1(new_n1130), .B2(new_n780), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT53), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n771), .B2(new_n378), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n795), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1131), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1127), .B(new_n1135), .C1(new_n845), .C2(new_n787), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1123), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n831), .B1(new_n1137), .B2(new_n805), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1119), .B(new_n1138), .C1(new_n1035), .C2(new_n853), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1117), .A2(new_n1118), .A3(new_n1139), .ZN(G378));
  INV_X1    g0940(.A(KEYINPUT119), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT117), .ZN(new_n1142));
  AND4_X1   g0942(.A1(new_n1142), .A2(new_n654), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1142), .B1(new_n913), .B2(new_n1110), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1114), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1111), .A2(KEYINPUT113), .A3(new_n1103), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1145), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n859), .A2(new_n863), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n889), .B2(new_n919), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n907), .B(G330), .C1(new_n1150), .C2(KEYINPUT40), .ZN(new_n1151));
  NOR3_X1   g0951(.A1(new_n643), .A2(KEYINPUT55), .A3(new_n652), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT55), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n389), .B2(new_n392), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n383), .A2(new_n867), .ZN(new_n1155));
  XOR2_X1   g0955(.A(new_n1155), .B(KEYINPUT56), .Z(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  OR3_X1    g0957(.A1(new_n1152), .A2(new_n1154), .A3(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1157), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1159));
  AND2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1151), .A2(new_n1161), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n896), .A2(G330), .A3(new_n1160), .A4(new_n907), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(KEYINPUT118), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n926), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT118), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1162), .A2(new_n1163), .A3(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1165), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1164), .A2(KEYINPUT118), .A3(new_n926), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT57), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n1148), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1141), .B1(new_n1173), .B2(new_n701), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1162), .A2(new_n1163), .A3(KEYINPUT116), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(new_n1166), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n1172), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1171), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1181), .A2(new_n1176), .A3(KEYINPUT57), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1182), .A2(KEYINPUT119), .A3(new_n700), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1174), .A2(new_n1180), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1160), .A2(new_n747), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n852), .A2(new_n202), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n759), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G116), .A2(new_n1187), .B1(new_n774), .B2(G97), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n798), .A2(G283), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1064), .A2(G58), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1188), .A2(new_n268), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1038), .B1(new_n783), .B2(new_n344), .C1(new_n465), .C2(new_n787), .ZN(new_n1192));
  NOR4_X1   g0992(.A1(new_n1191), .A2(new_n1192), .A3(G41), .A4(new_n990), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1193), .B(KEYINPUT114), .Z(new_n1194));
  NOR2_X1   g0994(.A1(new_n266), .A2(G41), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n1194), .A2(KEYINPUT58), .B1(G50), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT115), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1194), .A2(KEYINPUT58), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n787), .A2(new_n1125), .B1(new_n764), .B2(new_n378), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n795), .A2(new_n1128), .B1(new_n784), .B2(G137), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n845), .B2(new_n773), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1201), .B(new_n1203), .C1(G125), .C2(new_n1187), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT59), .ZN(new_n1205));
  AOI21_X1  g1005(.A(G41), .B1(new_n798), .B2(G124), .ZN(new_n1206));
  AOI21_X1  g1006(.A(G33), .B1(new_n1064), .B2(G159), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .A4(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n831), .B1(new_n1209), .B2(new_n805), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1185), .A2(new_n1186), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n1178), .B2(new_n755), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1184), .A2(new_n1213), .ZN(G375));
  AOI21_X1  g1014(.A(new_n1108), .B1(new_n913), .B2(new_n1110), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT120), .Z(new_n1216));
  OR3_X1    g1016(.A1(new_n1216), .A2(new_n963), .A3(new_n1111), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1083), .A2(new_n747), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n268), .B1(new_n1064), .B2(G58), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1219), .B1(new_n202), .B2(new_n764), .C1(new_n1125), .C2(new_n780), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(G137), .A2(new_n835), .B1(new_n784), .B2(G150), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1221), .B1(new_n845), .B2(new_n759), .C1(new_n800), .C2(new_n771), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n1220), .B(new_n1222), .C1(new_n774), .C2(new_n1128), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(G97), .A2(new_n795), .B1(new_n798), .B2(G303), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n465), .B2(new_n783), .C1(new_n762), .C2(new_n759), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n344), .A2(new_n764), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n773), .A2(new_n452), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n268), .B1(new_n769), .B2(new_n217), .C1(new_n770), .C2(new_n787), .ZN(new_n1228));
  NOR4_X1   g1028(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n805), .B1(new_n1223), .B2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n756), .B1(G68), .B2(new_n853), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1231), .B(KEYINPUT122), .ZN(new_n1232));
  AND3_X1   g1032(.A1(new_n1218), .A2(new_n1230), .A3(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n754), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1234), .A2(KEYINPUT121), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(KEYINPUT121), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1233), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1217), .A2(new_n1237), .ZN(G381));
  NAND3_X1  g1038(.A1(new_n989), .A2(new_n1079), .A3(new_n1011), .ZN(new_n1239));
  INV_X1    g1039(.A(G384), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1217), .A2(new_n1240), .A3(new_n1237), .ZN(new_n1241));
  NOR4_X1   g1041(.A1(new_n1239), .A2(G396), .A3(G393), .A4(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(G378), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1184), .A2(new_n1243), .A3(new_n1213), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1242), .A2(new_n1245), .ZN(G407));
  OAI21_X1  g1046(.A(new_n1245), .B1(new_n1242), .B2(new_n678), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(G213), .ZN(G409));
  XOR2_X1   g1048(.A(G393), .B(G396), .Z(new_n1249));
  INV_X1    g1049(.A(new_n1239), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1079), .B1(new_n989), .B2(new_n1011), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1249), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G387), .A2(G390), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1249), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1253), .A2(new_n1239), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1252), .A2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n678), .A2(G213), .A3(G2897), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1215), .A2(KEYINPUT60), .ZN(new_n1258));
  AND2_X1   g1058(.A1(new_n1113), .A2(KEYINPUT60), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n700), .B(new_n1258), .C1(new_n1216), .C2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1260), .A2(G384), .A3(new_n1237), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(G384), .B1(new_n1260), .B2(new_n1237), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1257), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1263), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1257), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1265), .A2(new_n1261), .A3(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1264), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1243), .B1(new_n1184), .B2(new_n1213), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1176), .A2(new_n960), .A3(new_n1178), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1181), .A2(new_n755), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1243), .A2(new_n1211), .A3(new_n1270), .A4(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n678), .A2(G213), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1268), .B1(new_n1269), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(G375), .A2(G378), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1276), .A2(new_n1277), .A3(new_n1278), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1256), .B(new_n1275), .C1(new_n1279), .C2(KEYINPUT62), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1279), .A2(KEYINPUT62), .ZN(new_n1281));
  XOR2_X1   g1081(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1282));
  NOR3_X1   g1082(.A1(new_n1280), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT63), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1279), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT123), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT61), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1276), .A2(KEYINPUT63), .A3(new_n1277), .A4(new_n1278), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT125), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1269), .A2(new_n1274), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1291), .A2(KEYINPUT125), .A3(KEYINPUT63), .A4(new_n1278), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT124), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1268), .A2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1264), .A2(new_n1267), .A3(KEYINPUT124), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1295), .B(new_n1296), .C1(new_n1269), .C2(new_n1274), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1279), .A2(KEYINPUT123), .A3(new_n1284), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1287), .A2(new_n1293), .A3(new_n1297), .A4(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1256), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1283), .B1(new_n1299), .B2(new_n1300), .ZN(G405));
  INV_X1    g1101(.A(KEYINPUT127), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1278), .A2(new_n1302), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(new_n1256), .B(new_n1303), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1276), .B(new_n1244), .C1(new_n1302), .C2(new_n1278), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(new_n1304), .B(new_n1305), .ZN(G402));
endmodule


