//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 1 0 0 0 0 0 0 1 1 0 1 1 1 0 1 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n551,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT64), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n461), .A2(G2105), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n464), .A2(G137), .B1(G101), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n467), .B1(new_n462), .B2(new_n463), .ZN(new_n468));
  AND2_X1   g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(G160));
  INV_X1    g047(.A(new_n463), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n464), .A2(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(new_n476), .B2(G112), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n478), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  OAI211_X1 g058(.A(G138), .B(new_n476), .C1(new_n473), .C2(new_n474), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n484), .B1(KEYINPUT65), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(G126), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n487), .B1(new_n462), .B2(new_n463), .ZN(new_n488));
  AND2_X1   g063(.A1(G114), .A2(G2104), .ZN(new_n489));
  OAI21_X1  g064(.A(G2105), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT65), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n464), .A2(new_n491), .A3(KEYINPUT4), .A4(G138), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n465), .A2(G102), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n486), .A2(new_n490), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G164));
  INV_X1    g070(.A(G543), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT5), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(KEYINPUT66), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT66), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(KEYINPUT5), .A3(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n501), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT6), .B(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G88), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G50), .ZN(new_n509));
  OAI22_X1  g084(.A1(new_n506), .A2(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n504), .A2(new_n510), .ZN(G166));
  AND3_X1   g086(.A1(new_n499), .A2(KEYINPUT5), .A3(G543), .ZN(new_n512));
  AOI21_X1  g087(.A(G543), .B1(new_n499), .B2(KEYINPUT5), .ZN(new_n513));
  OAI211_X1 g088(.A(G63), .B(G651), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT67), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT67), .ZN(new_n516));
  NAND4_X1  g091(.A1(new_n501), .A2(new_n516), .A3(G63), .A4(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n501), .A2(G89), .A3(new_n505), .ZN(new_n521));
  OR2_X1    g096(.A1(KEYINPUT68), .A2(G51), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT68), .A2(G51), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n505), .A2(G543), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n518), .A2(new_n520), .A3(new_n525), .ZN(G286));
  INV_X1    g101(.A(G286), .ZN(G168));
  INV_X1    g102(.A(KEYINPUT69), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n501), .A2(G64), .ZN(new_n529));
  NAND2_X1  g104(.A1(G77), .A2(G543), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n503), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n501), .A2(G90), .A3(new_n505), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n505), .A2(G52), .A3(G543), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n528), .B1(new_n531), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n536), .B1(new_n498), .B2(new_n500), .ZN(new_n537));
  INV_X1    g112(.A(new_n530), .ZN(new_n538));
  OAI21_X1  g113(.A(G651), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n539), .A2(KEYINPUT69), .A3(new_n533), .A4(new_n532), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n535), .A2(new_n540), .ZN(G171));
  AOI22_X1  g116(.A1(new_n501), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n503), .ZN(new_n543));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  INV_X1    g119(.A(G43), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n506), .A2(new_n544), .B1(new_n508), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT70), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n549), .A2(new_n553), .ZN(G188));
  INV_X1    g129(.A(G53), .ZN(new_n555));
  OAI21_X1  g130(.A(KEYINPUT9), .B1(new_n508), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n505), .A2(new_n557), .A3(G53), .A4(G543), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n560), .B1(new_n498), .B2(new_n500), .ZN(new_n561));
  AND2_X1   g136(.A1(G78), .A2(G543), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n506), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G91), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n559), .A2(new_n563), .A3(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  INV_X1    g142(.A(G166), .ZN(G303));
  NAND2_X1  g143(.A1(new_n564), .A2(G87), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n501), .B2(G74), .ZN(new_n570));
  INV_X1    g145(.A(new_n508), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G49), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(G288));
  AND2_X1   g148(.A1(G73), .A2(G543), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n501), .B2(G61), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n575), .A2(new_n503), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n564), .A2(G86), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n571), .A2(G48), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(G305));
  NOR2_X1   g154(.A1(new_n512), .A2(new_n513), .ZN(new_n580));
  INV_X1    g155(.A(G60), .ZN(new_n581));
  INV_X1    g156(.A(G72), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n580), .A2(new_n581), .B1(new_n582), .B2(new_n496), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT71), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI221_X1 g160(.A(KEYINPUT71), .B1(new_n582), .B2(new_n496), .C1(new_n580), .C2(new_n581), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n585), .A2(G651), .A3(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(G85), .ZN(new_n588));
  INV_X1    g163(.A(G47), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n506), .A2(new_n588), .B1(new_n508), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT72), .ZN(new_n591));
  AND2_X1   g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n590), .A2(new_n591), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n587), .B1(new_n592), .B2(new_n593), .ZN(G290));
  AND3_X1   g169(.A1(new_n501), .A2(G92), .A3(new_n505), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT10), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n508), .A2(KEYINPUT73), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n508), .A2(KEYINPUT73), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n597), .A2(G54), .A3(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n501), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n600), .A2(new_n503), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n596), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(new_n603), .B2(G171), .ZN(G321));
  XOR2_X1   g180(.A(G321), .B(KEYINPUT74), .Z(G284));
  NAND2_X1  g181(.A1(G299), .A2(new_n603), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G168), .B2(new_n603), .ZN(G297));
  OAI21_X1  g183(.A(new_n607), .B1(G168), .B2(new_n603), .ZN(G280));
  INV_X1    g184(.A(new_n602), .ZN(new_n610));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G860), .ZN(G148));
  INV_X1    g187(.A(new_n547), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(new_n603), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n602), .A2(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(new_n603), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n477), .A2(G123), .ZN(new_n618));
  OR2_X1    g193(.A1(G99), .A2(G2105), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n619), .B(G2104), .C1(G111), .C2(new_n476), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(G135), .B2(new_n464), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2096), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n476), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n627), .A2(G2100), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(G2100), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n623), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT75), .ZN(G156));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT77), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(KEYINPUT14), .ZN(new_n637));
  XOR2_X1   g212(.A(G2451), .B(G2454), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT76), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n636), .A2(KEYINPUT14), .A3(new_n640), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n642), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT78), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n644), .B1(new_n642), .B2(new_n645), .ZN(new_n651));
  OR3_X1    g226(.A1(new_n647), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n650), .B1(new_n647), .B2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(G14), .A3(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(G401));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2067), .B(G2678), .Z(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(new_n660), .A3(KEYINPUT17), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT18), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n659), .B2(KEYINPUT18), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n663), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2096), .B(G2100), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1956), .B(G2474), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT79), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1961), .B(G1966), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT80), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n672), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n673), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n674), .A2(new_n676), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n670), .A2(new_n672), .A3(KEYINPUT20), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n673), .A2(new_n679), .ZN(new_n680));
  OAI221_X1 g255(.A(new_n677), .B1(KEYINPUT20), .B2(new_n678), .C1(new_n680), .C2(new_n676), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT82), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1991), .B(G1996), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT81), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n686), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G229));
  NOR2_X1   g265(.A1(G16), .A2(G24), .ZN(new_n691));
  XOR2_X1   g266(.A(G290), .B(KEYINPUT85), .Z(new_n692));
  AOI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(G16), .ZN(new_n693));
  INV_X1    g268(.A(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G29), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n696), .A2(G25), .ZN(new_n697));
  OAI21_X1  g272(.A(G2104), .B1(new_n476), .B2(G107), .ZN(new_n698));
  INV_X1    g273(.A(G95), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(new_n476), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT84), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n464), .A2(G131), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n477), .A2(G119), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n697), .B1(new_n704), .B2(G29), .ZN(new_n705));
  MUX2_X1   g280(.A(new_n697), .B(new_n705), .S(KEYINPUT83), .Z(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT35), .B(G1991), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT87), .ZN(new_n709));
  AOI22_X1  g284(.A1(new_n707), .A2(new_n708), .B1(new_n709), .B2(KEYINPUT36), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n695), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n707), .A2(new_n708), .ZN(new_n712));
  MUX2_X1   g287(.A(G6), .B(G305), .S(G16), .Z(new_n713));
  XOR2_X1   g288(.A(KEYINPUT32), .B(G1981), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G22), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G166), .B2(new_n716), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(G1971), .Z(new_n719));
  NAND2_X1  g294(.A1(new_n716), .A2(G23), .ZN(new_n720));
  INV_X1    g295(.A(G288), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(new_n716), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT33), .B(G1976), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT86), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n722), .B(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n715), .A2(new_n719), .A3(new_n725), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT34), .Z(new_n727));
  NAND3_X1  g302(.A1(new_n711), .A2(new_n712), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n709), .A2(KEYINPUT36), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n622), .A2(G29), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT93), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT30), .B(G28), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n732), .B1(new_n696), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT31), .B(G11), .ZN(new_n735));
  OR2_X1    g310(.A1(KEYINPUT24), .A2(G34), .ZN(new_n736));
  NAND2_X1  g311(.A1(KEYINPUT24), .A2(G34), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n736), .A2(new_n696), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G160), .B2(new_n696), .ZN(new_n739));
  INV_X1    g314(.A(G2084), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n734), .A2(new_n735), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(G115), .A2(G2104), .ZN(new_n743));
  INV_X1    g318(.A(G127), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n475), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G2105), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT90), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n464), .A2(G139), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n465), .A2(G103), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT25), .Z(new_n750));
  NAND3_X1  g325(.A1(new_n747), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  MUX2_X1   g326(.A(G33), .B(new_n751), .S(G29), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G2072), .ZN(new_n753));
  NAND2_X1  g328(.A1(G168), .A2(G16), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT92), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G16), .B2(G21), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(KEYINPUT92), .B2(new_n754), .ZN(new_n758));
  INV_X1    g333(.A(G1966), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NOR3_X1   g335(.A1(new_n742), .A2(new_n753), .A3(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(G29), .A2(G32), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n477), .A2(G129), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n465), .A2(G105), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G141), .B2(new_n464), .ZN(new_n766));
  NAND3_X1  g341(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT91), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT26), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n762), .B1(new_n771), .B2(G29), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT27), .B(G1996), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n696), .A2(G27), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G164), .B2(new_n696), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT95), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT94), .B(G2078), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n777), .A2(new_n779), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n716), .A2(G5), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G171), .B2(new_n716), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n783), .A2(G1961), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n783), .A2(G1961), .ZN(new_n785));
  NOR4_X1   g360(.A1(new_n780), .A2(new_n781), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n761), .A2(new_n774), .A3(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT96), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n696), .A2(G26), .ZN(new_n790));
  OAI21_X1  g365(.A(G2104), .B1(new_n476), .B2(G116), .ZN(new_n791));
  INV_X1    g366(.A(G104), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(new_n476), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT88), .Z(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G128), .B2(new_n477), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n464), .A2(G140), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n790), .B1(new_n797), .B2(G29), .ZN(new_n798));
  MUX2_X1   g373(.A(new_n790), .B(new_n798), .S(KEYINPUT28), .Z(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT89), .B(G2067), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n716), .A2(G4), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n610), .B2(new_n716), .ZN(new_n803));
  INV_X1    g378(.A(G1348), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n716), .A2(G19), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n547), .B2(new_n716), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(G1341), .Z(new_n808));
  NAND2_X1  g383(.A1(new_n716), .A2(G20), .ZN(new_n809));
  INV_X1    g384(.A(G299), .ZN(new_n810));
  OAI211_X1 g385(.A(KEYINPUT23), .B(new_n809), .C1(new_n810), .C2(new_n716), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(KEYINPUT23), .B2(new_n809), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1956), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n801), .A2(new_n805), .A3(new_n808), .A4(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n787), .B2(new_n788), .ZN(new_n815));
  AND3_X1   g390(.A1(new_n730), .A2(new_n789), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n696), .A2(G35), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G162), .B2(new_n696), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT29), .B(G2090), .Z(new_n819));
  XOR2_X1   g394(.A(new_n818), .B(new_n819), .Z(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n729), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n711), .A2(new_n822), .A3(new_n712), .A4(new_n727), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n816), .A2(KEYINPUT97), .A3(new_n821), .A4(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT97), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n730), .A2(new_n789), .A3(new_n823), .A4(new_n815), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(new_n820), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n824), .A2(new_n827), .ZN(G311));
  NAND3_X1  g403(.A1(new_n816), .A2(new_n821), .A3(new_n823), .ZN(G150));
  NAND2_X1  g404(.A1(G80), .A2(G543), .ZN(new_n830));
  INV_X1    g405(.A(G67), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n580), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(G651), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n501), .A2(G93), .A3(new_n505), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n505), .A2(G55), .A3(G543), .ZN(new_n835));
  AND3_X1   g410(.A1(new_n834), .A2(KEYINPUT98), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(KEYINPUT98), .B1(new_n834), .B2(new_n835), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n833), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(G860), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT100), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT37), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n602), .A2(new_n611), .ZN(new_n842));
  XNOR2_X1  g417(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT99), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n834), .A2(new_n835), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT98), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n834), .A2(KEYINPUT98), .A3(new_n835), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n845), .B1(new_n850), .B2(new_n833), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n833), .B(new_n845), .C1(new_n836), .C2(new_n837), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n613), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n838), .A2(KEYINPUT99), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n855), .A2(new_n547), .A3(new_n852), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n844), .B(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n841), .B1(new_n858), .B2(G860), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT101), .Z(G145));
  NAND2_X1  g435(.A1(new_n751), .A2(KEYINPUT102), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n770), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n625), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n622), .B(new_n471), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(new_n704), .Z(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n863), .A2(new_n866), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n797), .B(G164), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n464), .A2(G142), .ZN(new_n871));
  AOI22_X1  g446(.A1(KEYINPUT103), .A2(new_n871), .B1(new_n477), .B2(G130), .ZN(new_n872));
  NOR2_X1   g447(.A1(G106), .A2(G2105), .ZN(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(new_n476), .B2(G118), .ZN(new_n874));
  OAI221_X1 g449(.A(new_n872), .B1(KEYINPUT103), .B2(new_n871), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(G162), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n870), .B(new_n876), .Z(new_n877));
  OR2_X1    g452(.A1(new_n869), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(G37), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n869), .A2(new_n877), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g457(.A(new_n857), .B(new_n615), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n610), .A2(G299), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n602), .A2(new_n810), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT41), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n884), .A2(KEYINPUT41), .A3(new_n885), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n883), .A2(new_n890), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n891), .B(KEYINPUT105), .Z(new_n892));
  INV_X1    g467(.A(new_n886), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n883), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT104), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n587), .B(G288), .C1(new_n592), .C2(new_n593), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n590), .B(new_n591), .ZN(new_n898));
  AOI21_X1  g473(.A(G288), .B1(new_n898), .B2(new_n587), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT106), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n576), .A2(new_n901), .A3(new_n577), .A4(new_n578), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n575), .A2(new_n503), .ZN(new_n903));
  INV_X1    g478(.A(G86), .ZN(new_n904));
  INV_X1    g479(.A(G48), .ZN(new_n905));
  OAI22_X1  g480(.A1(new_n506), .A2(new_n904), .B1(new_n508), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(KEYINPUT106), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(G166), .B1(new_n902), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n902), .A2(new_n907), .A3(G166), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT108), .B1(new_n900), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(G290), .A2(new_n721), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n896), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT108), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n914), .A2(new_n915), .A3(new_n910), .A4(new_n909), .ZN(new_n916));
  INV_X1    g491(.A(new_n910), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n913), .B(new_n896), .C1(new_n917), .C2(new_n908), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT107), .B1(new_n900), .B2(new_n911), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n912), .B(new_n916), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT42), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n892), .A2(new_n895), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n923), .B1(new_n892), .B2(new_n895), .ZN(new_n925));
  OAI21_X1  g500(.A(G868), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n838), .A2(new_n603), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(G295));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n927), .ZN(G331));
  NAND2_X1  g504(.A1(G286), .A2(KEYINPUT110), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT110), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n518), .A2(new_n525), .A3(new_n931), .A4(new_n520), .ZN(new_n932));
  NAND3_X1  g507(.A1(G301), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n521), .A2(new_n524), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n934), .B1(new_n515), .B2(new_n517), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n931), .B1(new_n935), .B2(new_n520), .ZN(new_n936));
  AND4_X1   g511(.A1(new_n931), .A2(new_n518), .A3(new_n520), .A4(new_n525), .ZN(new_n937));
  OAI21_X1  g512(.A(G171), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n855), .A2(new_n547), .A3(new_n852), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n547), .B1(new_n855), .B2(new_n852), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n933), .B(new_n938), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n936), .A2(new_n937), .A3(G171), .ZN(new_n942));
  AOI22_X1  g517(.A1(new_n930), .A2(new_n932), .B1(new_n540), .B2(new_n535), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n856), .B(new_n854), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n941), .A2(new_n944), .A3(KEYINPUT111), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT111), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n857), .A2(new_n946), .A3(new_n933), .A4(new_n938), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n886), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n941), .A2(new_n944), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n890), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n922), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n945), .A2(new_n890), .A3(new_n947), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n941), .A2(new_n944), .A3(new_n886), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n953), .A2(new_n922), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT112), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n922), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n893), .B1(new_n945), .B2(new_n947), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n890), .A2(new_n950), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n963));
  AOI21_X1  g538(.A(G37), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n956), .A2(new_n958), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n922), .B1(new_n953), .B2(new_n954), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n955), .A2(new_n966), .A3(G37), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n965), .B1(new_n958), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n879), .B1(new_n952), .B2(KEYINPUT112), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n953), .A2(new_n922), .A3(new_n954), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n963), .B1(new_n962), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT113), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT113), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n956), .A2(new_n975), .A3(new_n964), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n974), .A2(KEYINPUT43), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n969), .B1(new_n967), .B2(new_n958), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n977), .A2(KEYINPUT114), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT114), .B1(new_n977), .B2(new_n978), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n970), .B1(new_n979), .B2(new_n980), .ZN(G397));
  INV_X1    g556(.A(KEYINPUT124), .ZN(new_n982));
  INV_X1    g557(.A(G1384), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n494), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT50), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n466), .A2(new_n470), .A3(G40), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT116), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n466), .A2(new_n470), .A3(KEYINPUT116), .A4(G40), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n494), .A2(new_n991), .A3(new_n983), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n985), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n984), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n494), .A2(KEYINPUT45), .A3(new_n983), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(new_n990), .A3(new_n997), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n994), .A2(new_n740), .B1(new_n998), .B2(new_n759), .ZN(new_n999));
  NAND2_X1  g574(.A1(G286), .A2(G8), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n1002));
  INV_X1    g577(.A(G8), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n1002), .B(new_n1000), .C1(new_n999), .C2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n998), .ZN(new_n1005));
  OAI22_X1  g580(.A1(new_n1005), .A2(G1966), .B1(G2084), .B2(new_n993), .ZN(new_n1006));
  OAI211_X1 g581(.A(KEYINPUT51), .B(G8), .C1(new_n1006), .C2(G286), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1001), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n494), .A2(new_n983), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1003), .B1(new_n990), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n721), .A2(G1976), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT52), .ZN(new_n1013));
  OR3_X1    g588(.A1(new_n903), .A2(new_n906), .A3(G1981), .ZN(new_n1014));
  OAI21_X1  g589(.A(G1981), .B1(new_n903), .B2(new_n906), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT49), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1014), .A2(new_n1015), .A3(KEYINPUT49), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(new_n1010), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1976), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT52), .B1(G288), .B2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1010), .A2(new_n1011), .A3(new_n1022), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n1013), .A2(new_n1020), .A3(new_n1023), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n494), .A2(new_n991), .A3(new_n983), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n991), .B1(new_n494), .B2(new_n983), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G2090), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(new_n1028), .A3(new_n990), .ZN(new_n1029));
  XOR2_X1   g604(.A(KEYINPUT117), .B(G1971), .Z(new_n1030));
  NAND2_X1  g605(.A1(new_n998), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1003), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(G166), .A2(new_n1003), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1033), .B(KEYINPUT55), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n993), .A2(KEYINPUT119), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT119), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n985), .A2(new_n1037), .A3(new_n990), .A4(new_n992), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1036), .A2(new_n1028), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1003), .B1(new_n1039), .B2(new_n1031), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1024), .B(new_n1035), .C1(new_n1040), .C2(new_n1034), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1008), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT121), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n993), .A2(new_n1043), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n985), .A2(KEYINPUT121), .A3(new_n990), .A4(new_n992), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G1961), .ZN(new_n1047));
  INV_X1    g622(.A(G2078), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1005), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n1050));
  AOI22_X1  g625(.A1(new_n1046), .A2(new_n1047), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1005), .A2(KEYINPUT53), .A3(new_n1048), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1051), .A2(KEYINPUT123), .A3(G301), .A4(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT121), .B1(new_n1027), .B2(new_n990), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1045), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1047), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1050), .B1(new_n998), .B2(G2078), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1056), .A2(G301), .A3(new_n1057), .A4(new_n1052), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT123), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n1009), .A2(KEYINPUT115), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1009), .A2(KEYINPUT115), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(new_n995), .A3(new_n1062), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n997), .A2(KEYINPUT53), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n986), .A2(G2078), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1056), .A2(new_n1066), .A3(new_n1057), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(G171), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1053), .A2(new_n1060), .A3(KEYINPUT54), .A4(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n1070));
  AOI21_X1  g645(.A(G301), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1071));
  AND4_X1   g646(.A1(G301), .A2(new_n1056), .A3(new_n1057), .A4(new_n1066), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1042), .A2(new_n1069), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1956), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n993), .A2(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT56), .B(G2072), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n996), .A2(new_n990), .A3(new_n997), .A4(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(G299), .A2(KEYINPUT120), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n559), .A2(new_n565), .A3(new_n1081), .A4(new_n563), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1080), .A2(KEYINPUT57), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT57), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1079), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G2067), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n990), .A2(new_n1009), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1089), .B1(new_n1046), .B2(new_n804), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1086), .B1(new_n1090), .B2(new_n602), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1076), .B(new_n1078), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1046), .A2(new_n804), .ZN(new_n1094));
  OR2_X1    g669(.A1(new_n602), .A2(KEYINPUT122), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1094), .A2(KEYINPUT60), .A3(new_n1088), .A4(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n602), .A2(KEYINPUT122), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1090), .A2(KEYINPUT60), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1090), .A2(KEYINPUT60), .A3(new_n1095), .A4(new_n1097), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1086), .A2(KEYINPUT61), .A3(new_n1092), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT61), .B1(new_n1086), .B2(new_n1092), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n984), .B1(new_n988), .B2(new_n989), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT58), .B(G1341), .ZN(new_n1106));
  OAI22_X1  g681(.A1(new_n998), .A2(G1996), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT59), .B1(new_n1107), .B2(new_n547), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1103), .A2(new_n1104), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1107), .A2(KEYINPUT59), .A3(new_n547), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1102), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1074), .B1(new_n1093), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1113));
  NOR2_X1   g688(.A1(G288), .A2(G1976), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1114), .B(KEYINPUT118), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  AOI211_X1 g691(.A(new_n1003), .B(new_n1105), .C1(new_n1116), .C2(new_n1014), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT63), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1006), .A2(G8), .A3(G168), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1118), .B1(new_n1041), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1024), .A2(new_n1035), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT63), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1122));
  OR3_X1    g697(.A1(new_n1121), .A2(new_n1119), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1117), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1024), .A2(new_n1034), .A3(new_n1032), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n982), .B1(new_n1112), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1041), .B1(new_n1008), .B2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1129), .B(new_n1071), .C1(new_n1128), .C2(new_n1008), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1125), .ZN(new_n1131));
  AOI211_X1 g706(.A(new_n1131), .B(new_n1117), .C1(new_n1120), .C2(new_n1123), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1111), .A2(new_n1093), .ZN(new_n1133));
  OAI211_X1 g708(.A(KEYINPUT124), .B(new_n1132), .C1(new_n1133), .C2(new_n1074), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1127), .A2(new_n1130), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1063), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n990), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n797), .B(new_n1087), .ZN(new_n1139));
  XOR2_X1   g714(.A(new_n770), .B(G1996), .Z(new_n1140));
  AND2_X1   g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n704), .A2(new_n708), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n704), .A2(new_n708), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(G290), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1145), .B1(new_n694), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n694), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1138), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1135), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1137), .B1(new_n1139), .B2(new_n771), .ZN(new_n1152));
  XOR2_X1   g727(.A(new_n1152), .B(KEYINPUT126), .Z(new_n1153));
  NOR2_X1   g728(.A1(new_n1137), .A2(G1996), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT46), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1156), .B(KEYINPUT47), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1137), .A2(new_n1148), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1158), .B(KEYINPUT48), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1159), .B1(new_n1144), .B2(new_n1138), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1143), .B(KEYINPUT125), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1141), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n795), .A2(new_n1087), .A3(new_n796), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1137), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1157), .A2(new_n1160), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1151), .A2(new_n1165), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g741(.A(G227), .ZN(new_n1168));
  NAND3_X1  g742(.A1(new_n654), .A2(G319), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n1170));
  OAI21_X1  g744(.A(new_n689), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g745(.A(new_n1171), .B1(new_n1170), .B2(new_n1169), .ZN(new_n1172));
  NAND3_X1  g746(.A1(new_n1172), .A2(new_n881), .A3(new_n968), .ZN(G225));
  INV_X1    g747(.A(G225), .ZN(G308));
endmodule


