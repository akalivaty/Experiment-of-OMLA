//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 0 0 1 1 1 0 1 0 0 1 1 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n446, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n568, new_n570, new_n571,
    new_n572, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n586, new_n587,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n631, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1277, new_n1278, new_n1279, new_n1280;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT66), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT67), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT68), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT69), .Z(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  OR2_X1    g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(KEYINPUT70), .A3(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n466), .A2(new_n470), .A3(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n463), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT3), .B(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G137), .ZN(new_n475));
  NAND2_X1  g050(.A1(G101), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(G2105), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n473), .A2(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(new_n468), .A2(new_n469), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n479), .A2(new_n463), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  INV_X1    g062(.A(G2104), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G102), .ZN(new_n490));
  AOI22_X1  g065(.A1(new_n474), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(new_n463), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  OAI211_X1 g068(.A(G138), .B(new_n463), .C1(new_n468), .C2(new_n469), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n463), .A2(G138), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n474), .A2(KEYINPUT71), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  OR2_X1    g075(.A1(KEYINPUT72), .A2(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT72), .A2(KEYINPUT4), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n497), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(new_n470), .A3(new_n466), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n492), .B1(new_n500), .B2(new_n504), .ZN(G164));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT6), .B(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n512), .A2(KEYINPUT6), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  OAI211_X1 g096(.A(new_n517), .B(new_n519), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT73), .B(G88), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n515), .A2(new_n516), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n513), .A2(new_n524), .ZN(G166));
  NAND3_X1  g100(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n526));
  INV_X1    g101(.A(G51), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n515), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  INV_X1    g105(.A(G89), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n531), .B2(new_n522), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n528), .A2(new_n532), .ZN(G168));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n515), .A2(new_n534), .B1(new_n522), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n520), .A2(new_n521), .ZN(new_n537));
  INV_X1    g112(.A(G64), .ZN(new_n538));
  INV_X1    g113(.A(G77), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n537), .A2(new_n538), .B1(new_n539), .B2(new_n507), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(KEYINPUT74), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT74), .ZN(new_n542));
  OAI221_X1 g117(.A(new_n542), .B1(new_n539), .B2(new_n507), .C1(new_n537), .C2(new_n538), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n541), .A2(G651), .A3(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g121(.A1(new_n541), .A2(KEYINPUT75), .A3(new_n543), .A4(G651), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n536), .B1(new_n546), .B2(new_n547), .ZN(G171));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n537), .A2(new_n549), .ZN(new_n550));
  AND2_X1   g125(.A1(G68), .A2(G543), .ZN(new_n551));
  OAI21_X1  g126(.A(G651), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(KEYINPUT76), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT76), .ZN(new_n554));
  OAI211_X1 g129(.A(new_n554), .B(G651), .C1(new_n550), .C2(new_n551), .ZN(new_n555));
  INV_X1    g130(.A(G43), .ZN(new_n556));
  XNOR2_X1  g131(.A(KEYINPUT77), .B(G81), .ZN(new_n557));
  OAI22_X1  g132(.A1(new_n515), .A2(new_n556), .B1(new_n522), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n553), .A2(new_n555), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(KEYINPUT78), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n558), .B1(new_n552), .B2(KEYINPUT76), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT78), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n562), .A2(new_n563), .A3(new_n555), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n568));
  XOR2_X1   g143(.A(new_n568), .B(KEYINPUT79), .Z(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(new_n572));
  XOR2_X1   g147(.A(new_n572), .B(KEYINPUT80), .Z(G188));
  NAND2_X1  g148(.A1(new_n522), .A2(KEYINPUT81), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT81), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n510), .A2(new_n514), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(G91), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n514), .A2(G53), .A3(G543), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT9), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n510), .A2(KEYINPUT82), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT82), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n537), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n583), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n584));
  OAI211_X1 g159(.A(new_n577), .B(new_n579), .C1(new_n584), .C2(new_n512), .ZN(G299));
  NAND2_X1  g160(.A1(new_n546), .A2(new_n547), .ZN(new_n586));
  INV_X1    g161(.A(new_n536), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G301));
  INV_X1    g163(.A(G168), .ZN(G286));
  INV_X1    g164(.A(G166), .ZN(G303));
  INV_X1    g165(.A(G74), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n512), .B1(new_n537), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n515), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n592), .B1(new_n593), .B2(G49), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n574), .A2(G87), .A3(new_n576), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(G288));
  OAI21_X1  g171(.A(G61), .B1(new_n520), .B2(new_n521), .ZN(new_n597));
  NAND2_X1  g172(.A1(G73), .A2(G543), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n512), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AND2_X1   g174(.A1(G48), .A2(G543), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n599), .B1(new_n514), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n574), .A2(G86), .A3(new_n576), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(G305));
  AOI22_X1  g178(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(new_n512), .ZN(new_n605));
  INV_X1    g180(.A(G47), .ZN(new_n606));
  INV_X1    g181(.A(G85), .ZN(new_n607));
  OAI22_X1  g182(.A1(new_n515), .A2(new_n606), .B1(new_n522), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(G290));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NOR2_X1   g186(.A1(G301), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n574), .A2(G92), .A3(new_n576), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g190(.A1(new_n574), .A2(new_n576), .A3(KEYINPUT10), .A4(G92), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AND3_X1   g192(.A1(new_n514), .A2(G54), .A3(G543), .ZN(new_n618));
  NOR3_X1   g193(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT82), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n581), .B1(new_n508), .B2(new_n509), .ZN(new_n620));
  OAI21_X1  g195(.A(G66), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(G79), .A2(G543), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n618), .B1(new_n623), .B2(G651), .ZN(new_n624));
  AND3_X1   g199(.A1(new_n617), .A2(new_n624), .A3(KEYINPUT83), .ZN(new_n625));
  AOI21_X1  g200(.A(KEYINPUT83), .B1(new_n617), .B2(new_n624), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n612), .B1(new_n611), .B2(new_n627), .ZN(G284));
  AOI21_X1  g203(.A(new_n612), .B1(new_n611), .B2(new_n627), .ZN(G321));
  NAND2_X1  g204(.A1(G286), .A2(G868), .ZN(new_n630));
  INV_X1    g205(.A(G299), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(G868), .ZN(G297));
  OAI21_X1  g207(.A(new_n630), .B1(new_n631), .B2(G868), .ZN(G280));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n627), .B1(new_n634), .B2(G860), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT84), .Z(G148));
  NAND2_X1  g211(.A1(new_n566), .A2(new_n611), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n617), .A2(new_n624), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT83), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n617), .A2(new_n624), .A3(KEYINPUT83), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(new_n634), .A3(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n637), .B1(new_n642), .B2(new_n611), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT11), .Z(G282));
  INV_X1    g219(.A(new_n643), .ZN(G323));
  AND2_X1   g220(.A1(new_n466), .A2(new_n470), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(new_n489), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(KEYINPUT12), .ZN(new_n648));
  INV_X1    g223(.A(KEYINPUT12), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n646), .A2(new_n649), .A3(new_n489), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT13), .ZN(new_n652));
  INV_X1    g227(.A(G2100), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT85), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n480), .A2(G135), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n482), .A2(G123), .ZN(new_n657));
  NOR2_X1   g232(.A1(G99), .A2(G2105), .ZN(new_n658));
  OAI21_X1  g233(.A(G2104), .B1(new_n463), .B2(G111), .ZN(new_n659));
  OAI211_X1 g234(.A(new_n656), .B(new_n657), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2096), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n652), .B2(new_n653), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n655), .A2(new_n662), .ZN(G156));
  XOR2_X1   g238(.A(G2443), .B(G2446), .Z(new_n664));
  XNOR2_X1  g239(.A(G2451), .B(G2454), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(KEYINPUT15), .B(G2435), .Z(new_n670));
  INV_X1    g245(.A(G2438), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT15), .B(G2435), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(G2438), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2427), .B(G2430), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n677), .A2(KEYINPUT87), .A3(KEYINPUT14), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT87), .ZN(new_n679));
  INV_X1    g254(.A(new_n676), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n672), .B2(new_n674), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT14), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n679), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n672), .A2(new_n674), .A3(new_n680), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1341), .B(G1348), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT88), .ZN(new_n687));
  AND3_X1   g262(.A1(new_n684), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n687), .B1(new_n684), .B2(new_n685), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n669), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n684), .A2(new_n685), .ZN(new_n691));
  INV_X1    g266(.A(new_n687), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n684), .A2(new_n685), .A3(new_n687), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n693), .A2(new_n668), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n690), .A2(new_n695), .A3(G14), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT89), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g273(.A1(new_n690), .A2(new_n695), .A3(KEYINPUT89), .A4(G14), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n698), .A2(new_n700), .ZN(G401));
  XOR2_X1   g276(.A(G2084), .B(G2090), .Z(new_n702));
  XNOR2_X1  g277(.A(G2067), .B(G2678), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n702), .ZN(new_n705));
  XOR2_X1   g280(.A(G2072), .B(G2078), .Z(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(KEYINPUT17), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n702), .A2(new_n703), .ZN(new_n709));
  OAI221_X1 g284(.A(new_n704), .B1(new_n703), .B2(new_n707), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n704), .A2(new_n706), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT18), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(G2096), .B(G2100), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT90), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n713), .B(new_n715), .ZN(G227));
  XOR2_X1   g291(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n717));
  XNOR2_X1  g292(.A(G1956), .B(G2474), .ZN(new_n718));
  XNOR2_X1  g293(.A(G1961), .B(G1966), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(G1971), .B(G1976), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT19), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT20), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n718), .B(new_n719), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n728), .A2(new_n724), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n724), .A2(new_n718), .A3(new_n719), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR3_X1   g306(.A1(new_n727), .A2(G1986), .A3(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G1986), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n725), .B(KEYINPUT20), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n729), .A2(new_n730), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n717), .B1(new_n732), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(G1991), .B(G1996), .ZN(new_n738));
  INV_X1    g313(.A(G1981), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(G1986), .B1(new_n727), .B2(new_n731), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n734), .A2(new_n735), .A3(new_n733), .ZN(new_n742));
  INV_X1    g317(.A(new_n717), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  AND3_X1   g319(.A1(new_n737), .A2(new_n740), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n740), .B1(new_n737), .B2(new_n744), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n745), .A2(new_n746), .ZN(G229));
  MUX2_X1   g322(.A(G6), .B(G305), .S(G16), .Z(new_n748));
  XOR2_X1   g323(.A(KEYINPUT32), .B(G1981), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(G16), .A2(G23), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT91), .ZN(new_n752));
  INV_X1    g327(.A(G16), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(G288), .B2(new_n753), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT33), .B(G1976), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT92), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n754), .A2(new_n756), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n753), .A2(G22), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G166), .B2(new_n753), .ZN(new_n760));
  INV_X1    g335(.A(G1971), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n750), .A2(new_n757), .A3(new_n758), .A4(new_n762), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(KEYINPUT34), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(KEYINPUT34), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n753), .A2(G24), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n609), .B2(new_n753), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(new_n733), .ZN(new_n768));
  INV_X1    g343(.A(G29), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G25), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n480), .A2(G131), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n482), .A2(G119), .ZN(new_n772));
  OR2_X1    g347(.A1(G95), .A2(G2105), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n773), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n771), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n770), .B1(new_n776), .B2(new_n769), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT35), .B(G1991), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n764), .A2(new_n765), .A3(new_n768), .A4(new_n779), .ZN(new_n780));
  OR3_X1    g355(.A1(new_n780), .A2(KEYINPUT93), .A3(KEYINPUT36), .ZN(new_n781));
  OAI21_X1  g356(.A(KEYINPUT93), .B1(new_n780), .B2(KEYINPUT36), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n780), .A2(KEYINPUT36), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n769), .A2(G35), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G162), .B2(new_n769), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT29), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G2090), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n753), .A2(G19), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n565), .B2(G16), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n791), .A2(G1341), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n769), .A2(G33), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT25), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n480), .A2(G139), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n646), .A2(G127), .ZN(new_n798));
  INV_X1    g373(.A(G115), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(new_n488), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n797), .B1(new_n800), .B2(G2105), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n793), .B1(new_n801), .B2(new_n769), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G2072), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n788), .A2(new_n792), .A3(new_n803), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n769), .A2(G32), .ZN(new_n805));
  NAND3_X1  g380(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT26), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G129), .B2(new_n482), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n480), .A2(G141), .B1(G105), .B2(new_n489), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n805), .B1(new_n810), .B2(G29), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT27), .B(G1996), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT24), .ZN(new_n814));
  INV_X1    g389(.A(G34), .ZN(new_n815));
  AOI21_X1  g390(.A(G29), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n814), .B2(new_n815), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G160), .B2(new_n769), .ZN(new_n818));
  NOR2_X1   g393(.A1(G5), .A2(G16), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT99), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G171), .B2(G16), .ZN(new_n821));
  OAI221_X1 g396(.A(new_n813), .B1(G2084), .B2(new_n818), .C1(new_n821), .C2(G1961), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT100), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n791), .A2(G1341), .B1(G1961), .B2(new_n821), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n804), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n627), .A2(new_n753), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(G4), .B2(new_n753), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT94), .B(G1348), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n811), .A2(new_n812), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT97), .Z(new_n832));
  NAND2_X1  g407(.A1(new_n769), .A2(G27), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT101), .Z(new_n834));
  AOI21_X1  g409(.A(new_n497), .B1(new_n464), .B2(new_n465), .ZN(new_n835));
  OAI21_X1  g410(.A(KEYINPUT4), .B1(new_n835), .B2(KEYINPUT71), .ZN(new_n836));
  INV_X1    g411(.A(new_n499), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n504), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(G114), .A2(G2104), .ZN(new_n839));
  INV_X1    g414(.A(G126), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n479), .B2(new_n840), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n841), .A2(G2105), .B1(G102), .B2(new_n489), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n834), .B1(new_n843), .B2(G29), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(G2078), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n753), .A2(G21), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(G168), .B2(new_n753), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n847), .A2(G1966), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT98), .ZN(new_n849));
  NOR3_X1   g424(.A1(new_n832), .A2(new_n845), .A3(new_n849), .ZN(new_n850));
  XOR2_X1   g425(.A(KEYINPUT96), .B(KEYINPUT28), .Z(new_n851));
  NAND2_X1  g426(.A1(new_n769), .A2(G26), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  AOI22_X1  g428(.A1(G128), .A2(new_n482), .B1(new_n480), .B2(G140), .ZN(new_n854));
  OAI21_X1  g429(.A(G2104), .B1(new_n463), .B2(G116), .ZN(new_n855));
  NOR2_X1   g430(.A1(G104), .A2(G2105), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT95), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n853), .B1(new_n860), .B2(new_n769), .ZN(new_n861));
  INV_X1    g436(.A(G2067), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(G28), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n864), .A2(KEYINPUT30), .ZN(new_n865));
  AOI21_X1  g440(.A(G29), .B1(new_n864), .B2(KEYINPUT30), .ZN(new_n866));
  OR2_X1    g441(.A1(KEYINPUT31), .A2(G11), .ZN(new_n867));
  NAND2_X1  g442(.A1(KEYINPUT31), .A2(G11), .ZN(new_n868));
  AOI22_X1  g443(.A1(new_n865), .A2(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(new_n660), .B2(new_n769), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n870), .B1(new_n847), .B2(G1966), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n863), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n872), .B1(G2084), .B2(new_n818), .ZN(new_n873));
  XOR2_X1   g448(.A(KEYINPUT102), .B(KEYINPUT23), .Z(new_n874));
  NAND2_X1  g449(.A1(new_n753), .A2(G20), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(new_n631), .B2(new_n753), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n877), .B(G1956), .Z(new_n878));
  NAND4_X1  g453(.A1(new_n830), .A2(new_n850), .A3(new_n873), .A4(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n828), .A2(new_n829), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n822), .A2(new_n823), .ZN(new_n881));
  NOR4_X1   g456(.A1(new_n826), .A2(new_n879), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n784), .A2(new_n882), .ZN(G150));
  INV_X1    g458(.A(G150), .ZN(G311));
  INV_X1    g459(.A(KEYINPUT39), .ZN(new_n885));
  AOI22_X1  g460(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n886), .A2(new_n512), .ZN(new_n887));
  XNOR2_X1  g462(.A(KEYINPUT103), .B(G55), .ZN(new_n888));
  INV_X1    g463(.A(G93), .ZN(new_n889));
  OAI22_X1  g464(.A1(new_n515), .A2(new_n888), .B1(new_n522), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n560), .A2(KEYINPUT78), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n563), .B1(new_n562), .B2(new_n555), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n560), .A2(new_n892), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT38), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n891), .B1(new_n561), .B2(new_n564), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n900), .A2(new_n896), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT38), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n627), .A2(G559), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n899), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n905), .B1(new_n899), .B2(new_n903), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n885), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(G860), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n908), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n912), .A2(KEYINPUT39), .A3(new_n906), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(KEYINPUT104), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT104), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n912), .A2(new_n915), .A3(KEYINPUT39), .A4(new_n906), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n911), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n891), .A2(new_n910), .ZN(new_n919));
  XNOR2_X1  g494(.A(KEYINPUT105), .B(KEYINPUT37), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n919), .B(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  OR3_X1    g497(.A1(new_n917), .A2(new_n918), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n918), .B1(new_n917), .B2(new_n922), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(G145));
  XNOR2_X1  g500(.A(G160), .B(new_n660), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(G162), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n860), .A2(new_n843), .ZN(new_n928));
  NAND2_X1  g503(.A1(G164), .A2(new_n859), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n801), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n928), .A2(new_n801), .A3(new_n929), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n482), .A2(G130), .ZN(new_n934));
  OR2_X1    g509(.A1(G106), .A2(G2105), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n935), .B(G2104), .C1(G118), .C2(new_n463), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n937), .B1(G142), .B2(new_n480), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(new_n651), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n932), .A2(new_n933), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n939), .B1(new_n932), .B2(new_n933), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n810), .B(new_n775), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n941), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n932), .A2(new_n933), .ZN(new_n946));
  INV_X1    g521(.A(new_n939), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n943), .B1(new_n948), .B2(new_n940), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n927), .B1(new_n945), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G37), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n944), .B1(new_n941), .B2(new_n942), .ZN(new_n952));
  INV_X1    g527(.A(new_n927), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n948), .A2(new_n943), .A3(new_n940), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n950), .A2(new_n951), .A3(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n956), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g532(.A(G305), .B(new_n609), .ZN(new_n958));
  XNOR2_X1  g533(.A(G288), .B(G166), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n958), .B(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n964));
  INV_X1    g539(.A(new_n962), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n960), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n631), .A2(new_n638), .ZN(new_n969));
  NAND3_X1  g544(.A1(G299), .A2(new_n617), .A3(new_n624), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n642), .A2(KEYINPUT107), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT107), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n640), .A2(new_n973), .A3(new_n634), .A4(new_n641), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n972), .A2(new_n901), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n901), .B1(new_n972), .B2(new_n974), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n971), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n975), .A2(new_n976), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT41), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n971), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n969), .A2(new_n970), .A3(KEYINPUT41), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n977), .A2(new_n978), .B1(new_n979), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n971), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n973), .B1(new_n627), .B2(new_n634), .ZN(new_n986));
  INV_X1    g561(.A(new_n974), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n898), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n972), .A2(new_n901), .A3(new_n974), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n985), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT108), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n968), .B1(new_n984), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n988), .A2(new_n989), .A3(new_n983), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(new_n990), .B2(KEYINPUT108), .ZN(new_n994));
  AOI211_X1 g569(.A(new_n978), .B(new_n985), .C1(new_n988), .C2(new_n989), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n994), .A2(new_n967), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(G868), .B1(new_n992), .B2(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n891), .A2(G868), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n997), .A2(new_n999), .ZN(G295));
  INV_X1    g575(.A(KEYINPUT110), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n997), .A2(new_n1001), .A3(new_n999), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n967), .B1(new_n994), .B2(new_n995), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n977), .A2(new_n978), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n968), .A2(new_n1004), .A3(new_n991), .A4(new_n993), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n611), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT110), .B1(new_n1006), .B2(new_n998), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1002), .A2(new_n1007), .ZN(G331));
  AND3_X1   g583(.A1(new_n981), .A2(KEYINPUT112), .A3(new_n982), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT111), .ZN(new_n1010));
  NAND2_X1  g585(.A1(G168), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT111), .B1(new_n528), .B2(new_n532), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AND2_X1   g588(.A1(G171), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(G171), .A2(new_n1013), .ZN(new_n1015));
  OAI22_X1  g590(.A1(new_n1014), .A2(new_n1015), .B1(new_n900), .B2(new_n896), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n971), .A2(new_n1017), .A3(new_n980), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1013), .ZN(new_n1019));
  NAND2_X1  g594(.A1(G301), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(G171), .A2(new_n1013), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1020), .A2(new_n895), .A3(new_n897), .A4(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1016), .A2(new_n1018), .A3(new_n1022), .ZN(new_n1023));
  OR2_X1    g598(.A1(new_n1009), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1016), .A2(new_n1022), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n971), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n960), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n983), .A2(new_n1022), .A3(new_n1016), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1026), .A2(new_n1028), .A3(new_n960), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n951), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT43), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g608(.A(KEYINPUT113), .B(KEYINPUT43), .C1(new_n1027), .C2(new_n1030), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n960), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1035));
  OR3_X1    g610(.A1(new_n1030), .A2(KEYINPUT43), .A3(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1033), .A2(KEYINPUT44), .A3(new_n1034), .A4(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT43), .B1(new_n1030), .B2(new_n1035), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1009), .A2(new_n1023), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n985), .B1(new_n1016), .B2(new_n1022), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n961), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT43), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1041), .A2(new_n1042), .A3(new_n951), .A4(new_n1029), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1038), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT44), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1037), .A2(new_n1046), .ZN(G397));
  INV_X1    g622(.A(KEYINPUT45), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(G164), .B2(G1384), .ZN(new_n1049));
  INV_X1    g624(.A(new_n477), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n471), .A2(new_n472), .ZN(new_n1051));
  OAI211_X1 g626(.A(G40), .B(new_n1050), .C1(new_n1051), .C2(new_n463), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n860), .A2(new_n862), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n859), .A2(G2067), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G1996), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n810), .B(new_n1057), .ZN(new_n1058));
  OR2_X1    g633(.A1(new_n776), .A2(new_n778), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n776), .A2(new_n778), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1056), .A2(new_n1058), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n609), .B(new_n733), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1053), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT123), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT50), .ZN(new_n1065));
  INV_X1    g640(.A(G1384), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n843), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(G2084), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G40), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n473), .A2(new_n1070), .A3(new_n477), .ZN(new_n1071));
  AOI21_X1  g646(.A(G1384), .B1(new_n838), .B2(new_n842), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1071), .B1(new_n1072), .B2(new_n1065), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1069), .A2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1048), .A2(G1384), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1076), .B1(new_n838), .B2(new_n842), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(new_n1052), .ZN(new_n1078));
  AOI21_X1  g653(.A(G1966), .B1(new_n1078), .B2(new_n1049), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1064), .B1(new_n1074), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G1966), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1072), .A2(KEYINPUT45), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1071), .B1(G164), .B2(new_n1076), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AOI22_X1  g659(.A1(new_n499), .A2(new_n496), .B1(new_n646), .B2(new_n503), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1066), .B1(new_n1085), .B2(new_n492), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1052), .B1(new_n1086), .B2(KEYINPUT50), .ZN(new_n1087));
  AOI21_X1  g662(.A(G2084), .B1(new_n1072), .B2(new_n1065), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1084), .A2(new_n1089), .A3(KEYINPUT123), .ZN(new_n1090));
  AOI21_X1  g665(.A(G286), .B1(new_n1080), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G8), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT51), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(G168), .A2(new_n1092), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1080), .A2(new_n1090), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT51), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1084), .A2(new_n1089), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1096), .B(G8), .C1(new_n1097), .C2(G286), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1093), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT124), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n843), .A2(new_n1075), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1103), .B(new_n1071), .C1(KEYINPUT45), .C2(new_n1072), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1102), .B1(new_n1104), .B2(G2078), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT53), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1102), .B(new_n1107), .C1(new_n1104), .C2(G2078), .ZN(new_n1108));
  AOI21_X1  g683(.A(G1961), .B1(new_n1087), .B2(new_n1067), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  AND4_X1   g685(.A1(G301), .A2(new_n1106), .A3(new_n1108), .A4(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1109), .B1(new_n1105), .B2(KEYINPUT53), .ZN(new_n1112));
  AOI21_X1  g687(.A(G301), .B1(new_n1112), .B2(new_n1108), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1101), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(G303), .A2(G8), .ZN(new_n1115));
  XOR2_X1   g690(.A(new_n1115), .B(KEYINPUT55), .Z(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1067), .A2(KEYINPUT117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT117), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1072), .A2(new_n1119), .A3(new_n1065), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1073), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(G2090), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n1121), .A2(new_n1122), .B1(new_n761), .B2(new_n1104), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1117), .B1(new_n1123), .B2(new_n1092), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1104), .A2(new_n761), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1087), .A2(new_n1122), .A3(new_n1067), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1127), .A2(G8), .A3(new_n1116), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1092), .B1(new_n1072), .B2(new_n1071), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n594), .A2(G1976), .A3(new_n595), .ZN(new_n1130));
  INV_X1    g705(.A(G1976), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT52), .B1(G288), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1129), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1072), .A2(new_n1071), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n1134), .A2(G8), .A3(new_n1130), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT52), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1133), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1129), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT115), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n514), .A2(new_n600), .ZN(new_n1140));
  INV_X1    g715(.A(G86), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1140), .B1(new_n522), .B2(new_n1141), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n1142), .A2(KEYINPUT114), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n599), .B1(new_n1142), .B2(KEYINPUT114), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1139), .B1(new_n1145), .B2(new_n739), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n739), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT115), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n601), .A2(new_n602), .A3(new_n739), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1146), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT49), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1138), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1146), .A2(KEYINPUT49), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1137), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1124), .A2(new_n1128), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1106), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(G171), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1112), .A2(G301), .A3(new_n1108), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1157), .A2(KEYINPUT54), .A3(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1100), .A2(new_n1114), .A3(new_n1155), .A4(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT120), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1134), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1072), .A2(KEYINPUT120), .A3(new_n1071), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1087), .A2(new_n1067), .ZN(new_n1165));
  INV_X1    g740(.A(G1348), .ZN(new_n1166));
  AOI22_X1  g741(.A1(new_n862), .A2(new_n1164), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1167), .A2(KEYINPUT60), .A3(new_n638), .ZN(new_n1168));
  XNOR2_X1  g743(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1169), .ZN(new_n1170));
  XOR2_X1   g745(.A(KEYINPUT58), .B(G1341), .Z(new_n1171));
  NAND3_X1  g746(.A1(new_n1162), .A2(new_n1163), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1078), .A2(new_n1049), .A3(new_n1057), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1170), .B1(new_n1174), .B2(new_n566), .ZN(new_n1175));
  AOI211_X1 g750(.A(new_n565), .B(new_n1169), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1168), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1163), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT120), .B1(new_n1072), .B2(new_n1071), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n862), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1067), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1166), .B1(new_n1181), .B2(new_n1073), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1180), .A2(KEYINPUT60), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(KEYINPUT60), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1184));
  NOR3_X1   g759(.A1(new_n1183), .A2(new_n1184), .A3(new_n638), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1177), .A2(new_n1185), .ZN(new_n1186));
  OR2_X1    g761(.A1(new_n1121), .A2(G1956), .ZN(new_n1187));
  XNOR2_X1  g762(.A(KEYINPUT56), .B(G2072), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1078), .A2(new_n1049), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g765(.A(G299), .B(KEYINPUT57), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1191), .ZN(new_n1193));
  OAI211_X1 g768(.A(new_n1193), .B(new_n1189), .C1(G1956), .C2(new_n1121), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1192), .A2(KEYINPUT61), .A3(new_n1194), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1187), .A2(KEYINPUT119), .A3(new_n1193), .A4(new_n1189), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT119), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1194), .A2(new_n1197), .ZN(new_n1198));
  AOI22_X1  g773(.A1(new_n1196), .A2(new_n1198), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1199));
  OAI211_X1 g774(.A(new_n1186), .B(new_n1195), .C1(KEYINPUT61), .C2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1201));
  OAI21_X1  g776(.A(KEYINPUT121), .B1(new_n1167), .B2(new_n638), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1192), .A2(new_n1202), .ZN(new_n1203));
  NOR3_X1   g778(.A1(new_n1167), .A2(KEYINPUT121), .A3(new_n638), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1201), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1160), .B1(new_n1200), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(new_n1149), .ZN(new_n1207));
  INV_X1    g782(.A(new_n1148), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1149), .B1(new_n1147), .B2(KEYINPUT115), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1151), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1210), .A2(new_n1153), .A3(new_n1129), .ZN(new_n1211));
  NOR2_X1   g786(.A1(G288), .A2(G1976), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1207), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  XOR2_X1   g788(.A(new_n1129), .B(KEYINPUT116), .Z(new_n1214));
  AOI21_X1  g789(.A(new_n1136), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1215), .B1(new_n1135), .B2(new_n1132), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1211), .A2(new_n1216), .ZN(new_n1217));
  OAI22_X1  g792(.A1(new_n1213), .A2(new_n1214), .B1(new_n1217), .B2(new_n1128), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1116), .B1(new_n1127), .B2(G8), .ZN(new_n1219));
  INV_X1    g794(.A(new_n1219), .ZN(new_n1220));
  NAND3_X1  g795(.A1(new_n1220), .A2(new_n1154), .A3(KEYINPUT118), .ZN(new_n1221));
  INV_X1    g796(.A(KEYINPUT118), .ZN(new_n1222));
  OAI21_X1  g797(.A(new_n1222), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1223));
  AOI211_X1 g798(.A(new_n1092), .B(G286), .C1(new_n1084), .C2(new_n1089), .ZN(new_n1224));
  AND3_X1   g799(.A1(new_n1128), .A2(new_n1224), .A3(KEYINPUT63), .ZN(new_n1225));
  NAND3_X1  g800(.A1(new_n1221), .A2(new_n1223), .A3(new_n1225), .ZN(new_n1226));
  NAND4_X1  g801(.A1(new_n1124), .A2(new_n1154), .A3(new_n1128), .A4(new_n1224), .ZN(new_n1227));
  INV_X1    g802(.A(KEYINPUT63), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g804(.A(new_n1218), .B1(new_n1226), .B2(new_n1229), .ZN(new_n1230));
  AND3_X1   g805(.A1(new_n1084), .A2(new_n1089), .A3(KEYINPUT123), .ZN(new_n1231));
  AOI21_X1  g806(.A(KEYINPUT123), .B1(new_n1084), .B2(new_n1089), .ZN(new_n1232));
  OAI21_X1  g807(.A(G168), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g808(.A(new_n1096), .B1(new_n1233), .B2(G8), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1235));
  OAI21_X1  g810(.A(KEYINPUT62), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g811(.A(KEYINPUT62), .ZN(new_n1237));
  NAND3_X1  g812(.A1(new_n1093), .A2(new_n1099), .A3(new_n1237), .ZN(new_n1238));
  AND4_X1   g813(.A1(new_n1124), .A2(new_n1113), .A3(new_n1128), .A4(new_n1154), .ZN(new_n1239));
  NAND3_X1  g814(.A1(new_n1236), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g815(.A1(new_n1230), .A2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g816(.A(new_n1063), .B1(new_n1206), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g817(.A(new_n1056), .ZN(new_n1243));
  OAI21_X1  g818(.A(new_n1053), .B1(new_n1243), .B2(new_n810), .ZN(new_n1244));
  INV_X1    g819(.A(KEYINPUT46), .ZN(new_n1245));
  INV_X1    g820(.A(new_n1053), .ZN(new_n1246));
  OAI21_X1  g821(.A(new_n1245), .B1(new_n1246), .B2(G1996), .ZN(new_n1247));
  NAND3_X1  g822(.A1(new_n1053), .A2(KEYINPUT46), .A3(new_n1057), .ZN(new_n1248));
  NAND3_X1  g823(.A1(new_n1244), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  XNOR2_X1  g824(.A(new_n1249), .B(KEYINPUT47), .ZN(new_n1250));
  NAND2_X1  g825(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1251));
  OAI21_X1  g826(.A(new_n1054), .B1(new_n1251), .B2(new_n1060), .ZN(new_n1252));
  NAND2_X1  g827(.A1(new_n1252), .A2(new_n1053), .ZN(new_n1253));
  XNOR2_X1  g828(.A(new_n1253), .B(KEYINPUT125), .ZN(new_n1254));
  NAND2_X1  g829(.A1(new_n1061), .A2(new_n1053), .ZN(new_n1255));
  NOR2_X1   g830(.A1(G290), .A2(G1986), .ZN(new_n1256));
  NAND3_X1  g831(.A1(new_n1053), .A2(KEYINPUT48), .A3(new_n1256), .ZN(new_n1257));
  INV_X1    g832(.A(KEYINPUT48), .ZN(new_n1258));
  INV_X1    g833(.A(new_n1256), .ZN(new_n1259));
  OAI21_X1  g834(.A(new_n1258), .B1(new_n1246), .B2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g835(.A1(new_n1255), .A2(new_n1257), .A3(new_n1260), .ZN(new_n1261));
  AND3_X1   g836(.A1(new_n1250), .A2(new_n1254), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g837(.A1(new_n1242), .A2(new_n1262), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g838(.A1(G227), .A2(new_n461), .ZN(new_n1265));
  OAI21_X1  g839(.A(new_n1265), .B1(new_n698), .B2(new_n700), .ZN(new_n1266));
  INV_X1    g840(.A(KEYINPUT126), .ZN(new_n1267));
  NAND2_X1  g841(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g842(.A(new_n1265), .ZN(new_n1269));
  NAND2_X1  g843(.A1(new_n696), .A2(new_n697), .ZN(new_n1270));
  AOI21_X1  g844(.A(new_n1269), .B1(new_n1270), .B2(new_n699), .ZN(new_n1271));
  AOI21_X1  g845(.A(G229), .B1(new_n1271), .B2(KEYINPUT126), .ZN(new_n1272));
  AND3_X1   g846(.A1(new_n956), .A2(new_n1268), .A3(new_n1272), .ZN(new_n1273));
  AND3_X1   g847(.A1(new_n1044), .A2(new_n1273), .A3(KEYINPUT127), .ZN(new_n1274));
  AOI21_X1  g848(.A(KEYINPUT127), .B1(new_n1044), .B2(new_n1273), .ZN(new_n1275));
  NOR2_X1   g849(.A1(new_n1274), .A2(new_n1275), .ZN(G308));
  NAND2_X1  g850(.A1(new_n1044), .A2(new_n1273), .ZN(new_n1277));
  INV_X1    g851(.A(KEYINPUT127), .ZN(new_n1278));
  NAND2_X1  g852(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g853(.A1(new_n1044), .A2(new_n1273), .A3(KEYINPUT127), .ZN(new_n1280));
  NAND2_X1  g854(.A1(new_n1279), .A2(new_n1280), .ZN(G225));
endmodule


