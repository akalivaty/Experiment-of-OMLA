//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n555, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n578, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1231, new_n1232;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT66), .Z(new_n452));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n452), .A2(new_n457), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT67), .Z(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI211_X1 g038(.A(G137), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n464), .A2(KEYINPUT68), .A3(new_n465), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n462), .A2(new_n463), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(G2105), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(new_n472), .A2(new_n461), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  MUX2_X1   g055(.A(G100), .B(G112), .S(G2105), .Z(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n472), .A2(G2105), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(G136), .B2(new_n484), .ZN(G162));
  XNOR2_X1  g060(.A(KEYINPUT3), .B(G2104), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n486), .A2(G126), .A3(G2105), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n488));
  INV_X1    g063(.A(G2104), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n461), .A2(G102), .ZN(new_n490));
  NAND2_X1  g065(.A1(G114), .A2(G2105), .ZN(new_n491));
  AOI211_X1 g066(.A(new_n488), .B(new_n489), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G102), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n491), .B1(new_n493), .B2(G2105), .ZN(new_n494));
  AOI21_X1  g069(.A(KEYINPUT69), .B1(new_n494), .B2(G2104), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n487), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n486), .A2(KEYINPUT4), .A3(G138), .A4(new_n461), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n496), .A2(new_n501), .ZN(G164));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT70), .B1(new_n503), .B2(KEYINPUT6), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n505), .A2(new_n506), .A3(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n509));
  OR2_X1    g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n508), .A2(new_n509), .A3(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G88), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n510), .A2(new_n511), .ZN(new_n517));
  INV_X1    g092(.A(G62), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n508), .A2(G543), .A3(new_n509), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(new_n524), .A3(G50), .ZN(new_n525));
  INV_X1    g100(.A(G50), .ZN(new_n526));
  OAI21_X1  g101(.A(KEYINPUT71), .B1(new_n522), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n521), .B1(new_n525), .B2(new_n527), .ZN(G166));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT73), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n514), .A2(G89), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n523), .A2(G51), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n512), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n510), .A2(KEYINPUT72), .A3(new_n511), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n535), .A2(G63), .A3(G651), .A4(new_n536), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n531), .A2(new_n532), .A3(new_n533), .A4(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  NAND3_X1  g114(.A1(new_n535), .A2(G64), .A3(new_n536), .ZN(new_n540));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n503), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G52), .ZN(new_n543));
  XOR2_X1   g118(.A(KEYINPUT74), .B(G90), .Z(new_n544));
  OAI22_X1  g119(.A1(new_n543), .A2(new_n522), .B1(new_n513), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(G171));
  NAND3_X1  g121(.A1(new_n535), .A2(G56), .A3(new_n536), .ZN(new_n547));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n503), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  INV_X1    g125(.A(G81), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n550), .A2(new_n522), .B1(new_n513), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(G188));
  NAND4_X1  g134(.A1(new_n508), .A2(G53), .A3(G543), .A4(new_n509), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(KEYINPUT9), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n504), .A2(new_n507), .B1(KEYINPUT6), .B2(new_n503), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n562), .A2(new_n563), .A3(G53), .A4(G543), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n566), .B1(new_n510), .B2(new_n511), .ZN(new_n567));
  AND2_X1   g142(.A1(G78), .A2(G543), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n508), .A2(G91), .A3(new_n509), .A4(new_n512), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n565), .A2(new_n571), .ZN(G299));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n573));
  NAND2_X1  g148(.A1(G171), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT75), .B1(new_n542), .B2(new_n545), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G301));
  NAND2_X1  g152(.A1(new_n525), .A2(new_n527), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n578), .A2(new_n515), .A3(new_n520), .ZN(G303));
  NAND3_X1  g154(.A1(new_n562), .A2(G49), .A3(G543), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n562), .A2(G87), .A3(new_n512), .ZN(new_n581));
  AOI21_X1  g156(.A(G74), .B1(new_n535), .B2(new_n536), .ZN(new_n582));
  OAI211_X1 g157(.A(new_n580), .B(new_n581), .C1(new_n582), .C2(new_n503), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n583), .B(new_n584), .ZN(G288));
  NAND4_X1  g160(.A1(new_n508), .A2(G86), .A3(new_n509), .A4(new_n512), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n586), .A2(KEYINPUT77), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(KEYINPUT77), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n512), .A2(G61), .ZN(new_n589));
  AND2_X1   g164(.A1(G73), .A2(G543), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n562), .A2(G48), .A3(G543), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n587), .A2(new_n588), .A3(new_n591), .A4(new_n592), .ZN(G305));
  NAND3_X1  g168(.A1(new_n535), .A2(G60), .A3(new_n536), .ZN(new_n594));
  NAND2_X1  g169(.A1(G72), .A2(G543), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n503), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(G47), .ZN(new_n597));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  OAI22_X1  g173(.A1(new_n597), .A2(new_n522), .B1(new_n513), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G290));
  INV_X1    g176(.A(KEYINPUT78), .ZN(new_n602));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n576), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g179(.A1(G301), .A2(KEYINPUT78), .A3(G868), .ZN(new_n605));
  AND3_X1   g180(.A1(new_n562), .A2(G92), .A3(new_n512), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT10), .ZN(new_n607));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G66), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n517), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n523), .A2(G54), .B1(new_n610), .B2(G651), .ZN(new_n611));
  AND2_X1   g186(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT79), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n604), .B(new_n605), .C1(new_n613), .C2(G868), .ZN(G284));
  OAI211_X1 g189(.A(new_n604), .B(new_n605), .C1(new_n613), .C2(G868), .ZN(G321));
  MUX2_X1   g190(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g191(.A(G299), .B(G286), .S(G868), .Z(G280));
  XOR2_X1   g192(.A(KEYINPUT80), .B(G559), .Z(new_n618));
  OAI21_X1  g193(.A(new_n613), .B1(G860), .B2(new_n618), .ZN(G148));
  INV_X1    g194(.A(new_n553), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n613), .A2(new_n618), .ZN(new_n621));
  MUX2_X1   g196(.A(new_n620), .B(new_n621), .S(G868), .Z(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n486), .A2(new_n461), .ZN(new_n624));
  OR3_X1    g199(.A1(new_n624), .A2(KEYINPUT12), .A3(new_n489), .ZN(new_n625));
  OAI21_X1  g200(.A(KEYINPUT12), .B1(new_n624), .B2(new_n489), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  INV_X1    g203(.A(G2100), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n479), .A2(G123), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT81), .ZN(new_n632));
  MUX2_X1   g207(.A(G99), .B(G111), .S(G2105), .Z(new_n633));
  AOI22_X1  g208(.A1(new_n484), .A2(G135), .B1(G2104), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT82), .B(G2096), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n628), .A2(new_n629), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n630), .A2(new_n637), .A3(new_n638), .ZN(G156));
  XOR2_X1   g214(.A(G2451), .B(G2454), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT83), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT84), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2430), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  AND3_X1   g228(.A1(new_n652), .A2(KEYINPUT14), .A3(new_n653), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n646), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n646), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(G14), .A3(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G401));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  XNOR2_X1  g234(.A(G2072), .B(G2078), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT18), .Z(new_n663));
  INV_X1    g238(.A(new_n659), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n660), .A2(KEYINPUT17), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(new_n661), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(new_n664), .B2(new_n665), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n659), .A2(new_n661), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n660), .B1(new_n669), .B2(KEYINPUT17), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n663), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(G2096), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n671), .A2(G2096), .ZN(new_n674));
  OR3_X1    g249(.A1(new_n673), .A2(new_n629), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n629), .B1(new_n673), .B2(new_n674), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(G227));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1956), .B(G2474), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n681), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n681), .A2(new_n684), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT20), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR3_X1   g264(.A1(new_n681), .A2(KEYINPUT20), .A3(new_n684), .ZN(new_n690));
  OAI221_X1 g265(.A(new_n686), .B1(new_n681), .B2(new_n685), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT86), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n691), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G1991), .B(G1996), .Z(new_n695));
  XOR2_X1   g270(.A(G1981), .B(G1986), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n694), .A2(new_n697), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(G229));
  NOR2_X1   g276(.A1(G16), .A2(G22), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(G166), .B2(G16), .ZN(new_n703));
  INV_X1    g278(.A(G1971), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  OR2_X1    g280(.A1(G6), .A2(G16), .ZN(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(G305), .B2(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT88), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT32), .B(G1981), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT88), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n708), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(new_n710), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n707), .A2(G23), .ZN(new_n716));
  INV_X1    g291(.A(new_n583), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n716), .B1(new_n717), .B2(new_n707), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT33), .B(G1976), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n705), .A2(new_n712), .A3(new_n715), .A4(new_n720), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n721), .A2(KEYINPUT34), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(KEYINPUT34), .ZN(new_n723));
  NOR2_X1   g298(.A1(G25), .A2(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n484), .A2(G131), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n479), .A2(G119), .ZN(new_n726));
  MUX2_X1   g301(.A(G95), .B(G107), .S(G2105), .Z(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G2104), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n725), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n724), .B1(new_n730), .B2(G29), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT35), .B(G1991), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(G16), .A2(G24), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n600), .B2(G16), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT87), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1986), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n722), .A2(new_n723), .A3(new_n733), .A4(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT36), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n484), .A2(G141), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT96), .ZN(new_n741));
  NAND3_X1  g316(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT26), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT97), .ZN(new_n745));
  AOI211_X1 g320(.A(new_n743), .B(new_n745), .C1(G129), .C2(new_n479), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n741), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G29), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n748), .B2(G32), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT27), .B(G1996), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT98), .ZN(new_n753));
  NOR2_X1   g328(.A1(G29), .A2(G35), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G162), .B2(G29), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT29), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n756), .A2(G2090), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n757), .A2(KEYINPUT101), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(KEYINPUT101), .ZN(new_n759));
  NOR2_X1   g334(.A1(G5), .A2(G16), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT100), .Z(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G171), .B2(G16), .ZN(new_n762));
  INV_X1    g337(.A(G1961), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  AND4_X1   g339(.A1(new_n753), .A2(new_n758), .A3(new_n759), .A4(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(G168), .A2(new_n707), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n707), .B2(G21), .ZN(new_n767));
  INV_X1    g342(.A(G1966), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n769), .B(new_n770), .C1(G2090), .C2(new_n756), .ZN(new_n771));
  NOR2_X1   g346(.A1(G16), .A2(G19), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n553), .B2(G16), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1341), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT31), .B(G11), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT99), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n635), .A2(new_n748), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT30), .B(G28), .ZN(new_n778));
  AOI211_X1 g353(.A(new_n776), .B(new_n777), .C1(new_n748), .C2(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G27), .A2(G29), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G164), .B2(G29), .ZN(new_n781));
  INV_X1    g356(.A(G2078), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n779), .B(new_n783), .C1(new_n750), .C2(new_n751), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n771), .A2(new_n774), .A3(new_n784), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n748), .A2(G26), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  OAI211_X1 g363(.A(G128), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT90), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n486), .A2(KEYINPUT90), .A3(G128), .A4(G2105), .ZN(new_n792));
  MUX2_X1   g367(.A(G104), .B(G116), .S(G2105), .Z(new_n793));
  AOI22_X1  g368(.A1(new_n791), .A2(new_n792), .B1(G2104), .B2(new_n793), .ZN(new_n794));
  OAI211_X1 g369(.A(G140), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT89), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n486), .A2(KEYINPUT89), .A3(G140), .A4(new_n461), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n794), .A2(KEYINPUT91), .A3(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(KEYINPUT91), .B1(new_n794), .B2(new_n799), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n788), .B1(new_n804), .B2(G29), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G2067), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n748), .A2(G33), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n486), .A2(G127), .ZN(new_n808));
  NAND2_X1  g383(.A1(G115), .A2(G2104), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n461), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(KEYINPUT93), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(KEYINPUT93), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT25), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n814), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n484), .A2(G139), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n811), .A2(new_n812), .A3(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT94), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n807), .B1(new_n820), .B2(new_n748), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(G2072), .Z(new_n822));
  NAND4_X1  g397(.A1(new_n765), .A2(new_n785), .A3(new_n806), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n707), .A2(G4), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n613), .B2(new_n707), .ZN(new_n825));
  INV_X1    g400(.A(G1348), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n707), .A2(G20), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT102), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT23), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(G299), .B2(G16), .ZN(new_n831));
  INV_X1    g406(.A(G1956), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  AND2_X1   g408(.A1(KEYINPUT24), .A2(G34), .ZN(new_n834));
  NOR2_X1   g409(.A1(KEYINPUT24), .A2(G34), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n748), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n477), .B2(new_n748), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT95), .ZN(new_n838));
  INV_X1    g413(.A(G2084), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n833), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n827), .B(new_n840), .C1(new_n839), .C2(new_n838), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n823), .A2(new_n841), .ZN(new_n842));
  AND2_X1   g417(.A1(new_n739), .A2(new_n842), .ZN(G311));
  NAND2_X1  g418(.A1(new_n739), .A2(new_n842), .ZN(G150));
  INV_X1    g419(.A(KEYINPUT106), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT39), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n613), .A2(G559), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n607), .A2(new_n611), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT79), .ZN(new_n851));
  INV_X1    g426(.A(G559), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n847), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT104), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n553), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n535), .A2(G67), .A3(new_n536), .ZN(new_n856));
  NAND2_X1  g431(.A1(G80), .A2(G543), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n503), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(G55), .ZN(new_n859));
  INV_X1    g434(.A(G93), .ZN(new_n860));
  OAI22_X1  g435(.A1(new_n859), .A2(new_n522), .B1(new_n513), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(KEYINPUT104), .B1(new_n549), .B2(new_n552), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n855), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n553), .A2(new_n862), .A3(new_n854), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n849), .A2(new_n853), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n867), .B1(new_n849), .B2(new_n853), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n846), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(G860), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n868), .A2(new_n869), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT105), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n873), .A2(new_n874), .A3(KEYINPUT39), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n849), .A2(new_n853), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n865), .A2(new_n866), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n849), .A2(new_n853), .A3(new_n867), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(KEYINPUT39), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(KEYINPUT105), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n872), .B1(new_n875), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n863), .A2(G860), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(KEYINPUT37), .Z(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n845), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n870), .A2(new_n871), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n874), .B1(new_n873), .B2(KEYINPUT39), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n880), .A2(KEYINPUT105), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n890), .A2(KEYINPUT106), .A3(new_n884), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n886), .A2(new_n891), .ZN(G145));
  INV_X1    g467(.A(KEYINPUT110), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT109), .ZN(new_n894));
  INV_X1    g469(.A(new_n820), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n494), .A2(G2104), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(new_n488), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n494), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n899), .A2(new_n487), .A3(new_n499), .A4(new_n500), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n801), .A2(new_n900), .A3(new_n802), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n791), .A2(new_n792), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n793), .A2(G2104), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n799), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT91), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(G164), .B1(new_n906), .B2(new_n800), .ZN(new_n907));
  NOR3_X1   g482(.A1(new_n901), .A2(new_n907), .A3(new_n747), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n741), .A2(new_n746), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n900), .B1(new_n801), .B2(new_n802), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n906), .A2(G164), .A3(new_n800), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n895), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n747), .B1(new_n901), .B2(new_n907), .ZN(new_n914));
  INV_X1    g489(.A(new_n818), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n910), .A2(new_n909), .A3(new_n911), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n627), .B(new_n729), .ZN(new_n919));
  MUX2_X1   g494(.A(G106), .B(G118), .S(G2105), .Z(new_n920));
  AOI22_X1  g495(.A1(new_n484), .A2(G142), .B1(G2104), .B2(new_n920), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n479), .A2(KEYINPUT108), .A3(G130), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT108), .B1(new_n479), .B2(G130), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n919), .B(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n894), .B1(new_n918), .B2(new_n926), .ZN(new_n927));
  AOI211_X1 g502(.A(KEYINPUT109), .B(new_n925), .C1(new_n913), .C2(new_n917), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n893), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n908), .A2(new_n912), .A3(new_n818), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n820), .B1(new_n914), .B2(new_n916), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n926), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT109), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n918), .A2(new_n894), .A3(new_n926), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(KEYINPUT110), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n913), .A2(new_n925), .A3(new_n917), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n929), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n635), .B(KEYINPUT107), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n477), .B(G162), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n938), .B(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n933), .A2(new_n934), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n936), .A2(new_n940), .ZN(new_n944));
  AOI21_X1  g519(.A(G37), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n942), .A2(KEYINPUT40), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT40), .B1(new_n942), .B2(new_n945), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(G395));
  NOR2_X1   g523(.A1(new_n863), .A2(G868), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n850), .A2(G299), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n607), .A2(new_n565), .A3(new_n571), .A4(new_n611), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n950), .A2(KEYINPUT41), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(KEYINPUT41), .B1(new_n950), .B2(new_n951), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT111), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n621), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n613), .A2(KEYINPUT111), .A3(new_n618), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n956), .A2(new_n877), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n877), .B1(new_n956), .B2(new_n957), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n954), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n956), .A2(new_n957), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n867), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n956), .A2(new_n877), .A3(new_n957), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n950), .A2(new_n951), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n960), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n717), .B(new_n600), .ZN(new_n968));
  NAND2_X1  g543(.A1(G303), .A2(G305), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(G303), .A2(G305), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n968), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n971), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n600), .B(new_n583), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n973), .A2(new_n974), .A3(new_n969), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT112), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT112), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n972), .A2(new_n975), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT42), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n976), .A2(KEYINPUT42), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n967), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n960), .A2(new_n966), .A3(new_n983), .A4(new_n981), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n949), .B1(new_n987), .B2(G868), .ZN(G295));
  AOI21_X1  g563(.A(new_n949), .B1(new_n987), .B2(G868), .ZN(G331));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n574), .A2(G168), .A3(new_n575), .ZN(new_n991));
  NAND2_X1  g566(.A1(G286), .A2(G171), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n877), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n991), .A2(new_n992), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n867), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n954), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n999), .B1(new_n867), .B2(new_n995), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n993), .A2(KEYINPUT113), .A3(new_n877), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n1000), .A2(new_n1001), .A3(new_n965), .A4(new_n996), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT114), .ZN(new_n1004));
  INV_X1    g579(.A(new_n979), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n978), .B1(new_n972), .B2(new_n975), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1004), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n977), .A2(KEYINPUT114), .A3(new_n979), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1003), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G37), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1000), .A2(new_n1001), .A3(new_n996), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n954), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n995), .B(new_n877), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n965), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1012), .A2(new_n980), .A3(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1009), .A2(new_n1010), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT43), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1018), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1019));
  AOI22_X1  g594(.A1(new_n1011), .A2(new_n954), .B1(new_n1013), .B2(new_n965), .ZN(new_n1020));
  AOI21_X1  g595(.A(G37), .B1(new_n1020), .B2(new_n980), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT43), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1019), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n990), .B1(new_n1017), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1016), .A2(new_n1022), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1019), .A2(new_n1021), .A3(KEYINPUT43), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT44), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1024), .A2(new_n1027), .ZN(G397));
  INV_X1    g603(.A(G1384), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1029), .B1(new_n496), .B2(new_n501), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT45), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n476), .A2(new_n468), .A3(G40), .A4(new_n469), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n803), .B(G2067), .ZN(new_n1035));
  INV_X1    g610(.A(G1996), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n909), .B(new_n1036), .ZN(new_n1037));
  OR2_X1    g612(.A1(new_n730), .A2(new_n732), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n730), .A2(new_n732), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1035), .A2(new_n1037), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G1986), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n600), .B(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1034), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G2090), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1033), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT50), .B1(new_n900), .B2(new_n1029), .ZN(new_n1046));
  OAI211_X1 g621(.A(KEYINPUT50), .B(new_n1029), .C1(new_n496), .C2(new_n501), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1044), .B(new_n1045), .C1(new_n1046), .C2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT115), .ZN(new_n1050));
  OAI211_X1 g625(.A(KEYINPUT45), .B(new_n1029), .C1(new_n496), .C2(new_n501), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1032), .A2(new_n1045), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n704), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT50), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1030), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1033), .B1(new_n1055), .B2(new_n1047), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(new_n1057), .A3(new_n1044), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1050), .A2(new_n1053), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n1060));
  INV_X1    g635(.A(G8), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1060), .B1(G166), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1059), .A2(G8), .A3(new_n1064), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1044), .A2(new_n1056), .B1(new_n1052), .B2(new_n704), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1066), .B1(new_n1061), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(G8), .B1(new_n1030), .B2(new_n1033), .ZN(new_n1069));
  INV_X1    g644(.A(G1976), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n583), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT52), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1073), .A2(KEYINPUT116), .ZN(new_n1074));
  NOR2_X1   g649(.A1(KEYINPUT52), .A2(G1976), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1072), .A2(new_n1074), .B1(G288), .B2(new_n1075), .ZN(new_n1076));
  OAI22_X1  g651(.A1(new_n1069), .A2(new_n1071), .B1(KEYINPUT116), .B2(new_n1073), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n591), .A2(new_n586), .A3(new_n592), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(G1981), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1079), .B1(G305), .B2(G1981), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT49), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1069), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  OR2_X1    g657(.A1(G305), .A2(G1981), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1083), .A2(KEYINPUT49), .A3(new_n1079), .ZN(new_n1084));
  AOI22_X1  g659(.A1(new_n1076), .A2(new_n1077), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1065), .A2(new_n1068), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT51), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1052), .A2(new_n768), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n839), .B(new_n1045), .C1(new_n1046), .C2(new_n1048), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1061), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(G168), .A2(new_n1061), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1087), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1091), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n839), .A2(new_n1056), .B1(new_n1052), .B2(new_n768), .ZN(new_n1094));
  OAI211_X1 g669(.A(KEYINPUT51), .B(new_n1093), .C1(new_n1094), .C2(new_n1061), .ZN(new_n1095));
  NOR4_X1   g670(.A1(new_n1094), .A2(KEYINPUT120), .A3(new_n1061), .A4(G168), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1097), .B1(new_n1090), .B2(G286), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1092), .B(new_n1095), .C1(new_n1096), .C2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1045), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n763), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1032), .A2(new_n782), .A3(new_n1045), .A4(new_n1051), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1101), .B(new_n1102), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  OAI22_X1  g680(.A1(G1961), .A2(new_n1056), .B1(new_n1104), .B2(new_n1103), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT121), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1104), .A2(new_n1103), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1105), .A2(new_n1107), .A3(G301), .A4(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT45), .B1(new_n900), .B2(new_n1029), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1051), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n476), .A2(KEYINPUT53), .A3(G40), .A4(new_n782), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1114), .B1(KEYINPUT122), .B2(new_n470), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1113), .B(new_n1115), .C1(KEYINPUT122), .C2(new_n470), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1116), .A2(new_n1101), .A3(new_n1108), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1110), .B1(new_n1117), .B2(G171), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1109), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1086), .A2(new_n1099), .A3(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1105), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n576), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1117), .A2(new_n576), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT54), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1120), .A2(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT56), .B(G2072), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1032), .A2(new_n1045), .A3(new_n1051), .A4(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n1056), .B2(G1956), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT57), .ZN(new_n1129));
  NAND2_X1  g704(.A1(G299), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n565), .A2(KEYINPUT57), .A3(new_n571), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1128), .A2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1056), .A2(G1348), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1030), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n1045), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1137), .A2(G2067), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1134), .B1(new_n1139), .B2(new_n850), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1132), .B(new_n1127), .C1(new_n1056), .C2(G1956), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT61), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1100), .A2(new_n832), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1132), .B1(new_n1144), .B2(new_n1127), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1141), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1143), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT60), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1148), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1149));
  OAI221_X1 g724(.A(KEYINPUT60), .B1(new_n1137), .B2(G2067), .C1(new_n1056), .C2(G1348), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1149), .A2(new_n612), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1139), .A2(KEYINPUT60), .A3(new_n850), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1134), .A2(KEYINPUT61), .A3(new_n1141), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1147), .A2(new_n1151), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT59), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1155), .A2(KEYINPUT118), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g732(.A(KEYINPUT58), .B(G1341), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1158), .B1(new_n1136), .B2(new_n1045), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1113), .A2(KEYINPUT117), .A3(new_n1036), .A4(new_n1045), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1032), .A2(new_n1036), .A3(new_n1045), .A4(new_n1051), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT117), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1159), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1157), .B1(new_n1164), .B2(new_n620), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1161), .B(KEYINPUT117), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n553), .B(new_n1156), .C1(new_n1166), .C2(new_n1159), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g743(.A(KEYINPUT119), .B(new_n1142), .C1(new_n1154), .C2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1142), .B1(new_n1154), .B2(new_n1168), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT119), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  AND3_X1   g747(.A1(new_n1125), .A2(new_n1169), .A3(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1065), .A2(new_n1068), .A3(new_n1085), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1122), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT62), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1099), .A2(new_n1176), .ZN(new_n1177));
  AND2_X1   g752(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1090), .A2(G286), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(KEYINPUT120), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1090), .A2(new_n1097), .A3(G286), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(KEYINPUT62), .B1(new_n1178), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1175), .B1(new_n1177), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT63), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1090), .A2(G168), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1059), .A2(G8), .ZN(new_n1187));
  AOI211_X1 g762(.A(new_n1185), .B(new_n1186), .C1(new_n1187), .C2(new_n1066), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1188), .A2(new_n1065), .A3(new_n1085), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1185), .B1(new_n1174), .B2(new_n1186), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1192));
  INV_X1    g767(.A(G288), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1192), .A2(new_n1070), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1069), .B1(new_n1194), .B2(new_n1083), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1065), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1195), .B1(new_n1196), .B2(new_n1085), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1184), .A2(new_n1191), .A3(new_n1197), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1043), .B1(new_n1173), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1040), .A2(new_n1034), .ZN(new_n1200));
  OR2_X1    g775(.A1(new_n1200), .A2(KEYINPUT124), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1200), .A2(KEYINPUT124), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1034), .A2(new_n1041), .A3(new_n600), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1203), .B(KEYINPUT125), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1204), .B(KEYINPUT48), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1201), .A2(new_n1202), .A3(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(G2067), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n803), .B(new_n1207), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1034), .B1(new_n1208), .B2(new_n909), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n1210), .B(KEYINPUT46), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1212));
  XOR2_X1   g787(.A(KEYINPUT123), .B(KEYINPUT47), .Z(new_n1213));
  XNOR2_X1  g788(.A(new_n1212), .B(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1215));
  OAI22_X1  g790(.A1(new_n1215), .A2(new_n1039), .B1(G2067), .B2(new_n804), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1216), .A2(new_n1034), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n1206), .A2(new_n1214), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g793(.A(KEYINPUT126), .ZN(new_n1219));
  XNOR2_X1  g794(.A(new_n1218), .B(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1199), .A2(new_n1220), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g796(.A1(new_n677), .A2(G319), .ZN(new_n1223));
  NAND4_X1  g797(.A1(new_n1223), .A2(new_n657), .A3(KEYINPUT127), .A4(new_n700), .ZN(new_n1224));
  NAND3_X1  g798(.A1(new_n657), .A2(new_n700), .A3(new_n1223), .ZN(new_n1225));
  INV_X1    g799(.A(KEYINPUT127), .ZN(new_n1226));
  NAND2_X1  g800(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND4_X1  g801(.A1(new_n1025), .A2(new_n1026), .A3(new_n1224), .A4(new_n1227), .ZN(new_n1228));
  AND2_X1   g802(.A1(new_n942), .A2(new_n945), .ZN(new_n1229));
  NOR2_X1   g803(.A1(new_n1228), .A2(new_n1229), .ZN(G308));
  AND2_X1   g804(.A1(new_n1227), .A2(new_n1224), .ZN(new_n1231));
  NAND2_X1  g805(.A1(new_n942), .A2(new_n945), .ZN(new_n1232));
  NAND4_X1  g806(.A1(new_n1231), .A2(new_n1232), .A3(new_n1025), .A4(new_n1026), .ZN(G225));
endmodule


