//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 1 1 0 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962;
  INV_X1    g000(.A(KEYINPUT28), .ZN(new_n187));
  XNOR2_X1  g001(.A(G143), .B(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT0), .A2(G128), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  OR2_X1    g004(.A1(KEYINPUT0), .A2(G128), .ZN(new_n191));
  AND2_X1   g005(.A1(new_n191), .A2(new_n189), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n190), .B1(new_n192), .B2(new_n188), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  OAI22_X1  g009(.A1(new_n194), .A2(KEYINPUT11), .B1(new_n195), .B2(G137), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT11), .ZN(new_n197));
  INV_X1    g011(.A(G137), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n197), .A2(new_n198), .A3(KEYINPUT64), .A4(G134), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n196), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  AOI22_X1  g015(.A1(new_n194), .A2(KEYINPUT11), .B1(new_n195), .B2(G137), .ZN(new_n202));
  AND3_X1   g016(.A1(new_n200), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n201), .B1(new_n200), .B2(new_n202), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n193), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  AND4_X1   g019(.A1(KEYINPUT64), .A2(new_n197), .A3(new_n198), .A4(G134), .ZN(new_n206));
  AOI22_X1  g020(.A1(KEYINPUT64), .A2(new_n197), .B1(new_n198), .B2(G134), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n201), .B(new_n202), .C1(new_n206), .C2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT1), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n210), .A2(new_n212), .A3(new_n213), .A4(G128), .ZN(new_n214));
  INV_X1    g028(.A(G128), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(new_n211), .A3(G143), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n209), .B(G146), .C1(new_n215), .C2(KEYINPUT1), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n214), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n198), .A2(G134), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n195), .A2(G137), .ZN(new_n220));
  OAI21_X1  g034(.A(G131), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n208), .A2(new_n218), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n205), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT2), .B(G113), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(G116), .B(G119), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n226), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(new_n224), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n187), .B1(new_n223), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n223), .A2(new_n230), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT65), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n222), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n230), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n208), .A2(new_n218), .A3(KEYINPUT65), .A4(new_n221), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n234), .A2(new_n205), .A3(new_n235), .A4(new_n236), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n231), .B(new_n232), .C1(new_n187), .C2(new_n237), .ZN(new_n238));
  XOR2_X1   g052(.A(KEYINPUT66), .B(KEYINPUT27), .Z(new_n239));
  NOR2_X1   g053(.A1(G237), .A2(G953), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G210), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n239), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT26), .B(G101), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n242), .B(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n238), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n237), .A2(new_n247), .A3(new_n244), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n247), .B1(new_n237), .B2(new_n244), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n234), .A2(new_n205), .A3(new_n236), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT30), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT30), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n205), .A2(new_n253), .A3(new_n222), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(new_n230), .ZN(new_n256));
  AOI21_X1  g070(.A(KEYINPUT31), .B1(new_n250), .B2(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n235), .B1(new_n252), .B2(new_n254), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT31), .ZN(new_n259));
  NOR4_X1   g073(.A1(new_n258), .A2(new_n248), .A3(new_n249), .A4(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n246), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G472), .ZN(new_n262));
  INV_X1    g076(.A(G902), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT32), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n237), .A2(new_n244), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT67), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n237), .A2(new_n244), .A3(new_n247), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n259), .B1(new_n270), .B2(new_n258), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n250), .A2(KEYINPUT31), .A3(new_n256), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(G902), .B1(new_n273), .B2(new_n246), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n274), .A2(KEYINPUT32), .A3(new_n262), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n251), .A2(new_n230), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n237), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT28), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n278), .A2(new_n231), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT29), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n245), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(G902), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n256), .A2(new_n237), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n245), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n280), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n238), .A2(new_n245), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n282), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G472), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n266), .A2(new_n275), .A3(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(G119), .B(G128), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n290), .B(KEYINPUT68), .ZN(new_n291));
  XOR2_X1   g105(.A(KEYINPUT24), .B(G110), .Z(new_n292));
  OAI21_X1  g106(.A(KEYINPUT23), .B1(new_n215), .B2(G119), .ZN(new_n293));
  AOI21_X1  g107(.A(KEYINPUT69), .B1(new_n215), .B2(G119), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n293), .B(new_n294), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n291), .A2(new_n292), .B1(new_n295), .B2(G110), .ZN(new_n296));
  INV_X1    g110(.A(G140), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G125), .ZN(new_n298));
  INV_X1    g112(.A(G125), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G140), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n298), .A2(new_n300), .A3(KEYINPUT70), .A4(KEYINPUT16), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n298), .A2(new_n300), .A3(KEYINPUT16), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT16), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n297), .A3(G125), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT70), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n211), .B(new_n301), .C1(new_n302), .C2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n298), .A2(new_n300), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n305), .B(new_n304), .C1(new_n309), .C2(new_n303), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n211), .B1(new_n310), .B2(new_n301), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n296), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  OAI22_X1  g126(.A1(new_n291), .A2(new_n292), .B1(new_n295), .B2(G110), .ZN(new_n313));
  INV_X1    g127(.A(new_n311), .ZN(new_n314));
  INV_X1    g128(.A(new_n309), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n211), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n313), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G953), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(G221), .A3(G234), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(KEYINPUT22), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n321), .B(G137), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n312), .A2(new_n317), .A3(new_n322), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI22_X1  g140(.A1(new_n326), .A2(G902), .B1(KEYINPUT71), .B2(KEYINPUT25), .ZN(new_n327));
  INV_X1    g141(.A(G217), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n328), .B1(G234), .B2(new_n263), .ZN(new_n329));
  NOR2_X1   g143(.A1(KEYINPUT71), .A2(KEYINPUT25), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n324), .A2(new_n263), .A3(new_n325), .A4(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n327), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n329), .A2(G902), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n324), .A2(new_n325), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n308), .A2(new_n311), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT17), .ZN(new_n338));
  INV_X1    g152(.A(G237), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(new_n319), .A3(G214), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n209), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n240), .A2(G143), .A3(G214), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n201), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n342), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT84), .B1(new_n344), .B2(G131), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT84), .ZN(new_n346));
  AOI211_X1 g160(.A(new_n346), .B(new_n201), .C1(new_n341), .C2(new_n342), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n338), .B(new_n343), .C1(new_n345), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n344), .A2(G131), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n346), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n344), .A2(KEYINPUT84), .A3(G131), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(KEYINPUT17), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n337), .A2(new_n348), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n309), .A2(G146), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n316), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT18), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n356), .A2(new_n201), .ZN(new_n357));
  OAI221_X1 g171(.A(new_n355), .B1(new_n344), .B2(new_n357), .C1(new_n349), .C2(new_n356), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G113), .ZN(new_n360));
  INV_X1    g174(.A(G122), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(G113), .A2(G122), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OR2_X1    g178(.A1(new_n364), .A2(KEYINPUT86), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(KEYINPUT86), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n365), .A2(G104), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(G104), .B1(new_n365), .B2(new_n366), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n359), .A2(new_n369), .ZN(new_n370));
  XOR2_X1   g184(.A(KEYINPUT85), .B(KEYINPUT19), .Z(new_n371));
  NAND2_X1  g185(.A1(new_n315), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT85), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n309), .B1(new_n373), .B2(KEYINPUT19), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(G146), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n376), .A2(new_n311), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n343), .B1(new_n345), .B2(new_n347), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n369), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n358), .ZN(new_n380));
  INV_X1    g194(.A(G475), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n370), .A2(new_n380), .A3(new_n381), .A4(new_n263), .ZN(new_n382));
  XNOR2_X1  g196(.A(KEYINPUT83), .B(KEYINPUT20), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI22_X1  g198(.A1(new_n359), .A2(new_n369), .B1(new_n379), .B2(new_n358), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT20), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n385), .A2(new_n386), .A3(new_n381), .A4(new_n263), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G107), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT88), .ZN(new_n390));
  INV_X1    g204(.A(G116), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n390), .B1(new_n391), .B2(G122), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n361), .A2(KEYINPUT88), .A3(G116), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n391), .A2(G122), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n389), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n394), .A2(new_n389), .A3(new_n395), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(KEYINPUT89), .A2(KEYINPUT13), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n209), .A2(G128), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n215), .A2(G143), .ZN(new_n403));
  NAND2_X1  g217(.A1(KEYINPUT89), .A2(KEYINPUT13), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n401), .A2(new_n402), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n404), .ZN(new_n406));
  OAI211_X1 g220(.A(G128), .B(new_n209), .C1(new_n406), .C2(new_n400), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n405), .A2(new_n407), .A3(G134), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT90), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n402), .A2(new_n403), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n195), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT90), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n405), .A2(new_n407), .A3(new_n412), .A4(G134), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n399), .A2(new_n409), .A3(new_n411), .A4(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n410), .B(new_n195), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n395), .B(KEYINPUT14), .ZN(new_n416));
  INV_X1    g230(.A(new_n394), .ZN(new_n417));
  OAI21_X1  g231(.A(G107), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n415), .A2(new_n418), .A3(new_n398), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT9), .B(G234), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n420), .B(KEYINPUT72), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(G217), .A3(new_n319), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n414), .A2(new_n419), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n423), .B1(new_n414), .B2(new_n419), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n263), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G478), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n428), .A2(KEYINPUT15), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n427), .B(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(KEYINPUT87), .B1(new_n367), .B2(new_n368), .ZN(new_n432));
  OR2_X1    g246(.A1(new_n359), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(G902), .B1(new_n359), .B2(new_n432), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n381), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n388), .A2(new_n431), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n421), .A2(new_n263), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G221), .ZN(new_n439));
  XOR2_X1   g253(.A(new_n439), .B(KEYINPUT73), .Z(new_n440));
  INV_X1    g254(.A(G469), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT12), .ZN(new_n442));
  INV_X1    g256(.A(G104), .ZN(new_n443));
  OAI21_X1  g257(.A(KEYINPUT3), .B1(new_n443), .B2(G107), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT3), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(new_n389), .A3(G104), .ZN(new_n446));
  INV_X1    g260(.A(G101), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n443), .A2(G107), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n444), .A2(new_n446), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n389), .A2(G104), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n443), .A2(G107), .ZN(new_n451));
  OAI21_X1  g265(.A(G101), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(new_n218), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n203), .A2(new_n204), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n442), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OR2_X1    g270(.A1(new_n203), .A2(new_n204), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n218), .A2(new_n452), .A3(new_n449), .ZN(new_n458));
  INV_X1    g272(.A(new_n453), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n459), .A2(new_n218), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n457), .B(KEYINPUT12), .C1(new_n458), .C2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  OR2_X1    g276(.A1(new_n458), .A2(KEYINPUT10), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT76), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n449), .A2(new_n452), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n464), .B1(new_n449), .B2(new_n452), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(KEYINPUT10), .A3(new_n218), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n444), .A2(new_n446), .A3(new_n448), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT4), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(new_n470), .A3(G101), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT75), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n469), .A2(KEYINPUT75), .A3(new_n470), .A4(G101), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n469), .A2(G101), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n476), .A2(KEYINPUT4), .A3(new_n449), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n475), .A2(new_n193), .A3(new_n477), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n463), .A2(new_n468), .A3(new_n478), .A4(new_n455), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n462), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(G110), .B(G140), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT74), .ZN(new_n482));
  INV_X1    g296(.A(G227), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n483), .A2(G953), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n482), .B(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n480), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n463), .A2(new_n468), .A3(new_n478), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n457), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(new_n479), .A3(new_n485), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n441), .B1(new_n491), .B2(new_n263), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT77), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n440), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n479), .A2(new_n485), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n495), .A2(new_n489), .B1(new_n480), .B2(new_n486), .ZN(new_n496));
  OAI21_X1  g310(.A(G469), .B1(new_n496), .B2(G902), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n485), .B1(new_n489), .B2(new_n479), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n462), .A2(new_n479), .A3(new_n485), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n441), .B(new_n263), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n497), .A2(KEYINPUT77), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n437), .A2(new_n494), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(G214), .B1(G237), .B2(G902), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n319), .A2(G952), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n505), .B1(G234), .B2(G237), .ZN(new_n506));
  XOR2_X1   g320(.A(KEYINPUT21), .B(G898), .Z(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  AOI211_X1 g322(.A(new_n263), .B(new_n319), .C1(G234), .C2(G237), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n218), .A2(new_n299), .ZN(new_n512));
  AOI22_X1  g326(.A1(new_n210), .A2(new_n212), .B1(new_n191), .B2(new_n189), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n210), .A2(new_n212), .A3(new_n189), .ZN(new_n514));
  OAI21_X1  g328(.A(G125), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(G224), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n517), .A2(G953), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n516), .B(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n475), .A2(new_n230), .A3(new_n477), .ZN(new_n521));
  INV_X1    g335(.A(G119), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(G116), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n523), .A2(KEYINPUT5), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(new_n360), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n391), .A2(G119), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n523), .A2(new_n526), .A3(KEYINPUT5), .ZN(new_n527));
  AOI22_X1  g341(.A1(new_n525), .A2(new_n527), .B1(new_n225), .B2(new_n226), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n467), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n521), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(G110), .B(G122), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n521), .A2(new_n529), .A3(new_n531), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(KEYINPUT6), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n531), .B1(new_n521), .B2(new_n529), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT78), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT6), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n537), .B1(new_n536), .B2(new_n538), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n520), .B(new_n535), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT79), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n527), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n226), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n525), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n227), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n459), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n528), .A2(new_n453), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n531), .B(KEYINPUT8), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT80), .ZN(new_n551));
  OR2_X1    g365(.A1(new_n518), .A2(KEYINPUT81), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n512), .A2(new_n515), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n519), .A2(KEYINPUT7), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n553), .B(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT80), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n547), .A2(new_n548), .A3(new_n556), .A4(new_n549), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n551), .A2(new_n555), .A3(new_n534), .A4(new_n557), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n558), .A2(new_n263), .ZN(new_n559));
  OAI21_X1  g373(.A(G210), .B1(G237), .B2(G902), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT82), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n541), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n562), .B1(new_n541), .B2(new_n559), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n504), .B(new_n511), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n289), .A2(new_n336), .A3(new_n503), .A4(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(G101), .ZN(G3));
  NOR2_X1   g382(.A1(new_n262), .A2(KEYINPUT91), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n274), .B(new_n569), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n494), .A2(new_n501), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n336), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT33), .B1(new_n425), .B2(new_n426), .ZN(new_n573));
  INV_X1    g387(.A(new_n426), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT33), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n575), .A3(new_n424), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n573), .A2(new_n576), .A3(G478), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n428), .B(new_n263), .C1(new_n425), .C2(new_n426), .ZN(new_n578));
  NAND2_X1  g392(.A1(G478), .A2(G902), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n580), .B1(new_n388), .B2(new_n436), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n572), .A2(new_n565), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(KEYINPUT34), .B(G104), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n583), .B(new_n584), .ZN(G6));
  NOR2_X1   g399(.A1(new_n382), .A2(new_n383), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT92), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n435), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n431), .ZN(new_n589));
  INV_X1    g403(.A(new_n383), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n385), .A2(new_n381), .A3(new_n263), .A4(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n384), .A2(KEYINPUT92), .A3(new_n591), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n588), .A2(new_n511), .A3(new_n589), .A4(new_n592), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n593), .A2(KEYINPUT93), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n541), .A2(new_n559), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n561), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n541), .A2(new_n559), .A3(new_n562), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n593), .A2(KEYINPUT93), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n594), .A2(new_n504), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n600), .A2(new_n572), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT35), .B(G107), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G9));
  NOR2_X1   g417(.A1(new_n323), .A2(KEYINPUT36), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n318), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n333), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n332), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n503), .A2(new_n570), .A3(new_n566), .A4(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT94), .B(KEYINPUT37), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G110), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n608), .B(new_n610), .ZN(G12));
  OAI211_X1 g425(.A(new_n607), .B(new_n504), .C1(new_n563), .C2(new_n564), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT95), .B(G900), .Z(new_n614));
  AOI21_X1  g428(.A(new_n506), .B1(new_n509), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  AND4_X1   g430(.A1(new_n589), .A2(new_n588), .A3(new_n592), .A4(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n289), .A2(new_n571), .A3(new_n613), .A4(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT96), .B(G128), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G30));
  XNOR2_X1  g434(.A(new_n615), .B(KEYINPUT39), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n571), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(new_n623), .B(KEYINPUT40), .Z(new_n624));
  NOR2_X1   g438(.A1(new_n270), .A2(new_n258), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n245), .B2(new_n277), .ZN(new_n626));
  OAI21_X1  g440(.A(G472), .B1(new_n626), .B2(G902), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n266), .A2(new_n275), .A3(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n504), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n629), .A2(new_n630), .A3(new_n607), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n435), .B1(new_n384), .B2(new_n387), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n431), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n563), .A2(new_n564), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT97), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n598), .A2(KEYINPUT97), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT38), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n636), .A2(new_n637), .A3(KEYINPUT38), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n624), .A2(new_n631), .A3(new_n633), .A4(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G143), .ZN(G45));
  NOR2_X1   g458(.A1(new_n582), .A2(new_n615), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n289), .A2(new_n571), .A3(new_n613), .A4(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G146), .ZN(G48));
  NOR2_X1   g461(.A1(new_n565), .A2(new_n582), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n498), .A2(new_n499), .ZN(new_n649));
  NAND2_X1  g463(.A1(KEYINPUT98), .A2(G469), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n649), .A2(new_n263), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n263), .B1(new_n498), .B2(new_n499), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n652), .A2(KEYINPUT98), .A3(G469), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n651), .A2(new_n439), .A3(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n289), .A2(new_n648), .A3(new_n336), .A4(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT41), .B(G113), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT99), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n656), .B(new_n658), .ZN(G15));
  NAND3_X1  g473(.A1(new_n289), .A2(new_n336), .A3(new_n655), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n600), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT100), .B(G116), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G18));
  NOR2_X1   g477(.A1(new_n612), .A2(new_n654), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n388), .A2(new_n436), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n665), .A2(new_n510), .A3(new_n589), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n289), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT101), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(new_n522), .ZN(G21));
  OAI21_X1  g483(.A(new_n504), .B1(new_n563), .B2(new_n564), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n665), .A2(new_n589), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n670), .A2(new_n671), .A3(new_n654), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n261), .A2(new_n263), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n273), .B1(new_n244), .B2(new_n279), .ZN(new_n674));
  NOR2_X1   g488(.A1(G472), .A2(G902), .ZN(new_n675));
  AOI22_X1  g489(.A1(new_n673), .A2(G472), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n672), .A2(new_n336), .A3(new_n511), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G122), .ZN(G24));
  NOR2_X1   g492(.A1(new_n670), .A2(new_n654), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n645), .A2(new_n679), .A3(new_n607), .A4(new_n676), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G125), .ZN(G27));
  INV_X1    g495(.A(KEYINPUT103), .ZN(new_n682));
  AOI21_X1  g496(.A(KEYINPUT32), .B1(new_n274), .B2(new_n262), .ZN(new_n683));
  AOI22_X1  g497(.A1(new_n271), .A2(new_n272), .B1(new_n245), .B2(new_n238), .ZN(new_n684));
  NOR4_X1   g498(.A1(new_n684), .A2(new_n265), .A3(G472), .A4(G902), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n682), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n266), .A2(KEYINPUT103), .A3(new_n275), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n686), .A2(new_n288), .A3(new_n687), .ZN(new_n688));
  AOI22_X1  g502(.A1(new_n497), .A2(new_n500), .B1(G221), .B2(new_n438), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n689), .A2(new_n581), .A3(KEYINPUT42), .A4(new_n616), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT102), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n691), .B1(new_n634), .B2(new_n504), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n596), .A2(new_n691), .A3(new_n504), .A4(new_n597), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n690), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n688), .A2(new_n695), .A3(new_n336), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n289), .A2(new_n336), .ZN(new_n697));
  INV_X1    g511(.A(new_n645), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n596), .A2(new_n504), .A3(new_n597), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT102), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(new_n689), .A3(new_n693), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n697), .A2(new_n698), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n696), .B1(new_n702), .B2(KEYINPUT42), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G131), .ZN(G33));
  AND3_X1   g518(.A1(new_n700), .A2(new_n689), .A3(new_n693), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n705), .A2(new_n289), .A3(new_n336), .A4(new_n617), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G134), .ZN(G36));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n580), .A2(KEYINPUT104), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n580), .A2(KEYINPUT104), .ZN(new_n710));
  AND4_X1   g524(.A1(new_n708), .A2(new_n709), .A3(new_n632), .A4(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n665), .A2(KEYINPUT105), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n632), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n580), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n711), .B1(new_n717), .B2(KEYINPUT43), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n673), .B(new_n569), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n719), .A3(new_n607), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n692), .A2(new_n694), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n720), .A2(new_n721), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n491), .B(KEYINPUT45), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(G469), .ZN(new_n726));
  NAND2_X1  g540(.A1(G469), .A2(G902), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(KEYINPUT46), .A3(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT46), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n729), .B(G469), .C1(new_n725), .C2(G902), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n728), .A2(new_n500), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n439), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n621), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n722), .A2(new_n723), .A3(new_n724), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G137), .ZN(G39));
  INV_X1    g549(.A(new_n723), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n736), .A2(new_n289), .A3(new_n336), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT47), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n732), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n732), .A2(new_n738), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n645), .B(new_n737), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G140), .ZN(G42));
  NAND2_X1  g557(.A1(new_n688), .A2(new_n336), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n709), .A2(new_n708), .A3(new_n632), .A4(new_n710), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n580), .B1(new_n712), .B2(new_n714), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n746), .B(new_n506), .C1(new_n747), .C2(new_n708), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n736), .A2(new_n654), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n745), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(KEYINPUT48), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT50), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n676), .A2(new_n336), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n718), .A2(new_n506), .A3(new_n655), .A4(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n640), .A2(new_n641), .A3(new_n630), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n753), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n748), .A2(new_n754), .A3(new_n654), .ZN(new_n759));
  INV_X1    g573(.A(new_n757), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(new_n760), .A3(KEYINPUT50), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT116), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n750), .A2(new_n607), .A3(new_n676), .A4(new_n749), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n336), .A2(new_n506), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n665), .A2(new_n716), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n750), .A2(new_n629), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT116), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n758), .A2(new_n761), .A3(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n763), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OR3_X1    g587(.A1(new_n740), .A2(KEYINPUT114), .A3(new_n741), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n651), .A2(new_n653), .ZN(new_n775));
  XOR2_X1   g589(.A(new_n775), .B(KEYINPUT115), .Z(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n440), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT114), .B1(new_n740), .B2(new_n741), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n774), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n749), .A2(new_n755), .ZN(new_n780));
  OR3_X1    g594(.A1(new_n780), .A2(KEYINPUT113), .A3(new_n736), .ZN(new_n781));
  OAI21_X1  g595(.A(KEYINPUT113), .B1(new_n780), .B2(new_n736), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n779), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n763), .A2(KEYINPUT117), .A3(new_n768), .A4(new_n770), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n773), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n750), .A2(new_n581), .A3(new_n629), .A4(new_n765), .ZN(new_n788));
  INV_X1    g602(.A(new_n741), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n739), .A3(new_n777), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n781), .A2(new_n782), .A3(new_n790), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n791), .A2(KEYINPUT51), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n768), .A2(new_n762), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n505), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AND4_X1   g608(.A1(new_n752), .A2(new_n787), .A3(new_n788), .A4(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n588), .A2(new_n431), .A3(new_n592), .A4(new_n616), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n796), .A2(KEYINPUT108), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(KEYINPUT108), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n289), .A2(new_n797), .A3(new_n571), .A4(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n645), .A2(new_n676), .A3(new_n689), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n801), .A2(new_n607), .A3(new_n723), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n703), .A2(new_n706), .A3(new_n802), .ZN(new_n803));
  AND4_X1   g617(.A1(new_n504), .A2(new_n689), .A3(new_n633), .A4(new_n598), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n607), .A2(new_n615), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n628), .A3(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n618), .A2(new_n646), .A3(new_n806), .A4(new_n680), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n632), .A2(new_n589), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n565), .B1(new_n810), .B2(new_n582), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n811), .A2(new_n570), .A3(new_n336), .A4(new_n571), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n567), .A2(new_n812), .A3(new_n608), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(KEYINPUT107), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT107), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n567), .A2(new_n812), .A3(new_n608), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n677), .B(new_n656), .C1(new_n600), .C2(new_n660), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n668), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n803), .A2(new_n809), .A3(new_n817), .A4(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT110), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT110), .ZN(new_n824));
  INV_X1    g638(.A(new_n706), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n705), .A2(new_n289), .A3(new_n336), .A4(new_n645), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT42), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n825), .B1(new_n828), .B2(new_n696), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n819), .A2(new_n817), .A3(new_n829), .A4(new_n802), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n807), .B(KEYINPUT52), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n824), .B(new_n821), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n823), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT112), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n829), .A2(new_n802), .ZN(new_n836));
  OR3_X1    g650(.A1(new_n668), .A2(KEYINPUT111), .A3(new_n818), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT111), .B1(new_n668), .B2(new_n818), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n618), .A2(new_n680), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT109), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n841), .A2(new_n646), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n840), .A2(KEYINPUT109), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n806), .A2(KEYINPUT52), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n807), .A2(new_n808), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n839), .A2(new_n847), .A3(KEYINPUT53), .A4(new_n817), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n833), .A2(new_n834), .A3(new_n835), .A4(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n832), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n824), .B1(new_n820), .B2(new_n821), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n835), .B(new_n848), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT53), .B1(new_n845), .B2(new_n846), .ZN(new_n853));
  INV_X1    g667(.A(new_n830), .ZN(new_n854));
  AOI22_X1  g668(.A1(new_n853), .A2(new_n854), .B1(new_n820), .B2(KEYINPUT53), .ZN(new_n855));
  AOI22_X1  g669(.A1(new_n852), .A2(KEYINPUT112), .B1(KEYINPUT54), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n749), .A2(new_n755), .A3(new_n679), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n795), .A2(new_n849), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(G952), .A2(G953), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT118), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n642), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n775), .A2(KEYINPUT49), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(KEYINPUT106), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n628), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n440), .B1(new_n863), .B2(KEYINPUT106), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n630), .B1(new_n775), .B2(KEYINPUT49), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n747), .A2(new_n867), .A3(new_n336), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n862), .A2(new_n865), .A3(new_n866), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n861), .A2(new_n869), .ZN(G75));
  AOI21_X1  g684(.A(new_n263), .B1(new_n833), .B2(new_n848), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT56), .B1(new_n871), .B2(new_n561), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n535), .B1(new_n539), .B2(new_n540), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT119), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n520), .B(KEYINPUT55), .Z(new_n875));
  XNOR2_X1  g689(.A(new_n874), .B(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n876), .B1(KEYINPUT120), .B2(KEYINPUT56), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n872), .A2(new_n878), .ZN(new_n879));
  AOI211_X1 g693(.A(KEYINPUT56), .B(new_n877), .C1(new_n871), .C2(new_n561), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n319), .A2(G952), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(G51));
  OAI21_X1  g696(.A(new_n848), .B1(new_n850), .B2(new_n851), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT54), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n884), .A2(new_n885), .A3(new_n852), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n883), .A2(KEYINPUT121), .A3(KEYINPUT54), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n727), .B(KEYINPUT57), .Z(new_n888));
  NAND3_X1  g702(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n649), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT122), .ZN(new_n891));
  INV_X1    g705(.A(new_n726), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n891), .B1(new_n871), .B2(new_n892), .ZN(new_n893));
  AND4_X1   g707(.A1(new_n891), .A2(new_n883), .A3(G902), .A4(new_n892), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n881), .B1(new_n890), .B2(new_n895), .ZN(G54));
  NAND3_X1  g710(.A1(new_n871), .A2(KEYINPUT58), .A3(G475), .ZN(new_n897));
  INV_X1    g711(.A(new_n385), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n897), .A2(new_n898), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n899), .A2(new_n900), .A3(new_n881), .ZN(G60));
  XOR2_X1   g715(.A(new_n579), .B(KEYINPUT59), .Z(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n573), .B2(new_n576), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n886), .A2(new_n887), .A3(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n881), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n902), .B1(new_n856), .B2(new_n849), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n573), .A2(new_n576), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n904), .B(new_n905), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(G63));
  NAND2_X1  g723(.A1(G217), .A2(G902), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT123), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT60), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n883), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n326), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n605), .B(KEYINPUT124), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n883), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n914), .A2(new_n905), .A3(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n917), .B(new_n918), .ZN(G66));
  NAND2_X1  g733(.A1(new_n819), .A2(new_n817), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n319), .ZN(new_n921));
  OAI21_X1  g735(.A(G953), .B1(new_n508), .B2(new_n517), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n874), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n924), .B1(G898), .B2(new_n319), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n923), .B(new_n925), .ZN(G69));
  AND2_X1   g740(.A1(new_n734), .A2(new_n742), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n927), .A2(new_n843), .A3(new_n842), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n670), .A2(new_n671), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n745), .A2(new_n929), .A3(new_n733), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n829), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n319), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n255), .B(KEYINPUT125), .Z(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(new_n375), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n932), .B(new_n934), .C1(G900), .C2(new_n319), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n842), .A2(new_n643), .A3(new_n843), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT62), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n697), .B1(new_n582), .B2(new_n810), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n939), .A2(new_n571), .A3(new_n622), .A4(new_n723), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n938), .A2(new_n927), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n319), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n935), .B1(new_n934), .B2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(G900), .ZN(new_n944));
  OAI21_X1  g758(.A(G953), .B1(new_n483), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n943), .B(new_n945), .ZN(G72));
  NAND2_X1  g760(.A1(G472), .A2(G902), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT63), .Z(new_n948));
  OAI21_X1  g762(.A(new_n948), .B1(new_n941), .B2(new_n920), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n949), .A2(new_n244), .A3(new_n283), .ZN(new_n950));
  INV_X1    g764(.A(new_n283), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n928), .A2(new_n931), .A3(new_n920), .ZN(new_n952));
  INV_X1    g766(.A(new_n948), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n245), .B(new_n951), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n284), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n948), .B1(new_n955), .B2(new_n625), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT126), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n881), .B1(new_n855), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n950), .A2(new_n954), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(KEYINPUT127), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n950), .A2(new_n954), .A3(new_n961), .A4(new_n958), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n962), .ZN(G57));
endmodule


