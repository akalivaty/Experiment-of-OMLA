//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 0 1 1 1 0 0 0 1 1 0 0 1 0 0 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1243,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1305,
    new_n1306, new_n1307;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  OR3_X1    g0004(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT64), .ZN(new_n205));
  OAI21_X1  g0005(.A(KEYINPUT64), .B1(new_n203), .B2(new_n204), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  NAND2_X1  g0010(.A1(G107), .A2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n214), .B1(G50), .B2(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  INV_X1    g0017(.A(G97), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G116), .ZN(new_n221));
  INV_X1    g0021(.A(G270), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  INV_X1    g0024(.A(G250), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NOR3_X1   g0026(.A1(new_n220), .A2(new_n223), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G77), .A2(G244), .ZN(new_n228));
  AOI22_X1  g0028(.A1(new_n227), .A2(new_n228), .B1(new_n206), .B2(new_n205), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT1), .Z(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n231), .A2(new_n204), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n216), .A2(new_n212), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G50), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n210), .B(new_n230), .C1(new_n232), .C2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n217), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n222), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XNOR2_X1  g0044(.A(KEYINPUT65), .B(G107), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XOR2_X1   g0049(.A(G50), .B(G58), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(KEYINPUT70), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n203), .A2(G20), .ZN(new_n254));
  INV_X1    g0054(.A(G13), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n212), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n253), .B1(new_n257), .B2(KEYINPUT71), .ZN(new_n258));
  AOI211_X1 g0058(.A(KEYINPUT12), .B(new_n258), .C1(new_n253), .C2(new_n257), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(KEYINPUT12), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G50), .ZN(new_n262));
  INV_X1    g0062(.A(G77), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n204), .A2(G33), .ZN(new_n264));
  OAI221_X1 g0064(.A(new_n262), .B1(new_n204), .B2(G68), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n231), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n265), .A2(KEYINPUT11), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n267), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(new_n254), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n260), .B(new_n268), .C1(new_n212), .C2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(KEYINPUT11), .B1(new_n265), .B2(new_n267), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n259), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT72), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT14), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n203), .B(G274), .C1(G41), .C2(G45), .ZN(new_n278));
  XOR2_X1   g0078(.A(new_n278), .B(KEYINPUT69), .Z(new_n279));
  INV_X1    g0079(.A(G33), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  OAI211_X1 g0081(.A(G1), .B(G13), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n280), .A2(new_n218), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT66), .B(G1698), .ZN(new_n286));
  INV_X1    g0086(.A(G226), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  OAI22_X1  g0088(.A1(new_n286), .A2(new_n287), .B1(new_n217), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT3), .B(G33), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n285), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n279), .B1(new_n213), .B2(new_n284), .C1(new_n291), .C2(new_n282), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT13), .ZN(new_n293));
  OR2_X1    g0093(.A1(new_n291), .A2(new_n282), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT13), .ZN(new_n295));
  INV_X1    g0095(.A(new_n284), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G238), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n294), .A2(new_n295), .A3(new_n297), .A4(new_n279), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n277), .B1(new_n299), .B2(G169), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G169), .ZN(new_n302));
  AOI211_X1 g0102(.A(new_n302), .B(new_n276), .C1(new_n293), .C2(new_n298), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n299), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G179), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n301), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT73), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT73), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n301), .A2(new_n309), .A3(new_n304), .A4(new_n306), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n273), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G200), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n305), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G190), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n273), .B1(new_n299), .B2(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT8), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n216), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT68), .B(G58), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(new_n319), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(new_n270), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n323), .B1(new_n256), .B2(new_n322), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n280), .A2(KEYINPUT3), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT3), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G33), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT7), .B1(new_n329), .B2(new_n204), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT7), .ZN(new_n331));
  AOI211_X1 g0131(.A(new_n331), .B(G20), .C1(new_n326), .C2(new_n328), .ZN(new_n332));
  OAI21_X1  g0132(.A(G68), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n233), .B1(new_n321), .B2(new_n212), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n334), .A2(G20), .B1(G159), .B2(new_n261), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT16), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n269), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT74), .ZN(new_n339));
  AND3_X1   g0139(.A1(new_n326), .A2(new_n328), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n339), .B1(new_n326), .B2(new_n328), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n204), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n332), .B1(new_n342), .B2(new_n331), .ZN(new_n343));
  OAI211_X1 g0143(.A(KEYINPUT16), .B(new_n335), .C1(new_n343), .C2(new_n212), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n325), .B1(new_n338), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n278), .B1(new_n284), .B2(new_n217), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  XOR2_X1   g0147(.A(KEYINPUT76), .B(G190), .Z(new_n348));
  INV_X1    g0148(.A(G223), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n286), .A2(new_n349), .B1(new_n287), .B2(new_n288), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n350), .A2(new_n290), .B1(G33), .B2(G87), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n347), .B(new_n348), .C1(new_n351), .C2(new_n282), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT77), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n288), .A2(KEYINPUT66), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT66), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G1698), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n349), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n287), .A2(new_n288), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n290), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G33), .A2(G87), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n231), .B1(G33), .B2(G41), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT77), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n363), .A2(new_n364), .A3(new_n347), .A4(new_n348), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n282), .B1(new_n359), .B2(new_n360), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n312), .B1(new_n366), .B2(new_n346), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n353), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  AND2_X1   g0168(.A1(new_n345), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g0169(.A(new_n369), .B(KEYINPUT17), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n338), .A2(new_n344), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n324), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n363), .A2(G179), .A3(new_n347), .ZN(new_n373));
  OAI21_X1  g0173(.A(G169), .B1(new_n366), .B2(new_n346), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n372), .A2(KEYINPUT18), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT75), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n372), .A2(new_n375), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT18), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n379), .A2(new_n377), .A3(new_n380), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n370), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n354), .A2(new_n356), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G222), .ZN(new_n386));
  XOR2_X1   g0186(.A(KEYINPUT67), .B(G223), .Z(new_n387));
  OAI211_X1 g0187(.A(new_n386), .B(new_n290), .C1(new_n288), .C2(new_n387), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n388), .B(new_n362), .C1(G77), .C2(new_n290), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n296), .A2(G226), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n389), .A2(new_n390), .A3(new_n278), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G200), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT9), .ZN(new_n393));
  INV_X1    g0193(.A(G50), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n394), .A2(new_n216), .A3(new_n212), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n395), .A2(G20), .B1(G150), .B2(new_n261), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n322), .B2(new_n264), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n397), .A2(new_n267), .B1(new_n394), .B2(new_n256), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(new_n394), .B2(new_n270), .ZN(new_n399));
  OAI221_X1 g0199(.A(new_n392), .B1(new_n314), .B2(new_n391), .C1(new_n393), .C2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n400), .B1(new_n393), .B2(new_n399), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT10), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n401), .B(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n391), .A2(new_n302), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n404), .B(new_n399), .C1(G179), .C2(new_n391), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n270), .A2(new_n263), .ZN(new_n406));
  XOR2_X1   g0206(.A(KEYINPUT8), .B(G58), .Z(new_n407));
  AOI22_X1  g0207(.A1(new_n407), .A2(new_n261), .B1(G20), .B2(G77), .ZN(new_n408));
  XOR2_X1   g0208(.A(KEYINPUT15), .B(G87), .Z(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n408), .B1(new_n264), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n406), .B1(new_n411), .B2(new_n267), .ZN(new_n412));
  INV_X1    g0212(.A(new_n256), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n412), .B1(G77), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n278), .ZN(new_n415));
  INV_X1    g0215(.A(G244), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n284), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(G107), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n282), .B1(new_n329), .B2(new_n418), .ZN(new_n419));
  OAI221_X1 g0219(.A(new_n290), .B1(new_n213), .B2(new_n288), .C1(new_n286), .C2(new_n217), .ZN(new_n420));
  AOI211_X1 g0220(.A(new_n415), .B(new_n417), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(G179), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n414), .B(new_n423), .C1(G169), .C2(new_n421), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n384), .A2(new_n403), .A3(new_n405), .A4(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n414), .B1(G190), .B2(new_n421), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n312), .B2(new_n421), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n318), .A2(new_n425), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(G45), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n431), .A2(G1), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT5), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(G41), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n281), .A2(KEYINPUT5), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n432), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n436), .A2(G257), .A3(new_n282), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT82), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT82), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n436), .A2(new_n439), .A3(G257), .A4(new_n282), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n435), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n362), .A2(new_n442), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n432), .A2(KEYINPUT81), .A3(new_n434), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT81), .B1(new_n432), .B2(new_n434), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n443), .B(G274), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(KEYINPUT83), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n385), .A2(new_n290), .A3(G244), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT80), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT4), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT4), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n449), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n225), .A2(new_n288), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n290), .A2(new_n455), .B1(G33), .B2(G283), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n452), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n362), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT83), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n441), .A2(new_n459), .A3(new_n446), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n448), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G169), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n441), .A2(new_n459), .A3(new_n446), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n459), .B1(new_n441), .B2(new_n446), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n465), .A2(G179), .A3(new_n458), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n331), .B1(new_n290), .B2(G20), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n329), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G107), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT79), .ZN(new_n472));
  AND2_X1   g0272(.A1(KEYINPUT78), .A2(G97), .ZN(new_n473));
  NOR2_X1   g0273(.A1(KEYINPUT78), .A2(G97), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n475), .A2(KEYINPUT6), .A3(new_n418), .ZN(new_n476));
  XOR2_X1   g0276(.A(G97), .B(G107), .Z(new_n477));
  OAI21_X1  g0277(.A(new_n476), .B1(KEYINPUT6), .B2(new_n477), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n478), .A2(G20), .B1(G77), .B2(new_n261), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT79), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n470), .A2(new_n480), .A3(G107), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n472), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n267), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n256), .A2(new_n218), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n203), .A2(G33), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n413), .A2(new_n269), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G97), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n483), .A2(new_n484), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT84), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT84), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n483), .A2(new_n491), .A3(new_n484), .A4(new_n488), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n467), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n483), .A2(new_n484), .A3(new_n488), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n461), .A2(G200), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n494), .B(new_n495), .C1(new_n314), .C2(new_n461), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n290), .A2(new_n204), .A3(G87), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT22), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT22), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n290), .A2(new_n499), .A3(new_n204), .A4(G87), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n280), .A2(new_n221), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n498), .A2(new_n500), .B1(new_n204), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n204), .A2(G107), .ZN(new_n503));
  XNOR2_X1  g0303(.A(new_n503), .B(KEYINPUT23), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT24), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n502), .A2(KEYINPUT24), .A3(new_n504), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(new_n267), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n256), .A2(new_n418), .ZN(new_n510));
  XNOR2_X1  g0310(.A(new_n510), .B(KEYINPUT25), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n487), .A2(G107), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n436), .A2(G264), .A3(new_n282), .ZN(new_n515));
  OAI22_X1  g0315(.A1(new_n286), .A2(new_n225), .B1(new_n219), .B2(new_n288), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n516), .A2(new_n290), .B1(G33), .B2(G294), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n515), .B1(new_n517), .B2(new_n282), .ZN(new_n518));
  INV_X1    g0318(.A(new_n446), .ZN(new_n519));
  OAI21_X1  g0319(.A(G200), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n518), .A2(new_n519), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G190), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n513), .A2(new_n514), .A3(new_n520), .A4(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n493), .A2(new_n496), .A3(new_n523), .ZN(new_n524));
  OAI22_X1  g0324(.A1(new_n286), .A2(new_n213), .B1(new_n416), .B2(new_n288), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n290), .ZN(new_n526));
  INV_X1    g0326(.A(new_n501), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n282), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(G274), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n432), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n225), .B1(new_n431), .B2(G1), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(new_n282), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(KEYINPUT85), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT85), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n501), .B1(new_n525), .B2(new_n290), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n535), .B(new_n532), .C1(new_n536), .C2(new_n282), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n290), .A2(new_n204), .A3(G68), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT78), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n218), .ZN(new_n542));
  NAND2_X1  g0342(.A1(KEYINPUT78), .A2(G97), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n544), .A2(new_n264), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n544), .A2(new_n224), .A3(new_n418), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(G20), .B1(new_n285), .B2(KEYINPUT19), .ZN(new_n548));
  OAI221_X1 g0348(.A(new_n540), .B1(KEYINPUT19), .B2(new_n545), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n549), .A2(new_n267), .B1(new_n256), .B2(new_n410), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n487), .A2(new_n409), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n539), .A2(new_n302), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n538), .A2(new_n422), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT86), .ZN(new_n554));
  AOI211_X1 g0354(.A(KEYINPUT86), .B(G179), .C1(new_n534), .C2(new_n537), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n552), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n487), .A2(G87), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n550), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(G190), .B2(new_n538), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n539), .A2(G200), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n521), .A2(G169), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n564), .B1(new_n422), .B2(new_n521), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n509), .A2(new_n514), .A3(new_n512), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NOR3_X1   g0368(.A1(new_n524), .A2(new_n563), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n256), .A2(new_n221), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n413), .A2(G116), .A3(new_n269), .A4(new_n485), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n542), .A2(new_n280), .A3(new_n543), .ZN(new_n572));
  AOI21_X1  g0372(.A(G20), .B1(G33), .B2(G283), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n266), .A2(new_n231), .B1(G20), .B2(new_n221), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n574), .A2(KEYINPUT20), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT20), .B1(new_n574), .B2(new_n575), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n570), .B(new_n571), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT88), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT20), .ZN(new_n580));
  INV_X1    g0380(.A(new_n573), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n475), .B2(new_n280), .ZN(new_n582));
  INV_X1    g0382(.A(new_n575), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n580), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n574), .A2(KEYINPUT20), .A3(new_n575), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT88), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n586), .A2(new_n587), .A3(new_n570), .A4(new_n571), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n579), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n436), .A2(G270), .A3(new_n282), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n446), .A2(KEYINPUT87), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT87), .B1(new_n446), .B2(new_n590), .ZN(new_n592));
  AND2_X1   g0392(.A1(G264), .A2(G1698), .ZN(new_n593));
  AOI211_X1 g0393(.A(new_n593), .B(new_n329), .C1(G257), .C2(new_n385), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n362), .B1(new_n290), .B2(G303), .ZN(new_n595));
  OAI22_X1  g0395(.A1(new_n591), .A2(new_n592), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n589), .A2(KEYINPUT21), .A3(G169), .A4(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT89), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n594), .A2(new_n595), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n446), .A2(new_n590), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT87), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n446), .A2(KEYINPUT87), .A3(new_n590), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n600), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n605), .A2(new_n302), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n606), .A2(KEYINPUT89), .A3(KEYINPUT21), .A4(new_n589), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n589), .A2(G179), .A3(new_n605), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT90), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n589), .A2(KEYINPUT90), .A3(G179), .A4(new_n605), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n599), .A2(new_n607), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT91), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT21), .B1(new_n606), .B2(new_n589), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n599), .A2(new_n607), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n610), .A2(new_n611), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n615), .B1(new_n618), .B2(KEYINPUT91), .ZN(new_n619));
  INV_X1    g0419(.A(new_n589), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n596), .A2(G200), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n620), .B(new_n621), .C1(new_n348), .C2(new_n596), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n569), .A2(new_n614), .A3(new_n619), .A4(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n430), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g0424(.A(new_n624), .B(KEYINPUT92), .Z(G372));
  INV_X1    g0425(.A(new_n370), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n316), .A2(new_n424), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n626), .B1(new_n311), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n381), .A2(new_n376), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n403), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n631), .A2(new_n405), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT26), .ZN(new_n633));
  INV_X1    g0433(.A(new_n528), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n532), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(G200), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n560), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT93), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n467), .A2(new_n638), .A3(new_n489), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n638), .B1(new_n467), .B2(new_n489), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n633), .B(new_n637), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n550), .A2(new_n551), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n635), .A2(new_n302), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n553), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n615), .ZN(new_n645));
  AND4_X1   g0445(.A1(new_n616), .A2(new_n617), .A3(new_n645), .A4(new_n567), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n493), .A2(new_n496), .A3(new_n523), .A4(new_n637), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n641), .B(new_n644), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n563), .A2(new_n493), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(new_n633), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n632), .B1(new_n430), .B2(new_n652), .ZN(G369));
  NOR2_X1   g0453(.A1(new_n255), .A2(G20), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  OR3_X1    g0455(.A1(new_n655), .A2(KEYINPUT27), .A3(G1), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT27), .B1(new_n655), .B2(G1), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(G213), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(G343), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n567), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n566), .A2(new_n660), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n523), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n661), .B1(new_n567), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT94), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n664), .B(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n660), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n620), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n618), .B2(new_n615), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n619), .A2(new_n614), .A3(new_n622), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n669), .B1(new_n670), .B2(new_n668), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(G330), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n645), .B1(new_n612), .B2(new_n613), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n618), .A2(KEYINPUT91), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(new_n660), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n666), .B1(new_n673), .B2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n661), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(G399));
  INV_X1    g0480(.A(new_n208), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(G41), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n546), .A2(G116), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G1), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n234), .B2(new_n683), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT28), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n651), .A2(new_n667), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT29), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT86), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n538), .B2(new_n422), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(new_n555), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n693), .A2(new_n552), .B1(new_n561), .B2(new_n560), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n490), .A2(new_n492), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n694), .A2(new_n633), .A3(new_n467), .A4(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n644), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n618), .A2(KEYINPUT91), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n698), .A2(new_n614), .A3(new_n645), .A4(new_n567), .ZN(new_n699));
  INV_X1    g0499(.A(new_n647), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n697), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT26), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n660), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT29), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n690), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(G330), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n465), .A2(new_n605), .A3(G179), .A4(new_n458), .ZN(new_n709));
  INV_X1    g0509(.A(new_n518), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n538), .A2(new_n710), .ZN(new_n711));
  OAI211_X1 g0511(.A(KEYINPUT95), .B(new_n708), .C1(new_n709), .C2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n711), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n461), .A2(new_n422), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n708), .A2(KEYINPUT95), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n713), .A2(new_n714), .A3(new_n605), .A4(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n605), .A2(new_n521), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n717), .A2(new_n422), .A3(new_n461), .A4(new_n635), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n712), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(KEYINPUT31), .B1(new_n719), .B2(new_n660), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n660), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n720), .B1(KEYINPUT96), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n719), .A2(new_n660), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(KEYINPUT96), .A3(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n676), .A2(new_n622), .A3(new_n569), .A4(new_n667), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n707), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n706), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n687), .B1(new_n732), .B2(G1), .ZN(G364));
  NOR2_X1   g0533(.A1(G13), .A2(G33), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G20), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n671), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n681), .A2(new_n329), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G355), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n340), .A2(new_n341), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n681), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(G45), .B2(new_n234), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n251), .A2(G45), .ZN(new_n745));
  OAI221_X1 g0545(.A(new_n740), .B1(G116), .B2(new_n208), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n204), .B1(KEYINPUT97), .B2(new_n302), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n302), .A2(KEYINPUT97), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n231), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n736), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n203), .B1(new_n654), .B2(G45), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n682), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n204), .A2(new_n422), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n312), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n348), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT98), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n348), .A2(new_n756), .A3(KEYINPUT98), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n755), .A2(new_n314), .A3(new_n312), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n761), .A2(new_n321), .B1(new_n263), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n755), .A2(G200), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n348), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G179), .A2(G200), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n204), .B1(new_n767), .B2(G190), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n766), .A2(new_n394), .B1(new_n218), .B2(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n204), .A2(new_n312), .A3(G179), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(new_n314), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G107), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n764), .A2(G190), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n773), .B1(new_n775), .B2(new_n212), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n763), .A2(new_n769), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n770), .A2(G190), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G87), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n767), .A2(G20), .A3(new_n314), .ZN(new_n781));
  INV_X1    g0581(.A(G159), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT32), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n777), .A2(new_n290), .A3(new_n780), .A4(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G322), .ZN(new_n786));
  XOR2_X1   g0586(.A(KEYINPUT33), .B(G317), .Z(new_n787));
  OAI22_X1  g0587(.A1(new_n761), .A2(new_n786), .B1(new_n775), .B2(new_n787), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n788), .B(KEYINPUT99), .Z(new_n789));
  INV_X1    g0589(.A(G283), .ZN(new_n790));
  INV_X1    g0590(.A(G311), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n771), .A2(new_n790), .B1(new_n762), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n781), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n290), .B(new_n792), .C1(G329), .C2(new_n793), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n789), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G294), .ZN(new_n796));
  INV_X1    g0596(.A(G303), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n795), .B1(new_n796), .B2(new_n768), .C1(new_n797), .C2(new_n778), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n765), .A2(G326), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n785), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n749), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n738), .A2(new_n751), .A3(new_n754), .A4(new_n801), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n671), .A2(G330), .ZN(new_n803));
  INV_X1    g0603(.A(new_n754), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n803), .A2(new_n672), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n802), .A2(new_n805), .ZN(G396));
  AND2_X1   g0606(.A1(new_n414), .A2(new_n660), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n424), .B1(new_n428), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n424), .A2(new_n660), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT103), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n688), .A2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT104), .Z(new_n814));
  INV_X1    g0614(.A(new_n811), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n667), .B(new_n815), .C1(new_n648), .C2(new_n650), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n730), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n814), .A2(new_n729), .A3(new_n816), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n818), .A2(new_n804), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n778), .A2(new_n418), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n772), .A2(G87), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n791), .B2(new_n781), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(G283), .B2(new_n774), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n797), .B2(new_n766), .ZN(new_n825));
  INV_X1    g0625(.A(new_n762), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n821), .B(new_n825), .C1(G116), .C2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n768), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n290), .B1(new_n828), .B2(G97), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n827), .B(new_n829), .C1(new_n796), .C2(new_n761), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT101), .Z(new_n831));
  NOR2_X1   g0631(.A1(new_n768), .A2(new_n321), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G137), .A2(new_n765), .B1(new_n774), .B2(G150), .ZN(new_n833));
  INV_X1    g0633(.A(G143), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n833), .B1(new_n782), .B2(new_n762), .C1(new_n761), .C2(new_n834), .ZN(new_n835));
  XOR2_X1   g0635(.A(KEYINPUT102), .B(KEYINPUT34), .Z(new_n836));
  OR2_X1    g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n772), .A2(G68), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n835), .A2(new_n836), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n741), .B1(G132), .B2(new_n793), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n837), .A2(new_n838), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n832), .B(new_n841), .C1(G50), .C2(new_n779), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n749), .B1(new_n831), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n749), .A2(new_n734), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT100), .Z(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n804), .B1(new_n846), .B2(new_n263), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n843), .B(new_n847), .C1(new_n735), .C2(new_n815), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n820), .A2(new_n848), .ZN(G384));
  OAI21_X1  g0649(.A(new_n335), .B1(new_n343), .B2(new_n212), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n337), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n851), .A2(new_n267), .A3(new_n344), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n324), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n375), .ZN(new_n854));
  INV_X1    g0654(.A(new_n658), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n345), .A2(new_n368), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(KEYINPUT37), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n369), .A2(KEYINPUT37), .ZN(new_n860));
  OR3_X1    g0660(.A1(new_n345), .A2(KEYINPUT105), .A3(new_n658), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT105), .B1(new_n345), .B2(new_n658), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n860), .A2(new_n863), .A3(new_n379), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n865), .B(KEYINPUT38), .C1(new_n384), .C2(new_n856), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT106), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n345), .A2(new_n368), .A3(new_n867), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n373), .A2(new_n374), .ZN(new_n869));
  OAI21_X1  g0669(.A(KEYINPUT106), .B1(new_n345), .B2(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(KEYINPUT107), .B(new_n868), .C1(new_n369), .C2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n863), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n379), .A2(KEYINPUT106), .A3(new_n857), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT107), .B1(new_n873), .B2(new_n868), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT37), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n875), .A2(KEYINPUT108), .A3(new_n864), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT108), .B1(new_n875), .B2(new_n864), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n863), .B1(new_n626), .B2(new_n629), .ZN(new_n878));
  NOR3_X1   g0678(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n866), .B1(new_n879), .B2(KEYINPUT38), .ZN(new_n880));
  OR2_X1    g0680(.A1(new_n273), .A2(new_n667), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n317), .A2(new_n881), .B1(new_n311), .B2(new_n660), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n882), .A2(new_n811), .ZN(new_n883));
  INV_X1    g0683(.A(new_n720), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n728), .A2(new_n884), .A3(new_n721), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n880), .A2(KEYINPUT40), .A3(new_n883), .A4(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n865), .B1(new_n384), .B2(new_n856), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT38), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n866), .ZN(new_n890));
  INV_X1    g0690(.A(new_n311), .ZN(new_n891));
  INV_X1    g0691(.A(new_n316), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n891), .A2(new_n892), .A3(new_n881), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n311), .A2(new_n660), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n885), .A2(new_n890), .A3(new_n895), .A4(new_n815), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT40), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n886), .A2(new_n429), .A3(new_n898), .A4(new_n885), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n886), .A2(G330), .A3(new_n898), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n885), .A2(G330), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n430), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n899), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n311), .A2(new_n667), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n889), .A2(KEYINPUT39), .A3(new_n866), .ZN(new_n906));
  INV_X1    g0706(.A(new_n866), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n875), .A2(new_n864), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT108), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n878), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n875), .A2(KEYINPUT108), .A3(new_n864), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n907), .B1(new_n913), .B2(new_n888), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n905), .B(new_n906), .C1(new_n914), .C2(KEYINPUT39), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n629), .A2(new_n855), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n882), .B1(new_n810), .B2(new_n816), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n916), .B1(new_n917), .B2(new_n890), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  XOR2_X1   g0719(.A(new_n903), .B(new_n919), .Z(new_n920));
  NAND3_X1  g0720(.A1(new_n690), .A2(new_n429), .A3(new_n705), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n632), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n920), .B(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n203), .B2(new_n654), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n221), .B1(new_n478), .B2(KEYINPUT35), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n925), .B(new_n232), .C1(KEYINPUT35), .C2(new_n478), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT36), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n235), .B1(new_n321), .B2(new_n212), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n928), .A2(new_n263), .B1(G50), .B2(new_n212), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(G1), .A3(new_n255), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n924), .A2(new_n927), .A3(new_n930), .ZN(G367));
  OAI221_X1 g0731(.A(new_n741), .B1(new_n544), .B2(new_n771), .C1(new_n766), .C2(new_n791), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n778), .A2(new_n221), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n933), .A2(KEYINPUT46), .B1(G317), .B2(new_n793), .ZN(new_n934));
  OAI221_X1 g0734(.A(new_n934), .B1(KEYINPUT46), .B2(new_n933), .C1(new_n790), .C2(new_n762), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n932), .B(new_n935), .C1(G107), .C2(new_n828), .ZN(new_n936));
  OAI221_X1 g0736(.A(new_n936), .B1(new_n796), .B2(new_n775), .C1(new_n797), .C2(new_n761), .ZN(new_n937));
  INV_X1    g0737(.A(G150), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n761), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n778), .A2(new_n321), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n771), .A2(new_n263), .ZN(new_n941));
  AOI211_X1 g0741(.A(new_n940), .B(new_n941), .C1(G143), .C2(new_n765), .ZN(new_n942));
  INV_X1    g0742(.A(G137), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n762), .A2(new_n394), .B1(new_n943), .B2(new_n781), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n329), .B(new_n944), .C1(G159), .C2(new_n774), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n828), .A2(G68), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n942), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n937), .B1(new_n939), .B2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT47), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n749), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n559), .A2(new_n660), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n637), .A2(new_n644), .A3(new_n951), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n644), .A2(new_n951), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n952), .A2(new_n736), .A3(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n743), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n750), .B1(new_n208), .B2(new_n410), .C1(new_n955), .C2(new_n243), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n950), .A2(new_n754), .A3(new_n954), .A4(new_n956), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n493), .A2(new_n496), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n489), .A2(new_n660), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n666), .A2(new_n677), .A3(new_n958), .A4(new_n959), .ZN(new_n960));
  OR3_X1    g0760(.A1(new_n960), .A2(KEYINPUT109), .A3(KEYINPUT42), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n958), .A2(new_n959), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n467), .A2(new_n489), .A3(new_n660), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n568), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n660), .B1(new_n965), .B2(new_n493), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(new_n960), .B2(KEYINPUT42), .ZN(new_n967));
  OAI21_X1  g0767(.A(KEYINPUT109), .B1(new_n960), .B2(KEYINPUT42), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n961), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n952), .A2(new_n953), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT110), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n969), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n972), .B1(new_n969), .B2(new_n974), .ZN(new_n977));
  INV_X1    g0777(.A(new_n666), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n672), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n964), .ZN(new_n980));
  NOR3_X1   g0780(.A1(new_n976), .A2(new_n977), .A3(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n980), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n969), .A2(new_n974), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n971), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n982), .B1(new_n984), .B2(new_n975), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n666), .A2(new_n677), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n987), .A2(new_n679), .A3(new_n964), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(KEYINPUT111), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT111), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n987), .A2(new_n990), .A3(new_n679), .A4(new_n964), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT45), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n964), .B1(new_n987), .B2(new_n679), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT44), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n989), .A2(KEYINPUT45), .A3(new_n991), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n994), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n672), .B(new_n978), .C1(new_n676), .C2(new_n660), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n678), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n731), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n682), .B(KEYINPUT41), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n752), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  AND3_X1   g0804(.A1(new_n986), .A2(new_n1004), .A3(KEYINPUT112), .ZN(new_n1005));
  AOI21_X1  g0805(.A(KEYINPUT112), .B1(new_n986), .B2(new_n1004), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n957), .B1(new_n1005), .B2(new_n1006), .ZN(G387));
  NAND2_X1  g0807(.A1(new_n732), .A2(new_n1000), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n678), .A2(new_n999), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n731), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1008), .A2(new_n682), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1000), .A2(new_n753), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n322), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n1013), .A2(new_n774), .B1(new_n826), .B2(G68), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT113), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n742), .B1(new_n761), .B2(new_n394), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n779), .A2(G77), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1017), .B1(new_n938), .B2(new_n781), .C1(new_n766), .C2(new_n782), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n218), .B2(new_n771), .C1(new_n410), .C2(new_n768), .ZN(new_n1020));
  INV_X1    g0820(.A(G317), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n761), .A2(new_n1021), .B1(new_n797), .B2(new_n762), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT114), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n791), .B2(new_n775), .C1(new_n786), .C2(new_n766), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT48), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n828), .A2(G283), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n779), .A2(G294), .ZN(new_n1027));
  AND3_X1   g0827(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(KEYINPUT49), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n793), .A2(G326), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n772), .A2(G116), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1029), .A2(new_n741), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1028), .A2(KEYINPUT49), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1020), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n749), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n978), .A2(new_n736), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n955), .B1(new_n240), .B2(G45), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n684), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1037), .B1(new_n1038), .B2(new_n739), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n407), .ZN(new_n1040));
  OR3_X1    g0840(.A1(new_n1040), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1041));
  OAI21_X1  g0841(.A(KEYINPUT50), .B1(new_n1040), .B2(G50), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1041), .A2(new_n431), .A3(new_n1042), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1038), .B(new_n1043), .C1(G68), .C2(G77), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n1039), .A2(new_n1044), .B1(G107), .B2(new_n208), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n804), .B1(new_n1045), .B2(new_n750), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1035), .A2(new_n1036), .A3(new_n1046), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1012), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1011), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(KEYINPUT115), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT115), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1011), .A2(new_n1048), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1052), .ZN(G393));
  INV_X1    g0853(.A(new_n749), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n761), .A2(new_n791), .B1(new_n1021), .B2(new_n766), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT52), .Z(new_n1056));
  NOR2_X1   g0856(.A1(new_n768), .A2(new_n221), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n773), .B1(new_n796), .B2(new_n762), .C1(new_n790), .C2(new_n778), .ZN(new_n1058));
  NOR4_X1   g0858(.A1(new_n1056), .A2(new_n290), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1059), .B1(new_n797), .B2(new_n775), .C1(new_n786), .C2(new_n781), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n822), .B1(new_n1040), .B2(new_n762), .C1(new_n394), .C2(new_n775), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n742), .B1(new_n834), .B2(new_n781), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n778), .A2(new_n212), .B1(new_n263), .B2(new_n768), .ZN(new_n1063));
  NOR3_X1   g0863(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n761), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n1065), .A2(G159), .B1(G150), .B2(new_n765), .ZN(new_n1066));
  XOR2_X1   g0866(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1064), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT117), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1054), .B1(new_n1060), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n750), .B1(new_n208), .B2(new_n544), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n248), .B2(new_n743), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n1073), .A2(new_n804), .A3(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n737), .B2(new_n964), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n998), .A2(new_n979), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n979), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n994), .A2(new_n996), .A3(new_n997), .A4(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1077), .B1(new_n1081), .B2(new_n752), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n998), .A2(new_n732), .A3(new_n1000), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n1081), .B2(new_n1008), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1082), .B1(new_n1084), .B2(new_n682), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(G390));
  OAI21_X1  g0886(.A(new_n882), .B1(new_n901), .B2(new_n812), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n809), .B1(new_n704), .B2(new_n808), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n729), .A2(new_n815), .A3(new_n895), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT119), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n623), .A2(new_n660), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n721), .A2(KEYINPUT96), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n884), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n725), .ZN(new_n1095));
  OAI211_X1 g0895(.A(G330), .B(new_n815), .C1(new_n1092), .C2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n882), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n885), .A2(new_n895), .A3(G330), .A4(new_n815), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n816), .A2(new_n810), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1091), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1100), .ZN(new_n1102));
  AOI211_X1 g0902(.A(KEYINPUT119), .B(new_n1102), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1090), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n922), .A2(new_n902), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n906), .B1(new_n914), .B2(KEYINPUT39), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n904), .B1(new_n1102), .B2(new_n882), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n904), .B(KEYINPUT118), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1110), .B(new_n880), .C1(new_n1088), .C2(new_n882), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1089), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n1109), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1098), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1106), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n906), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT39), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1118), .B1(new_n880), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n917), .A2(new_n905), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1111), .B(new_n1112), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n699), .A2(new_n700), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n697), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1123), .A2(new_n703), .A3(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1125), .A2(new_n667), .A3(new_n808), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n810), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n914), .B1(new_n1127), .B2(new_n895), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1128), .A2(new_n1110), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1122), .B1(new_n1129), .B2(new_n1114), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1130), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1117), .A2(new_n682), .A3(new_n1131), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1065), .A2(G116), .B1(G77), .B2(new_n828), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n772), .A2(G68), .B1(new_n826), .B2(new_n475), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n329), .B1(new_n775), .B2(new_n418), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G294), .B2(new_n793), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1133), .A2(new_n780), .A3(new_n1134), .A4(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(G283), .B2(new_n765), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n290), .B1(new_n771), .B2(new_n394), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT120), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1139), .A2(new_n1140), .B1(G137), .B2(new_n774), .ZN(new_n1141));
  INV_X1    g0941(.A(G128), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1141), .B1(new_n1140), .B2(new_n1139), .C1(new_n1142), .C2(new_n766), .ZN(new_n1143));
  XOR2_X1   g0943(.A(KEYINPUT54), .B(G143), .Z(new_n1144));
  AOI22_X1  g0944(.A1(new_n826), .A2(new_n1144), .B1(new_n828), .B2(G159), .ZN(new_n1145));
  OAI21_X1  g0945(.A(KEYINPUT53), .B1(new_n778), .B2(new_n938), .ZN(new_n1146));
  INV_X1    g0946(.A(G132), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1145), .B(new_n1146), .C1(new_n761), .C2(new_n1147), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n778), .A2(KEYINPUT53), .A3(new_n938), .ZN(new_n1149));
  INV_X1    g0949(.A(G125), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n781), .A2(new_n1150), .ZN(new_n1151));
  NOR4_X1   g0951(.A1(new_n1143), .A2(new_n1148), .A3(new_n1149), .A4(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n749), .B1(new_n1138), .B2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1153), .B(new_n754), .C1(new_n1013), .C2(new_n845), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(new_n1107), .B2(new_n734), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(new_n1130), .B2(new_n753), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1132), .A2(new_n1156), .ZN(G378));
  INV_X1    g0957(.A(new_n1090), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(KEYINPUT119), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1099), .A2(new_n1091), .A3(new_n1100), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1158), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1105), .B1(new_n1116), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n886), .A2(G330), .A3(new_n898), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n403), .A2(new_n405), .ZN(new_n1165));
  XOR2_X1   g0965(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1166));
  XNOR2_X1  g0966(.A(new_n1165), .B(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n399), .A2(new_n855), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1167), .B(new_n1168), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n915), .A2(new_n918), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1169), .B1(new_n915), .B2(new_n918), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1164), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1169), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n919), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n915), .A2(new_n918), .A3(new_n1169), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1174), .A2(new_n900), .A3(new_n1175), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n1172), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1163), .A2(KEYINPUT57), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT57), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1105), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n1130), .B2(new_n1104), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1172), .A2(new_n1176), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1179), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1178), .A2(new_n682), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1177), .A2(new_n753), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n804), .B1(new_n846), .B2(new_n394), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n762), .A2(new_n943), .B1(new_n768), .B2(new_n938), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n775), .A2(new_n1147), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1187), .B(new_n1188), .C1(new_n779), .C2(new_n1144), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1189), .B1(new_n1150), .B2(new_n766), .C1(new_n1142), .C2(new_n761), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1191), .A2(G33), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n772), .A2(G159), .ZN(new_n1194));
  AOI21_X1  g0994(.A(G41), .B1(new_n793), .B2(G124), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n742), .A2(G33), .ZN(new_n1197));
  AOI21_X1  g0997(.A(G50), .B1(new_n1197), .B2(new_n281), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT121), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n771), .A2(new_n321), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n410), .A2(new_n762), .B1(new_n790), .B2(new_n781), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(G97), .C2(new_n774), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n765), .A2(G116), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1202), .A2(new_n946), .A3(new_n1017), .A4(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n281), .B1(new_n761), .B2(new_n418), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n1204), .A2(new_n742), .A3(new_n1205), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT58), .Z(new_n1207));
  AND3_X1   g1007(.A1(new_n1196), .A2(new_n1199), .A3(new_n1207), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1186), .B1(new_n1054), .B2(new_n1208), .C1(new_n1173), .C2(new_n735), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1185), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1184), .A2(new_n1210), .ZN(G375));
  NAND2_X1  g1011(.A1(new_n1162), .A2(new_n1180), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1212), .A2(new_n1106), .A3(new_n1002), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n766), .A2(new_n796), .B1(new_n410), .B2(new_n768), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n775), .A2(new_n221), .B1(new_n762), .B2(new_n418), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT122), .Z(new_n1216));
  AOI211_X1 g1016(.A(new_n1214), .B(new_n1216), .C1(G283), .C2(new_n1065), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n218), .B2(new_n778), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n781), .A2(new_n797), .ZN(new_n1219));
  NOR4_X1   g1019(.A1(new_n1218), .A2(new_n290), .A3(new_n941), .A4(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1065), .A2(G137), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n774), .A2(new_n1144), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n762), .A2(new_n938), .B1(new_n768), .B2(new_n394), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1223), .B(new_n741), .C1(G132), .C2(new_n765), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n771), .A2(new_n321), .B1(new_n1142), .B2(new_n781), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1221), .A2(new_n1222), .A3(new_n1224), .A4(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(G159), .B2(new_n779), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n749), .B1(new_n1220), .B2(new_n1228), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1229), .B(new_n754), .C1(G68), .C2(new_n845), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n882), .B2(new_n734), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n1104), .B2(new_n753), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1213), .A2(new_n1232), .ZN(new_n1233));
  XOR2_X1   g1033(.A(new_n1233), .B(KEYINPUT123), .Z(G381));
  XOR2_X1   g1034(.A(G375), .B(KEYINPUT124), .Z(new_n1235));
  INV_X1    g1035(.A(G378), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1085), .B(new_n957), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1237));
  INV_X1    g1037(.A(G396), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1050), .A2(new_n1238), .A3(new_n1052), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(G381), .A2(G384), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1235), .A2(new_n1236), .A3(new_n1240), .A4(new_n1241), .ZN(G407));
  NAND3_X1  g1042(.A1(new_n1235), .A2(new_n659), .A3(new_n1236), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(G407), .A2(G213), .A3(new_n1243), .ZN(G409));
  NAND2_X1  g1044(.A1(G387), .A2(G390), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1050), .A2(new_n1238), .A3(new_n1052), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1238), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1247));
  OAI21_X1  g1047(.A(KEYINPUT127), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(G393), .A2(G396), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT127), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1249), .A2(new_n1239), .A3(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1245), .A2(new_n1252), .A3(new_n1237), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1251), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n1245), .B2(new_n1237), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1253), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT60), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1212), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1162), .A2(KEYINPUT60), .A3(new_n1180), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1258), .A2(new_n682), .A3(new_n1106), .A4(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(G384), .B1(new_n1260), .B2(new_n1232), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1260), .A2(G384), .A3(new_n1232), .ZN(new_n1263));
  INV_X1    g1063(.A(G213), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1264), .A2(G343), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(G2897), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1262), .A2(new_n1263), .A3(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1263), .ZN(new_n1268));
  OAI211_X1 g1068(.A(G2897), .B(new_n1265), .C1(new_n1268), .C2(new_n1261), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1182), .A2(KEYINPUT126), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT126), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1172), .A2(new_n1176), .A3(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(new_n753), .A3(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1163), .A2(new_n1002), .A3(new_n1177), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1273), .A2(new_n1274), .A3(new_n1209), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1236), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1184), .A2(G378), .A3(new_n1210), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT125), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1184), .A2(new_n1210), .A3(G378), .A4(KEYINPUT125), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1276), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1267), .B(new_n1269), .C1(new_n1281), .C2(new_n1265), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1268), .A2(new_n1261), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1281), .A2(new_n1265), .A3(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT62), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1282), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1276), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1265), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1290), .A2(new_n1286), .A3(new_n1291), .A4(new_n1283), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT61), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1256), .B1(new_n1287), .B2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1290), .A2(new_n1291), .A3(new_n1283), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1269), .A2(new_n1267), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1297), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT63), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1296), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1293), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1301), .B1(KEYINPUT63), .B2(new_n1285), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1300), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1295), .A2(new_n1303), .ZN(G405));
  NAND2_X1  g1104(.A1(G375), .A2(new_n1236), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1288), .A2(new_n1305), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1306), .B(new_n1283), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(new_n1307), .B(new_n1256), .ZN(G402));
endmodule


