//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 1 1 0 1 1 0 0 0 1 0 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1154, new_n1155, new_n1156, new_n1158, new_n1159,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1224, new_n1225;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OR2_X1    g0008(.A1(new_n206), .A2(KEYINPUT66), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n206), .A2(KEYINPUT66), .ZN(new_n210));
  NAND3_X1  g0010(.A1(new_n209), .A2(G50), .A3(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G20), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT65), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT0), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  AOI22_X1  g0021(.A1(new_n212), .A2(new_n217), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n222), .B1(new_n218), .B2(new_n221), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT67), .ZN(new_n224));
  AND2_X1   g0024(.A1(G107), .A2(G264), .ZN(new_n225));
  INV_X1    g0025(.A(G87), .ZN(new_n226));
  INV_X1    g0026(.A(G250), .ZN(new_n227));
  INV_X1    g0027(.A(G97), .ZN(new_n228));
  INV_X1    g0028(.A(G257), .ZN(new_n229));
  OAI22_X1  g0029(.A1(new_n226), .A2(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n225), .B(new_n230), .C1(G68), .C2(G238), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G50), .A2(G226), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G77), .A2(G244), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G116), .A2(G270), .ZN(new_n234));
  NAND4_X1  g0034(.A1(new_n231), .A2(new_n232), .A3(new_n233), .A4(new_n234), .ZN(new_n235));
  AND2_X1   g0035(.A1(G58), .A2(G232), .ZN(new_n236));
  OAI21_X1  g0036(.A(new_n219), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT1), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n224), .A2(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G264), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n241), .B(G270), .Z(new_n242));
  XOR2_X1   g0042(.A(G238), .B(G244), .Z(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G226), .B(G232), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n242), .B(new_n247), .ZN(G358));
  XNOR2_X1  g0048(.A(G68), .B(G77), .ZN(new_n249));
  INV_X1    g0049(.A(G50), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(G58), .ZN(new_n252));
  XOR2_X1   g0052(.A(G107), .B(G116), .Z(new_n253));
  XNOR2_X1  g0053(.A(G87), .B(G97), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n252), .B(new_n255), .ZN(G351));
  OAI21_X1  g0056(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT8), .B(G58), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G20), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n259), .A2(new_n261), .B1(G150), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n213), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G13), .ZN(new_n268));
  INV_X1    g0068(.A(G20), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n264), .A2(new_n266), .B1(new_n250), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n266), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n272), .B1(G1), .B2(new_n269), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n271), .B1(new_n250), .B2(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n274), .B(KEYINPUT9), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT3), .B(G33), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G222), .ZN(new_n278));
  INV_X1    g0078(.A(G223), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n276), .B(new_n278), .C1(new_n279), .C2(new_n277), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n214), .B1(new_n260), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n280), .B(new_n283), .C1(G77), .C2(new_n276), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n285));
  AND2_X1   g0085(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G226), .ZN(new_n287));
  INV_X1    g0087(.A(G274), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n284), .A2(new_n287), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G200), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT72), .ZN(new_n293));
  INV_X1    g0093(.A(G190), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(KEYINPUT10), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n275), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n297), .A2(KEYINPUT73), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(KEYINPUT73), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n275), .B(new_n292), .C1(new_n294), .C2(new_n291), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n298), .A2(new_n299), .B1(KEYINPUT10), .B2(new_n300), .ZN(new_n301));
  OR3_X1    g0101(.A1(new_n291), .A2(KEYINPUT69), .A3(G179), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n291), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT69), .B1(new_n291), .B2(G179), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n302), .A2(new_n274), .A3(new_n304), .A4(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(G58), .A2(G68), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n203), .A2(new_n205), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G20), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n262), .A2(G159), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT77), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AND2_X1   g0114(.A1(KEYINPUT3), .A2(G33), .ZN(new_n315));
  NOR2_X1   g0115(.A1(KEYINPUT3), .A2(G33), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(KEYINPUT7), .B1(new_n317), .B2(new_n269), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT7), .ZN(new_n319));
  NOR4_X1   g0119(.A1(new_n315), .A2(new_n316), .A3(new_n319), .A4(G20), .ZN(new_n320));
  OAI21_X1  g0120(.A(G68), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n310), .A2(KEYINPUT77), .A3(new_n311), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n314), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT16), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n314), .A2(KEYINPUT16), .A3(new_n321), .A4(new_n322), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(new_n266), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n270), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n258), .ZN(new_n329));
  INV_X1    g0129(.A(new_n273), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n329), .B1(new_n330), .B2(new_n258), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n279), .A2(new_n277), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n276), .B(new_n333), .C1(G226), .C2(new_n277), .ZN(new_n334));
  NAND2_X1  g0134(.A1(G33), .A2(G87), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n283), .ZN(new_n337));
  INV_X1    g0137(.A(G179), .ZN(new_n338));
  AND3_X1   g0138(.A1(new_n282), .A2(G232), .A3(new_n285), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n337), .A2(new_n338), .A3(new_n290), .A4(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n282), .B1(new_n334), .B2(new_n335), .ZN(new_n342));
  NOR3_X1   g0142(.A1(new_n342), .A2(new_n289), .A3(new_n339), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n341), .B1(new_n343), .B2(G169), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT18), .B1(new_n332), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT18), .ZN(new_n347));
  AOI211_X1 g0147(.A(new_n347), .B(new_n344), .C1(new_n327), .C2(new_n331), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n343), .A2(new_n294), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n343), .B2(G200), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n327), .A2(new_n351), .A3(new_n331), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT78), .B(KEYINPUT17), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT17), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n355), .A2(KEYINPUT78), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n327), .A2(new_n351), .A3(new_n331), .A4(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  NOR4_X1   g0158(.A1(new_n301), .A2(new_n307), .A3(new_n349), .A4(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(G226), .B(new_n277), .C1(new_n315), .C2(new_n316), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT74), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n276), .A2(KEYINPUT74), .A3(G226), .A4(new_n277), .ZN(new_n363));
  NAND2_X1  g0163(.A1(G33), .A2(G97), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n276), .A2(G232), .A3(G1698), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n362), .A2(new_n363), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n289), .B1(new_n366), .B2(new_n283), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT13), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n286), .A2(G238), .ZN(new_n369));
  AND3_X1   g0169(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n368), .B1(new_n367), .B2(new_n369), .ZN(new_n371));
  OAI21_X1  g0171(.A(G169), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(KEYINPUT76), .A2(KEYINPUT14), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n366), .A2(new_n283), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n376), .A2(new_n369), .A3(new_n290), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT13), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n380), .A2(G169), .A3(new_n373), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n370), .A2(new_n371), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G179), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n375), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n261), .A2(G77), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n202), .A2(G20), .ZN(new_n386));
  INV_X1    g0186(.A(new_n262), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n385), .B(new_n386), .C1(new_n250), .C2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n266), .ZN(new_n389));
  XOR2_X1   g0189(.A(new_n389), .B(KEYINPUT11), .Z(new_n390));
  NOR2_X1   g0190(.A1(new_n268), .A2(new_n386), .ZN(new_n391));
  XOR2_X1   g0191(.A(new_n391), .B(KEYINPUT12), .Z(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n202), .B2(new_n273), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n384), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT75), .B1(new_n380), .B2(G200), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n378), .A2(G190), .A3(new_n379), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n380), .A2(KEYINPUT75), .A3(G200), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n398), .A2(new_n394), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n276), .A2(G232), .A3(new_n277), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT70), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n276), .A2(G238), .A3(G1698), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n317), .A2(G107), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n276), .A2(KEYINPUT70), .A3(G232), .A4(new_n277), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n404), .A2(new_n405), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n283), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n286), .A2(G244), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n409), .A2(new_n290), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n338), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n328), .A2(G77), .ZN(new_n413));
  XOR2_X1   g0213(.A(KEYINPUT15), .B(G87), .Z(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n261), .ZN(new_n415));
  INV_X1    g0215(.A(G77), .ZN(new_n416));
  OAI221_X1 g0216(.A(new_n415), .B1(new_n269), .B2(new_n416), .C1(new_n387), .C2(new_n258), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n413), .B1(new_n417), .B2(new_n266), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n330), .A2(G77), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n409), .A2(new_n290), .A3(new_n410), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n303), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n412), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G200), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n420), .B1(new_n411), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT71), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT71), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n420), .B(new_n428), .C1(new_n411), .C2(new_n425), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n427), .B(new_n429), .C1(new_n294), .C2(new_n422), .ZN(new_n430));
  AND4_X1   g0230(.A1(new_n396), .A2(new_n401), .A3(new_n424), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n359), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  AOI211_X1 g0233(.A(new_n266), .B(new_n270), .C1(new_n267), .C2(G33), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(G116), .ZN(new_n435));
  AOI21_X1  g0235(.A(G20), .B1(G33), .B2(G283), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(G33), .B2(new_n228), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n437), .B(new_n266), .C1(new_n269), .C2(G116), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT85), .ZN(new_n439));
  OR2_X1    g0239(.A1(new_n439), .A2(KEYINPUT20), .ZN(new_n440));
  OR2_X1    g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n268), .A2(new_n269), .A3(G116), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n439), .A2(KEYINPUT20), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n438), .A2(new_n440), .A3(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n435), .A2(new_n441), .A3(new_n443), .A4(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(G45), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(G1), .ZN(new_n448));
  AND2_X1   g0248(.A1(KEYINPUT5), .A2(G41), .ZN(new_n449));
  NOR2_X1   g0249(.A1(KEYINPUT5), .A2(G41), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n451), .A2(new_n282), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G270), .ZN(new_n453));
  OR2_X1    g0253(.A1(new_n451), .A2(new_n288), .ZN(new_n454));
  INV_X1    g0254(.A(G303), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n317), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G264), .A2(G1698), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n457), .B1(new_n229), .B2(G1698), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n283), .B(new_n456), .C1(new_n317), .C2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n453), .A2(new_n454), .A3(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(new_n338), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n446), .A2(new_n461), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n460), .A2(G200), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n460), .A2(new_n294), .ZN(new_n464));
  OR3_X1    g0264(.A1(new_n463), .A2(new_n446), .A3(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n446), .A2(KEYINPUT21), .A3(G169), .A4(new_n460), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n446), .A2(G169), .A3(new_n460), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT21), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AND4_X1   g0269(.A1(new_n462), .A2(new_n465), .A3(new_n466), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n267), .A2(G45), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n260), .A2(new_n281), .ZN(new_n472));
  OAI211_X1 g0272(.A(G250), .B(new_n471), .C1(new_n472), .C2(new_n213), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n448), .A2(KEYINPUT82), .A3(G274), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT82), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(new_n471), .B2(new_n288), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n473), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n276), .A2(G238), .A3(new_n277), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n276), .A2(G244), .A3(G1698), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G116), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n477), .B1(new_n481), .B2(new_n283), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n482), .A2(KEYINPUT84), .A3(G190), .ZN(new_n483));
  AOI21_X1  g0283(.A(KEYINPUT84), .B1(new_n482), .B2(G190), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(G97), .A2(G107), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n226), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n364), .A2(new_n269), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n487), .A2(KEYINPUT19), .A3(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n269), .B(G68), .C1(new_n315), .C2(new_n316), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n364), .A2(G20), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n489), .B(new_n490), .C1(KEYINPUT19), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n266), .ZN(new_n493));
  INV_X1    g0293(.A(new_n414), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n270), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT83), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT83), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n493), .A2(new_n498), .A3(new_n495), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n497), .A2(new_n499), .B1(G87), .B2(new_n434), .ZN(new_n500));
  OR2_X1    g0300(.A1(new_n482), .A2(new_n425), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n485), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT23), .B1(new_n269), .B2(G107), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT23), .ZN(new_n504));
  INV_X1    g0304(.A(G107), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n504), .A2(new_n505), .A3(G20), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n269), .A2(G33), .A3(G116), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n503), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT86), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT86), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n503), .A2(new_n506), .A3(new_n507), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n269), .B(G87), .C1(new_n315), .C2(new_n316), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT22), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT22), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n276), .A2(new_n515), .A3(new_n269), .A4(G87), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT24), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n512), .A2(new_n517), .A3(KEYINPUT24), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n520), .A2(new_n266), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n434), .A2(G107), .ZN(new_n523));
  NOR2_X1   g0323(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(new_n328), .B2(G107), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n270), .B(new_n505), .C1(KEYINPUT87), .C2(KEYINPUT25), .ZN(new_n526));
  NAND2_X1  g0326(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n522), .A2(new_n523), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G294), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n276), .B1(G257), .B2(new_n277), .ZN(new_n531));
  NOR2_X1   g0331(.A1(G250), .A2(G1698), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n533), .A2(new_n283), .B1(new_n452), .B2(G264), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n454), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n303), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n534), .A2(new_n454), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n338), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n529), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n434), .A2(new_n414), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n493), .A2(new_n498), .A3(new_n495), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n498), .B1(new_n493), .B2(new_n495), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n482), .A2(new_n338), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n543), .B(new_n544), .C1(G169), .C2(new_n482), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n502), .A2(new_n539), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n434), .A2(G97), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n270), .A2(new_n228), .ZN(new_n548));
  XNOR2_X1  g0348(.A(new_n548), .B(KEYINPUT80), .ZN(new_n549));
  OAI21_X1  g0349(.A(G107), .B1(new_n318), .B2(new_n320), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT6), .ZN(new_n551));
  AND2_X1   g0351(.A1(G97), .A2(G107), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n551), .B1(new_n552), .B2(new_n486), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n505), .A2(KEYINPUT6), .A3(G97), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n555), .A2(G20), .B1(G77), .B2(new_n262), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n272), .B1(new_n550), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n557), .A2(KEYINPUT79), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT79), .ZN(new_n559));
  AOI211_X1 g0359(.A(new_n559), .B(new_n272), .C1(new_n550), .C2(new_n556), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n547), .B(new_n549), .C1(new_n558), .C2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(G250), .B(G1698), .C1(new_n315), .C2(new_n316), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT81), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n562), .A2(new_n563), .B1(G33), .B2(G283), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n276), .A2(KEYINPUT81), .A3(G250), .A4(G1698), .ZN(new_n565));
  OAI211_X1 g0365(.A(G244), .B(new_n277), .C1(new_n315), .C2(new_n316), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT4), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n276), .A2(KEYINPUT4), .A3(G244), .A4(new_n277), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n564), .A2(new_n565), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n283), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n452), .A2(G257), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n454), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n303), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n570), .A2(new_n283), .B1(G257), .B2(new_n452), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n575), .A2(new_n338), .A3(new_n454), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n561), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n547), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n555), .A2(G20), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n262), .A2(G77), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n319), .B1(new_n276), .B2(G20), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n317), .A2(KEYINPUT7), .A3(new_n269), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n505), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n266), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n559), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n557), .A2(KEYINPUT79), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n578), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n573), .A2(G200), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n575), .A2(G190), .A3(new_n454), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n588), .A2(new_n549), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n528), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n512), .A2(new_n517), .A3(KEYINPUT24), .ZN(new_n593));
  AOI21_X1  g0393(.A(KEYINPUT24), .B1(new_n512), .B2(new_n517), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n592), .B1(new_n595), .B2(new_n266), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n537), .A2(G190), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n535), .A2(G200), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n596), .A2(new_n597), .A3(new_n523), .A4(new_n598), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n577), .A2(new_n591), .A3(new_n599), .ZN(new_n600));
  AND4_X1   g0400(.A1(new_n433), .A2(new_n470), .A3(new_n546), .A4(new_n600), .ZN(G372));
  INV_X1    g0401(.A(new_n346), .ZN(new_n602));
  INV_X1    g0402(.A(new_n348), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT75), .ZN(new_n605));
  AOI211_X1 g0405(.A(new_n605), .B(new_n425), .C1(new_n378), .C2(new_n379), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n399), .A2(new_n394), .ZN(new_n607));
  NOR3_X1   g0407(.A1(new_n397), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT91), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n424), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n412), .A2(new_n421), .A3(KEYINPUT91), .A4(new_n423), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n608), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n612), .B1(new_n395), .B2(new_n384), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n604), .B1(new_n613), .B2(new_n358), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n298), .A2(new_n299), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n300), .A2(KEYINPUT10), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n307), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n543), .A2(new_n544), .ZN(new_n619));
  INV_X1    g0419(.A(new_n477), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n481), .A2(KEYINPUT88), .A3(new_n283), .ZN(new_n621));
  AOI21_X1  g0421(.A(KEYINPUT88), .B1(new_n481), .B2(new_n283), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n303), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n623), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n500), .B1(new_n626), .B2(new_n425), .ZN(new_n627));
  OR2_X1    g0427(.A1(new_n627), .A2(KEYINPUT89), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n627), .A2(KEYINPUT89), .B1(G190), .B2(new_n482), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n625), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n469), .A2(new_n466), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n462), .ZN(new_n632));
  INV_X1    g0432(.A(new_n539), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n630), .B(new_n600), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n502), .A2(new_n545), .ZN(new_n635));
  OAI21_X1  g0435(.A(KEYINPUT26), .B1(new_n635), .B2(new_n577), .ZN(new_n636));
  INV_X1    g0436(.A(new_n625), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  XNOR2_X1  g0438(.A(new_n577), .B(KEYINPUT90), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n630), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n634), .A2(new_n636), .A3(new_n637), .A4(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n618), .B1(new_n432), .B2(new_n642), .ZN(G369));
  OR3_X1    g0443(.A1(new_n268), .A2(KEYINPUT27), .A3(G20), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT27), .B1(new_n268), .B2(G20), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(G213), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(G343), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n446), .A2(new_n649), .ZN(new_n650));
  MUX2_X1   g0450(.A(new_n632), .B(new_n470), .S(new_n650), .Z(new_n651));
  AND2_X1   g0451(.A1(new_n651), .A2(G330), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n599), .A2(new_n539), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n648), .B1(new_n596), .B2(new_n523), .ZN(new_n654));
  OAI22_X1  g0454(.A1(new_n653), .A2(new_n654), .B1(new_n539), .B2(new_n648), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n632), .A2(new_n648), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(new_n653), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n648), .B(KEYINPUT92), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n658), .B1(new_n633), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n656), .A2(new_n660), .ZN(G399));
  NOR3_X1   g0461(.A1(new_n635), .A2(KEYINPUT26), .A3(new_n577), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n630), .A2(new_n639), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n662), .B1(new_n663), .B2(KEYINPUT26), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n664), .A2(new_n637), .A3(new_n634), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n665), .A2(KEYINPUT29), .A3(new_n648), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(KEYINPUT95), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT95), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n641), .A2(new_n659), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT29), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n667), .B1(new_n666), .B2(new_n671), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n600), .A2(new_n546), .A3(new_n470), .A4(new_n659), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n453), .A2(new_n454), .A3(new_n459), .ZN(new_n674));
  NOR4_X1   g0474(.A1(new_n626), .A2(new_n537), .A3(G179), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n573), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n674), .A2(G179), .A3(new_n534), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT30), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n677), .A2(new_n678), .A3(new_n482), .A4(new_n575), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n461), .A2(new_n575), .A3(new_n482), .A4(new_n534), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(KEYINPUT30), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n676), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n659), .ZN(new_n684));
  XNOR2_X1  g0484(.A(KEYINPUT94), .B(KEYINPUT31), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n675), .A2(new_n573), .B1(new_n681), .B2(new_n679), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(new_n648), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n673), .B(new_n686), .C1(KEYINPUT31), .C2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G330), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n672), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n267), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT93), .ZN(new_n693));
  INV_X1    g0493(.A(new_n220), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n693), .B1(new_n694), .B2(G41), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n220), .A2(KEYINPUT93), .A3(new_n281), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G116), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n486), .A2(new_n226), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n697), .A2(G1), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n211), .B2(new_n697), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT28), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n692), .A2(new_n703), .ZN(G364));
  INV_X1    g0504(.A(new_n697), .ZN(new_n705));
  INV_X1    g0505(.A(G13), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G20), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n267), .B1(new_n707), .B2(G45), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n651), .A2(G330), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n711), .B1(new_n713), .B2(new_n652), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n213), .B1(G20), .B2(new_n303), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n269), .A2(G190), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(new_n338), .A3(G200), .ZN(new_n717));
  OR2_X1    g0517(.A1(new_n717), .A2(KEYINPUT100), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(KEYINPUT100), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n505), .ZN(new_n721));
  NAND3_X1  g0521(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT99), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G190), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n721), .B1(G68), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n723), .A2(new_n294), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n725), .B(new_n276), .C1(new_n250), .C2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n269), .A2(new_n294), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n730), .A2(new_n425), .A3(G179), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n226), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n730), .A2(new_n338), .A3(G200), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G179), .A2(G200), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G190), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G20), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n734), .A2(G58), .B1(G97), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n716), .A2(G179), .A3(new_n425), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT98), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n739), .A2(new_n740), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n738), .B1(new_n744), .B2(new_n416), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n716), .A2(new_n735), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G159), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT32), .ZN(new_n749));
  NOR4_X1   g0549(.A1(new_n728), .A2(new_n733), .A3(new_n745), .A4(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n720), .ZN(new_n751));
  XNOR2_X1  g0551(.A(KEYINPUT33), .B(G317), .ZN(new_n752));
  AOI22_X1  g0552(.A1(new_n751), .A2(G283), .B1(new_n724), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(G311), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n753), .B1(new_n754), .B2(new_n744), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n726), .A2(G326), .ZN(new_n756));
  INV_X1    g0556(.A(new_n734), .ZN(new_n757));
  INV_X1    g0557(.A(G322), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n731), .A2(G303), .B1(G329), .B2(new_n747), .ZN(new_n760));
  INV_X1    g0560(.A(G294), .ZN(new_n761));
  INV_X1    g0561(.A(new_n737), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n760), .B(new_n317), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  NOR4_X1   g0563(.A1(new_n755), .A2(new_n756), .A3(new_n759), .A4(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n715), .B1(new_n750), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G13), .A2(G33), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n765), .B1(new_n651), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n768), .A2(new_n715), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n771), .B(KEYINPUT97), .Z(new_n772));
  NAND3_X1  g0572(.A1(new_n276), .A2(G355), .A3(new_n220), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n252), .A2(new_n447), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n317), .A2(new_n220), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT96), .Z(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(new_n211), .B2(G45), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n773), .B1(G116), .B2(new_n220), .C1(new_n774), .C2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n770), .B1(new_n772), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n714), .B1(new_n711), .B2(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT101), .Z(G396));
  NOR2_X1   g0581(.A1(new_n420), .A2(new_n648), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(new_n430), .B2(new_n424), .ZN(new_n783));
  AND3_X1   g0583(.A1(new_n610), .A2(new_n611), .A3(new_n782), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n641), .A2(new_n659), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(KEYINPUT102), .ZN(new_n787));
  INV_X1    g0587(.A(new_n785), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n669), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n787), .B(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(new_n690), .Z(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n711), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n727), .A2(new_n455), .B1(new_n762), .B2(new_n228), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(G283), .B2(new_n724), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n276), .B1(new_n731), .B2(G107), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n720), .A2(new_n226), .ZN(new_n796));
  INV_X1    g0596(.A(new_n744), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n796), .B1(G116), .B2(new_n797), .ZN(new_n798));
  AND3_X1   g0598(.A1(new_n794), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n799), .B1(new_n761), .B2(new_n757), .C1(new_n754), .C2(new_n746), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n724), .A2(G150), .B1(G143), .B2(new_n734), .ZN(new_n801));
  INV_X1    g0601(.A(G137), .ZN(new_n802));
  INV_X1    g0602(.A(G159), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n801), .B1(new_n802), .B2(new_n727), .C1(new_n803), .C2(new_n744), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT34), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n720), .A2(new_n202), .B1(new_n201), .B2(new_n762), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(G132), .B2(new_n747), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n805), .A2(new_n276), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n732), .A2(new_n250), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n800), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n711), .B1(new_n810), .B2(new_n715), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n715), .A2(new_n766), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n811), .B1(G77), .B2(new_n813), .C1(new_n767), .C2(new_n785), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n792), .A2(new_n814), .ZN(G384));
  OAI21_X1  g0615(.A(new_n618), .B1(new_n672), .B2(new_n432), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n395), .B(new_n649), .C1(new_n608), .C2(new_n384), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n395), .A2(new_n649), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n396), .A2(new_n401), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n424), .A2(new_n649), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n821), .B1(new_n786), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n332), .A2(new_n345), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n332), .A2(new_n647), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n825), .A2(new_n826), .A3(new_n352), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(KEYINPUT37), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT37), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n825), .A2(new_n826), .A3(new_n829), .A4(new_n352), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n646), .B1(new_n327), .B2(new_n331), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n349), .B2(new_n358), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT38), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n831), .A2(new_n833), .A3(KEYINPUT38), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n824), .A2(new_n838), .B1(new_n349), .B2(new_n646), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT103), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n838), .B1(new_n840), .B2(KEYINPUT39), .ZN(new_n841));
  XNOR2_X1  g0641(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n841), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n396), .A2(new_n649), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n839), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n816), .B(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n683), .A2(KEYINPUT31), .A3(new_n649), .ZN(new_n849));
  INV_X1    g0649(.A(new_n685), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n687), .B2(new_n648), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n673), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n433), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT40), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n831), .A2(new_n833), .A3(KEYINPUT38), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT38), .B1(new_n831), .B2(new_n833), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n820), .A2(new_n852), .A3(new_n785), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n854), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AND3_X1   g0659(.A1(new_n820), .A2(new_n852), .A3(new_n785), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n838), .A2(new_n860), .A3(KEYINPUT40), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n853), .B(new_n862), .Z(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(G330), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n848), .B(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n267), .B2(new_n707), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n698), .B1(new_n555), .B2(KEYINPUT35), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n217), .B(new_n867), .C1(KEYINPUT35), .C2(new_n555), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT36), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n212), .A2(G77), .A3(new_n308), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(G50), .B2(new_n202), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n871), .A2(G1), .A3(new_n706), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n866), .A2(new_n869), .A3(new_n872), .ZN(G367));
  NAND4_X1  g0673(.A1(new_n561), .A2(new_n684), .A3(new_n574), .A4(new_n576), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n874), .A2(KEYINPUT104), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n561), .A2(new_n684), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n577), .A2(new_n591), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n874), .A2(KEYINPUT104), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n875), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n660), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g0680(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n881));
  XNOR2_X1  g0681(.A(new_n880), .B(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n660), .A2(new_n879), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT45), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n656), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n885), .B(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n652), .A2(new_n655), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n657), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n658), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n691), .B1(new_n887), .B2(new_n892), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n697), .B(KEYINPUT41), .Z(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n708), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n500), .A2(new_n648), .ZN(new_n897));
  MUX2_X1   g0697(.A(new_n630), .B(new_n625), .S(new_n897), .Z(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT43), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n658), .A2(new_n879), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT42), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n879), .A2(new_n633), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n684), .B1(new_n902), .B2(new_n577), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n899), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n886), .A2(new_n879), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n904), .B(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n898), .A2(KEYINPUT43), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n906), .B(new_n907), .Z(new_n908));
  NAND2_X1  g0708(.A1(new_n896), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n776), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n771), .B1(new_n242), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n694), .B2(new_n414), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n746), .A2(new_n802), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n744), .A2(new_n250), .B1(new_n720), .B2(new_n416), .ZN(new_n914));
  INV_X1    g0714(.A(G143), .ZN(new_n915));
  INV_X1    g0715(.A(new_n724), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n915), .A2(new_n727), .B1(new_n916), .B2(new_n803), .ZN(new_n917));
  AOI211_X1 g0717(.A(new_n914), .B(new_n917), .C1(G68), .C2(new_n737), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n918), .B(new_n276), .C1(new_n201), .C2(new_n732), .ZN(new_n919));
  AOI211_X1 g0719(.A(new_n913), .B(new_n919), .C1(G150), .C2(new_n734), .ZN(new_n920));
  INV_X1    g0720(.A(G283), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n317), .B1(new_n744), .B2(new_n921), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n751), .A2(G97), .B1(G311), .B2(new_n726), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n747), .A2(G317), .B1(new_n737), .B2(G107), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n923), .B(new_n924), .C1(new_n455), .C2(new_n757), .ZN(new_n925));
  AOI211_X1 g0725(.A(new_n922), .B(new_n925), .C1(G294), .C2(new_n724), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n731), .A2(G116), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT46), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n920), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT47), .Z(new_n930));
  AOI21_X1  g0730(.A(new_n912), .B1(new_n930), .B2(new_n715), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n931), .B(new_n710), .C1(new_n769), .C2(new_n898), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n909), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(G387));
  NAND2_X1  g0734(.A1(new_n691), .A2(new_n891), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n672), .A2(new_n690), .A3(new_n892), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n935), .A2(new_n705), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n276), .A2(new_n699), .A3(new_n220), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n247), .A2(new_n447), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT106), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n700), .B(new_n447), .C1(new_n202), .C2(new_n416), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n258), .A2(G50), .ZN(new_n942));
  XOR2_X1   g0742(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n943));
  XNOR2_X1  g0743(.A(new_n942), .B(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n776), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  OAI221_X1 g0745(.A(new_n938), .B1(G107), .B2(new_n220), .C1(new_n940), .C2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n711), .B1(new_n946), .B2(new_n772), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT108), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n797), .A2(G303), .B1(new_n726), .B2(G322), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n734), .A2(G317), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n949), .B(new_n950), .C1(new_n754), .C2(new_n916), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT48), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n952), .B1(new_n921), .B2(new_n762), .C1(new_n761), .C2(new_n732), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT49), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n276), .B1(new_n747), .B2(G326), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n954), .B(new_n955), .C1(new_n698), .C2(new_n720), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n317), .B1(new_n747), .B2(G150), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n957), .B1(new_n732), .B2(new_n416), .C1(new_n720), .C2(new_n228), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT109), .Z(new_n959));
  NOR2_X1   g0759(.A1(new_n762), .A2(new_n494), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n744), .A2(new_n202), .B1(new_n727), .B2(new_n803), .ZN(new_n961));
  NOR3_X1   g0761(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n962), .B1(new_n250), .B2(new_n757), .C1(new_n258), .C2(new_n916), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n956), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n715), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n948), .B1(new_n655), .B2(new_n769), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n937), .B(new_n966), .C1(new_n708), .C2(new_n891), .ZN(G393));
  NAND2_X1  g0767(.A1(new_n887), .A2(new_n709), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n771), .B1(new_n228), .B2(new_n220), .C1(new_n910), .C2(new_n255), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n710), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT110), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n726), .A2(G150), .B1(G159), .B2(new_n734), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT111), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT51), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n796), .B1(G50), .B2(new_n724), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n731), .A2(G68), .B1(G77), .B2(new_n737), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n975), .A2(new_n276), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(new_n259), .B2(new_n797), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n974), .B(new_n978), .C1(new_n915), .C2(new_n746), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n721), .B1(G294), .B2(new_n797), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n698), .B2(new_n762), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n726), .A2(G317), .B1(G311), .B2(new_n734), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT52), .ZN(new_n983));
  NOR3_X1   g0783(.A1(new_n981), .A2(new_n276), .A3(new_n983), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n984), .B1(new_n921), .B2(new_n732), .C1(new_n455), .C2(new_n916), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n746), .A2(new_n758), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n979), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT112), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n971), .B1(new_n769), .B2(new_n879), .C1(new_n988), .C2(new_n965), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n887), .B(new_n936), .Z(new_n990));
  OAI211_X1 g0790(.A(new_n968), .B(new_n989), .C1(new_n990), .C2(new_n697), .ZN(G390));
  NOR2_X1   g0791(.A1(new_n857), .A2(new_n844), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n665), .A2(new_n648), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n822), .B1(new_n993), .B2(new_n785), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n992), .B1(new_n994), .B2(new_n821), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n841), .B1(new_n838), .B2(new_n842), .C1(new_n824), .C2(new_n844), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n689), .A2(G330), .A3(new_n785), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n998), .A2(new_n821), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n821), .A2(new_n788), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n852), .A2(G330), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n995), .B2(new_n996), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1001), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n821), .B1(new_n1003), .B2(new_n788), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n994), .A2(new_n999), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n998), .A2(new_n821), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1005), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n786), .A2(new_n823), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n433), .A2(G330), .A3(new_n852), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n618), .B(new_n1017), .C1(new_n672), .C2(new_n432), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1008), .A2(new_n1020), .A3(KEYINPUT113), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT113), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1007), .B1(new_n1022), .B2(new_n1019), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1021), .A2(new_n705), .A3(new_n1023), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n843), .A2(new_n767), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n731), .A2(G150), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT53), .Z(new_n1027));
  AOI22_X1  g0827(.A1(new_n1027), .A2(KEYINPUT114), .B1(G50), .B2(new_n751), .ZN(new_n1028));
  INV_X1    g0828(.A(G125), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1028), .B(new_n276), .C1(new_n1029), .C2(new_n746), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G137), .B2(new_n724), .ZN(new_n1031));
  XOR2_X1   g0831(.A(KEYINPUT54), .B(G143), .Z(new_n1032));
  NAND2_X1  g0832(.A1(new_n797), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n737), .A2(G159), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n726), .A2(G128), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n1027), .B2(KEYINPUT114), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(G132), .B2(new_n734), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .A4(new_n1037), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n720), .A2(new_n202), .B1(new_n416), .B2(new_n762), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n744), .A2(new_n228), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n317), .B1(new_n746), .B2(new_n761), .ZN(new_n1041));
  OR4_X1    g0841(.A1(new_n733), .A2(new_n1039), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(G107), .B2(new_n724), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n698), .B2(new_n757), .C1(new_n921), .C2(new_n727), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n965), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n711), .B(new_n1045), .C1(new_n258), .C2(new_n812), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n1007), .A2(new_n709), .B1(new_n1025), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1024), .A2(new_n1047), .ZN(G378));
  INV_X1    g0848(.A(KEYINPUT57), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n859), .A2(G330), .A3(new_n861), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(KEYINPUT119), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT119), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n859), .A2(new_n861), .A3(new_n1052), .A4(G330), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  XOR2_X1   g0854(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n617), .A2(new_n306), .A3(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1055), .B1(new_n301), .B2(new_n307), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n274), .A2(new_n647), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT117), .Z(new_n1060));
  AND3_X1   g0860(.A1(new_n1057), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1060), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1054), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1063), .B1(new_n1050), .B2(KEYINPUT119), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(KEYINPUT120), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1063), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT120), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1069), .A2(new_n1070), .A3(new_n1065), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n846), .B1(new_n1067), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT121), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1064), .A2(KEYINPUT120), .A3(new_n1066), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1070), .B1(new_n1069), .B2(new_n1065), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1077), .A2(KEYINPUT121), .A3(new_n846), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1079));
  OAI21_X1  g0879(.A(KEYINPUT122), .B1(new_n1079), .B2(new_n846), .ZN(new_n1080));
  OR4_X1    g0880(.A1(KEYINPUT122), .A2(new_n1069), .A3(new_n846), .A4(new_n1065), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1074), .A2(new_n1078), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1018), .B1(new_n1007), .B2(new_n1015), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1049), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT123), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1079), .B(new_n847), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n697), .B1(new_n1088), .B2(KEYINPUT57), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1081), .A2(new_n1080), .ZN(new_n1090));
  AOI21_X1  g0890(.A(KEYINPUT121), .B1(new_n1077), .B2(new_n846), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1073), .B(new_n847), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1090), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1083), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1095), .A2(KEYINPUT123), .A3(new_n1049), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1086), .A2(new_n1089), .A3(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n710), .B1(G50), .B2(new_n813), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n250), .B1(new_n315), .B2(G41), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n916), .A2(new_n228), .B1(new_n762), .B2(new_n202), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n746), .A2(new_n921), .ZN(new_n1101));
  NOR4_X1   g0901(.A1(new_n1100), .A2(G41), .A3(new_n276), .A4(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n726), .A2(G116), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n720), .A2(new_n201), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n416), .A2(new_n732), .B1(new_n757), .B2(new_n505), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n414), .B2(new_n797), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1102), .A2(new_n1103), .A3(new_n1105), .A4(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT58), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n797), .A2(G137), .B1(G128), .B2(new_n734), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n737), .A2(G150), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G132), .B2(new_n724), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n731), .A2(new_n1032), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT115), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1113), .B(new_n1115), .C1(new_n1029), .C2(new_n727), .ZN(new_n1116));
  AOI21_X1  g0916(.A(G33), .B1(new_n1116), .B2(KEYINPUT59), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n751), .A2(G159), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT116), .ZN(new_n1119));
  OR2_X1    g0919(.A1(new_n1119), .A2(G124), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(G124), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n747), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1117), .A2(new_n281), .A3(new_n1118), .A4(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1116), .A2(KEYINPUT59), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1099), .B(new_n1109), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1098), .B1(new_n1125), .B2(new_n715), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n1068), .B2(new_n767), .ZN(new_n1127));
  XOR2_X1   g0927(.A(new_n1127), .B(KEYINPUT118), .Z(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n1093), .B2(new_n709), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1097), .A2(new_n1129), .ZN(G375));
  NAND2_X1  g0930(.A1(new_n821), .A2(new_n766), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n813), .A2(G68), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n317), .B(new_n1104), .C1(G137), .C2(new_n734), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n724), .A2(new_n1032), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n747), .A2(G128), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n726), .A2(G132), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n250), .B2(new_n762), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(G150), .B2(new_n797), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .A4(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n732), .A2(new_n803), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n757), .A2(new_n921), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n746), .A2(new_n455), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1142), .B(new_n960), .C1(G116), .C2(new_n724), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n276), .B1(new_n797), .B2(G107), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n751), .A2(G77), .B1(G97), .B2(new_n731), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n726), .A2(G294), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n1139), .A2(new_n1140), .B1(new_n1141), .B2(new_n1147), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n711), .B(new_n1132), .C1(new_n1148), .C2(new_n715), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1015), .A2(new_n709), .B1(new_n1131), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1018), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n894), .B1(new_n1151), .B2(new_n1015), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1150), .B1(new_n1152), .B2(new_n1019), .ZN(G381));
  OR4_X1    g0953(.A1(G396), .A2(G387), .A3(G393), .A4(G390), .ZN(new_n1154));
  NOR3_X1   g0954(.A1(new_n1154), .A2(G384), .A3(G381), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(G375), .A2(G378), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(G407));
  INV_X1    g0957(.A(G343), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1156), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(G213), .ZN(G409));
  INV_X1    g0960(.A(G378), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1128), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1093), .A2(new_n894), .A3(new_n1094), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1087), .A2(new_n708), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1158), .A2(G213), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G375), .B2(G378), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1016), .A2(new_n1018), .A3(KEYINPUT60), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(KEYINPUT124), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT124), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1016), .A2(new_n1018), .A3(new_n1171), .A4(KEYINPUT60), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n697), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT125), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT60), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1175), .A2(new_n1019), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1173), .A2(new_n1174), .A3(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1174), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1150), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(G384), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  OAI211_X1 g0982(.A(G384), .B(new_n1150), .C1(new_n1178), .C2(new_n1179), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1168), .A2(new_n1184), .ZN(new_n1185));
  OR2_X1    g0985(.A1(new_n1185), .A2(KEYINPUT62), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT61), .ZN(new_n1187));
  AOI21_X1  g0987(.A(KEYINPUT123), .B1(new_n1095), .B2(new_n1049), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1085), .B(KEYINPUT57), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1089), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1129), .ZN(new_n1192));
  OAI21_X1  g0992(.A(G378), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1167), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1158), .A2(G213), .A3(G2897), .ZN(new_n1196));
  AND3_X1   g0996(.A1(new_n1182), .A2(new_n1183), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1196), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1195), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1185), .A2(KEYINPUT62), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1186), .A2(new_n1187), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n933), .B(G390), .ZN(new_n1203));
  XOR2_X1   g1003(.A(G393), .B(G396), .Z(new_n1204));
  XOR2_X1   g1004(.A(new_n1203), .B(new_n1204), .Z(new_n1205));
  NAND2_X1  g1005(.A1(new_n1202), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT127), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1200), .A2(KEYINPUT63), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT61), .B1(new_n1208), .B2(new_n1185), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1193), .A2(KEYINPUT63), .A3(new_n1184), .A4(new_n1194), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(KEYINPUT126), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT126), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1168), .A2(new_n1212), .A3(KEYINPUT63), .A4(new_n1184), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1205), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n1211), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1207), .B1(new_n1209), .B2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT63), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n1195), .B2(new_n1199), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1168), .A2(new_n1184), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1187), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1211), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n1220), .A2(new_n1221), .A3(KEYINPUT127), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1206), .B1(new_n1216), .B2(new_n1222), .ZN(G405));
  XNOR2_X1  g1023(.A(G375), .B(new_n1161), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(new_n1184), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1225), .B(new_n1205), .ZN(G402));
endmodule


