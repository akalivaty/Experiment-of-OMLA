

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589;

  XNOR2_X1 U322 ( .A(n426), .B(KEYINPUT48), .ZN(n556) );
  XNOR2_X1 U323 ( .A(n384), .B(n291), .ZN(n385) );
  NOR2_X1 U324 ( .A1(n540), .A2(n463), .ZN(n572) );
  INV_X1 U325 ( .A(n556), .ZN(n557) );
  AND2_X1 U326 ( .A1(G232GAT), .A2(G233GAT), .ZN(n290) );
  XOR2_X1 U327 ( .A(n383), .B(n382), .Z(n291) );
  INV_X1 U328 ( .A(KEYINPUT65), .ZN(n417) );
  XNOR2_X1 U329 ( .A(n417), .B(KEYINPUT45), .ZN(n418) );
  XNOR2_X1 U330 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U331 ( .A(n336), .B(n290), .ZN(n343) );
  XNOR2_X1 U332 ( .A(KEYINPUT54), .B(KEYINPUT123), .ZN(n443) );
  XNOR2_X1 U333 ( .A(n343), .B(n367), .ZN(n344) );
  XNOR2_X1 U334 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U335 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U336 ( .A(n354), .B(n353), .ZN(n414) );
  XOR2_X1 U337 ( .A(n388), .B(n580), .Z(n562) );
  XNOR2_X1 U338 ( .A(n467), .B(G190GAT), .ZN(n468) );
  XNOR2_X1 U339 ( .A(n469), .B(n468), .ZN(G1351GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT85), .B(KEYINPUT0), .Z(n293) );
  XNOR2_X1 U341 ( .A(KEYINPUT86), .B(G127GAT), .ZN(n292) );
  XNOR2_X1 U342 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U343 ( .A(G113GAT), .B(n294), .Z(n321) );
  XOR2_X1 U344 ( .A(KEYINPUT20), .B(G176GAT), .Z(n296) );
  XNOR2_X1 U345 ( .A(G15GAT), .B(KEYINPUT87), .ZN(n295) );
  XNOR2_X1 U346 ( .A(n296), .B(n295), .ZN(n308) );
  XOR2_X1 U347 ( .A(G120GAT), .B(G71GAT), .Z(n383) );
  XOR2_X1 U348 ( .A(G99GAT), .B(G190GAT), .Z(n298) );
  XNOR2_X1 U349 ( .A(G43GAT), .B(G134GAT), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U351 ( .A(n383), .B(n299), .Z(n301) );
  NAND2_X1 U352 ( .A1(G227GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U353 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U354 ( .A(n302), .B(KEYINPUT88), .Z(n306) );
  XOR2_X1 U355 ( .A(G183GAT), .B(KEYINPUT18), .Z(n304) );
  XNOR2_X1 U356 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n303) );
  XNOR2_X1 U357 ( .A(n304), .B(n303), .ZN(n439) );
  XNOR2_X1 U358 ( .A(G169GAT), .B(n439), .ZN(n305) );
  XNOR2_X1 U359 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U360 ( .A(n308), .B(n307), .Z(n309) );
  XOR2_X1 U361 ( .A(n321), .B(n309), .Z(n540) );
  XOR2_X1 U362 ( .A(G134GAT), .B(KEYINPUT79), .Z(n336) );
  XOR2_X1 U363 ( .A(G85GAT), .B(G162GAT), .Z(n311) );
  XNOR2_X1 U364 ( .A(G29GAT), .B(G148GAT), .ZN(n310) );
  XNOR2_X1 U365 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U366 ( .A(n336), .B(n312), .Z(n314) );
  NAND2_X1 U367 ( .A1(G225GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U368 ( .A(n314), .B(n313), .ZN(n333) );
  XOR2_X1 U369 ( .A(KEYINPUT97), .B(KEYINPUT93), .Z(n316) );
  XNOR2_X1 U370 ( .A(KEYINPUT96), .B(KEYINPUT1), .ZN(n315) );
  XNOR2_X1 U371 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U372 ( .A(G57GAT), .B(G155GAT), .Z(n318) );
  XNOR2_X1 U373 ( .A(G1GAT), .B(G120GAT), .ZN(n317) );
  XNOR2_X1 U374 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U375 ( .A(n320), .B(n319), .Z(n327) );
  INV_X1 U376 ( .A(n321), .ZN(n325) );
  XOR2_X1 U377 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n323) );
  XNOR2_X1 U378 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n322) );
  XNOR2_X1 U379 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U380 ( .A(n325), .B(n324), .Z(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U382 ( .A(n328), .B(KEYINPUT92), .Z(n331) );
  XNOR2_X1 U383 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n329) );
  XNOR2_X1 U384 ( .A(n329), .B(KEYINPUT2), .ZN(n446) );
  XNOR2_X1 U385 ( .A(n446), .B(KEYINPUT6), .ZN(n330) );
  XNOR2_X1 U386 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n513) );
  INV_X1 U388 ( .A(n513), .ZN(n528) );
  INV_X1 U389 ( .A(KEYINPUT47), .ZN(n413) );
  XOR2_X1 U390 ( .A(G99GAT), .B(G85GAT), .Z(n377) );
  XOR2_X1 U391 ( .A(G36GAT), .B(G190GAT), .Z(n437) );
  XOR2_X1 U392 ( .A(n377), .B(n437), .Z(n335) );
  XNOR2_X1 U393 ( .A(G218GAT), .B(G106GAT), .ZN(n334) );
  XNOR2_X1 U394 ( .A(n335), .B(n334), .ZN(n345) );
  INV_X1 U395 ( .A(G43GAT), .ZN(n337) );
  NAND2_X1 U396 ( .A1(n337), .A2(G29GAT), .ZN(n340) );
  INV_X1 U397 ( .A(G29GAT), .ZN(n338) );
  NAND2_X1 U398 ( .A1(n338), .A2(G43GAT), .ZN(n339) );
  NAND2_X1 U399 ( .A1(n340), .A2(n339), .ZN(n342) );
  XNOR2_X1 U400 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n341) );
  XNOR2_X1 U401 ( .A(n342), .B(n341), .ZN(n367) );
  XOR2_X1 U402 ( .A(n345), .B(n344), .Z(n354) );
  XOR2_X1 U403 ( .A(G50GAT), .B(G162GAT), .Z(n447) );
  XOR2_X1 U404 ( .A(KEYINPUT67), .B(KEYINPUT66), .Z(n347) );
  XNOR2_X1 U405 ( .A(KEYINPUT77), .B(KEYINPUT9), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n447), .B(n348), .ZN(n352) );
  XOR2_X1 U408 ( .A(KEYINPUT78), .B(KEYINPUT10), .Z(n350) );
  XNOR2_X1 U409 ( .A(G92GAT), .B(KEYINPUT11), .ZN(n349) );
  XOR2_X1 U410 ( .A(n350), .B(n349), .Z(n351) );
  XOR2_X1 U411 ( .A(KEYINPUT69), .B(KEYINPUT29), .Z(n356) );
  NAND2_X1 U412 ( .A1(G229GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U413 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U414 ( .A(n357), .B(KEYINPUT70), .Z(n365) );
  XOR2_X1 U415 ( .A(G22GAT), .B(G141GAT), .Z(n359) );
  XNOR2_X1 U416 ( .A(G50GAT), .B(G36GAT), .ZN(n358) );
  XNOR2_X1 U417 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U418 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n361) );
  XNOR2_X1 U419 ( .A(G197GAT), .B(G113GAT), .ZN(n360) );
  XNOR2_X1 U420 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U421 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U422 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U423 ( .A(G15GAT), .B(G1GAT), .Z(n393) );
  XOR2_X1 U424 ( .A(n366), .B(n393), .Z(n369) );
  XOR2_X1 U425 ( .A(G169GAT), .B(G8GAT), .Z(n440) );
  XNOR2_X1 U426 ( .A(n367), .B(n440), .ZN(n368) );
  XOR2_X1 U427 ( .A(n369), .B(n368), .Z(n510) );
  INV_X1 U428 ( .A(n510), .ZN(n576) );
  XNOR2_X1 U429 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n388) );
  XOR2_X1 U430 ( .A(G92GAT), .B(G64GAT), .Z(n371) );
  XNOR2_X1 U431 ( .A(G204GAT), .B(KEYINPUT74), .ZN(n370) );
  XNOR2_X1 U432 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U433 ( .A(G176GAT), .B(n372), .Z(n434) );
  XOR2_X1 U434 ( .A(G78GAT), .B(G148GAT), .Z(n374) );
  XNOR2_X1 U435 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n373) );
  XNOR2_X1 U436 ( .A(n374), .B(n373), .ZN(n450) );
  XOR2_X1 U437 ( .A(KEYINPUT71), .B(n450), .Z(n376) );
  NAND2_X1 U438 ( .A1(G230GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U439 ( .A(n376), .B(n375), .ZN(n386) );
  XOR2_X1 U440 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n379) );
  XOR2_X1 U441 ( .A(KEYINPUT13), .B(G57GAT), .Z(n396) );
  XNOR2_X1 U442 ( .A(n377), .B(n396), .ZN(n378) );
  XNOR2_X1 U443 ( .A(n379), .B(n378), .ZN(n384) );
  XOR2_X1 U444 ( .A(KEYINPUT76), .B(KEYINPUT73), .Z(n381) );
  XNOR2_X1 U445 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n380) );
  XNOR2_X1 U446 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U447 ( .A(n434), .B(n387), .Z(n580) );
  NAND2_X1 U448 ( .A1(n576), .A2(n562), .ZN(n389) );
  XNOR2_X1 U449 ( .A(KEYINPUT46), .B(n389), .ZN(n410) );
  XOR2_X1 U450 ( .A(G64GAT), .B(G78GAT), .Z(n391) );
  XNOR2_X1 U451 ( .A(G183GAT), .B(G211GAT), .ZN(n390) );
  XNOR2_X1 U452 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U453 ( .A(n392), .B(G71GAT), .Z(n395) );
  XNOR2_X1 U454 ( .A(n393), .B(G127GAT), .ZN(n394) );
  XNOR2_X1 U455 ( .A(n395), .B(n394), .ZN(n409) );
  XOR2_X1 U456 ( .A(n396), .B(KEYINPUT82), .Z(n398) );
  NAND2_X1 U457 ( .A1(G231GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U458 ( .A(n398), .B(n397), .ZN(n402) );
  XOR2_X1 U459 ( .A(KEYINPUT81), .B(KEYINPUT14), .Z(n400) );
  XNOR2_X1 U460 ( .A(KEYINPUT83), .B(KEYINPUT15), .ZN(n399) );
  XNOR2_X1 U461 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U462 ( .A(n402), .B(n401), .Z(n407) );
  XOR2_X1 U463 ( .A(G22GAT), .B(G155GAT), .Z(n448) );
  XOR2_X1 U464 ( .A(KEYINPUT84), .B(KEYINPUT12), .Z(n404) );
  XNOR2_X1 U465 ( .A(G8GAT), .B(KEYINPUT80), .ZN(n403) );
  XNOR2_X1 U466 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U467 ( .A(n448), .B(n405), .ZN(n406) );
  XNOR2_X1 U468 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U469 ( .A(n409), .B(n408), .ZN(n584) );
  INV_X1 U470 ( .A(n584), .ZN(n470) );
  NAND2_X1 U471 ( .A1(n410), .A2(n470), .ZN(n411) );
  NOR2_X1 U472 ( .A1(n414), .A2(n411), .ZN(n412) );
  XNOR2_X1 U473 ( .A(n413), .B(n412), .ZN(n425) );
  OR2_X1 U474 ( .A1(n414), .A2(KEYINPUT36), .ZN(n416) );
  NAND2_X1 U475 ( .A1(n414), .A2(KEYINPUT36), .ZN(n415) );
  NAND2_X1 U476 ( .A1(n416), .A2(n415), .ZN(n492) );
  NAND2_X1 U477 ( .A1(n492), .A2(n584), .ZN(n419) );
  NOR2_X1 U478 ( .A1(n580), .A2(n420), .ZN(n421) );
  XNOR2_X1 U479 ( .A(n421), .B(KEYINPUT113), .ZN(n422) );
  NOR2_X1 U480 ( .A1(n422), .A2(n576), .ZN(n423) );
  XNOR2_X1 U481 ( .A(KEYINPUT114), .B(n423), .ZN(n424) );
  NOR2_X1 U482 ( .A1(n425), .A2(n424), .ZN(n426) );
  XOR2_X1 U483 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n428) );
  NAND2_X1 U484 ( .A1(G226GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U485 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U486 ( .A(n429), .B(KEYINPUT80), .Z(n436) );
  XNOR2_X1 U487 ( .A(G211GAT), .B(KEYINPUT89), .ZN(n430) );
  XNOR2_X1 U488 ( .A(n430), .B(KEYINPUT21), .ZN(n431) );
  XOR2_X1 U489 ( .A(n431), .B(KEYINPUT90), .Z(n433) );
  XNOR2_X1 U490 ( .A(G197GAT), .B(G218GAT), .ZN(n432) );
  XNOR2_X1 U491 ( .A(n433), .B(n432), .ZN(n458) );
  XNOR2_X1 U492 ( .A(n458), .B(n434), .ZN(n435) );
  XNOR2_X1 U493 ( .A(n436), .B(n435), .ZN(n438) );
  XOR2_X1 U494 ( .A(n438), .B(n437), .Z(n442) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U496 ( .A(n442), .B(n441), .Z(n530) );
  INV_X1 U497 ( .A(n530), .ZN(n518) );
  NOR2_X1 U498 ( .A1(n556), .A2(n518), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n445) );
  NOR2_X1 U500 ( .A1(n528), .A2(n445), .ZN(n575) );
  XNOR2_X1 U501 ( .A(n447), .B(n446), .ZN(n449) );
  XNOR2_X1 U502 ( .A(n449), .B(n448), .ZN(n454) );
  XOR2_X1 U503 ( .A(n450), .B(KEYINPUT24), .Z(n452) );
  NAND2_X1 U504 ( .A1(G228GAT), .A2(G233GAT), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U506 ( .A(n454), .B(n453), .Z(n460) );
  XOR2_X1 U507 ( .A(KEYINPUT91), .B(G204GAT), .Z(n456) );
  XNOR2_X1 U508 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n455) );
  XNOR2_X1 U509 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U510 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U511 ( .A(n460), .B(n459), .ZN(n475) );
  NAND2_X1 U512 ( .A1(n575), .A2(n475), .ZN(n462) );
  XOR2_X1 U513 ( .A(KEYINPUT55), .B(KEYINPUT124), .Z(n461) );
  XNOR2_X1 U514 ( .A(n462), .B(n461), .ZN(n463) );
  NAND2_X1 U515 ( .A1(n572), .A2(n562), .ZN(n466) );
  XOR2_X1 U516 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n464) );
  XNOR2_X1 U517 ( .A(n464), .B(G176GAT), .ZN(n465) );
  XNOR2_X1 U518 ( .A(n466), .B(n465), .ZN(G1349GAT) );
  NAND2_X1 U519 ( .A1(n572), .A2(n414), .ZN(n469) );
  XOR2_X1 U520 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n467) );
  OR2_X1 U521 ( .A1(n510), .A2(n580), .ZN(n496) );
  NOR2_X1 U522 ( .A1(n414), .A2(n470), .ZN(n471) );
  XNOR2_X1 U523 ( .A(n471), .B(KEYINPUT16), .ZN(n483) );
  XNOR2_X1 U524 ( .A(n530), .B(KEYINPUT27), .ZN(n477) );
  NAND2_X1 U525 ( .A1(n477), .A2(n528), .ZN(n472) );
  XNOR2_X1 U526 ( .A(n472), .B(KEYINPUT100), .ZN(n559) );
  XNOR2_X1 U527 ( .A(n475), .B(KEYINPUT28), .ZN(n522) );
  INV_X1 U528 ( .A(n522), .ZN(n536) );
  NOR2_X1 U529 ( .A1(n559), .A2(n536), .ZN(n542) );
  NAND2_X1 U530 ( .A1(n540), .A2(n542), .ZN(n482) );
  INV_X1 U531 ( .A(n540), .ZN(n533) );
  NAND2_X1 U532 ( .A1(n533), .A2(n530), .ZN(n473) );
  NAND2_X1 U533 ( .A1(n475), .A2(n473), .ZN(n474) );
  XOR2_X1 U534 ( .A(KEYINPUT25), .B(n474), .Z(n479) );
  NOR2_X1 U535 ( .A1(n533), .A2(n475), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n476), .B(KEYINPUT26), .ZN(n574) );
  NAND2_X1 U537 ( .A1(n477), .A2(n574), .ZN(n478) );
  NAND2_X1 U538 ( .A1(n479), .A2(n478), .ZN(n480) );
  NAND2_X1 U539 ( .A1(n480), .A2(n513), .ZN(n481) );
  NAND2_X1 U540 ( .A1(n482), .A2(n481), .ZN(n493) );
  NAND2_X1 U541 ( .A1(n483), .A2(n493), .ZN(n511) );
  NOR2_X1 U542 ( .A1(n496), .A2(n511), .ZN(n484) );
  XOR2_X1 U543 ( .A(KEYINPUT101), .B(n484), .Z(n490) );
  NAND2_X1 U544 ( .A1(n490), .A2(n528), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n485), .B(KEYINPUT34), .ZN(n486) );
  XNOR2_X1 U546 ( .A(G1GAT), .B(n486), .ZN(G1324GAT) );
  NAND2_X1 U547 ( .A1(n530), .A2(n490), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n487), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U549 ( .A(G15GAT), .B(KEYINPUT35), .Z(n489) );
  NAND2_X1 U550 ( .A1(n490), .A2(n533), .ZN(n488) );
  XNOR2_X1 U551 ( .A(n489), .B(n488), .ZN(G1326GAT) );
  NAND2_X1 U552 ( .A1(n490), .A2(n536), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n491), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT104), .B(KEYINPUT39), .Z(n501) );
  NAND2_X1 U555 ( .A1(n492), .A2(n493), .ZN(n494) );
  NOR2_X1 U556 ( .A1(n584), .A2(n494), .ZN(n495) );
  XNOR2_X1 U557 ( .A(KEYINPUT37), .B(n495), .ZN(n527) );
  NOR2_X1 U558 ( .A1(n527), .A2(n496), .ZN(n499) );
  XOR2_X1 U559 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n497) );
  XNOR2_X1 U560 ( .A(KEYINPUT38), .B(n497), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n499), .B(n498), .ZN(n508) );
  NAND2_X1 U562 ( .A1(n508), .A2(n528), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U564 ( .A(G29GAT), .B(n502), .ZN(G1328GAT) );
  NAND2_X1 U565 ( .A1(n530), .A2(n508), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n503), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U567 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n507) );
  XOR2_X1 U568 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n505) );
  NAND2_X1 U569 ( .A1(n508), .A2(n533), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(G1330GAT) );
  NAND2_X1 U572 ( .A1(n508), .A2(n536), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n509), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U574 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n517) );
  NAND2_X1 U575 ( .A1(n510), .A2(n562), .ZN(n526) );
  NOR2_X1 U576 ( .A1(n526), .A2(n511), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(KEYINPUT107), .ZN(n521) );
  NOR2_X1 U578 ( .A1(n513), .A2(n521), .ZN(n515) );
  XNOR2_X1 U579 ( .A(G57GAT), .B(KEYINPUT109), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(G1332GAT) );
  NOR2_X1 U582 ( .A1(n518), .A2(n521), .ZN(n519) );
  XOR2_X1 U583 ( .A(G64GAT), .B(n519), .Z(G1333GAT) );
  NOR2_X1 U584 ( .A1(n540), .A2(n521), .ZN(n520) );
  XOR2_X1 U585 ( .A(G71GAT), .B(n520), .Z(G1334GAT) );
  NOR2_X1 U586 ( .A1(n522), .A2(n521), .ZN(n524) );
  XNOR2_X1 U587 ( .A(KEYINPUT43), .B(KEYINPUT110), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U589 ( .A(G78GAT), .B(n525), .ZN(G1335GAT) );
  NOR2_X1 U590 ( .A1(n527), .A2(n526), .ZN(n537) );
  NAND2_X1 U591 ( .A1(n528), .A2(n537), .ZN(n529) );
  XNOR2_X1 U592 ( .A(G85GAT), .B(n529), .ZN(G1336GAT) );
  XOR2_X1 U593 ( .A(G92GAT), .B(KEYINPUT111), .Z(n532) );
  NAND2_X1 U594 ( .A1(n537), .A2(n530), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n532), .B(n531), .ZN(G1337GAT) );
  NAND2_X1 U596 ( .A1(n533), .A2(n537), .ZN(n534) );
  XNOR2_X1 U597 ( .A(n534), .B(KEYINPUT112), .ZN(n535) );
  XNOR2_X1 U598 ( .A(G99GAT), .B(n535), .ZN(G1338GAT) );
  NAND2_X1 U599 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U600 ( .A(n538), .B(KEYINPUT44), .ZN(n539) );
  XNOR2_X1 U601 ( .A(G106GAT), .B(n539), .ZN(G1339GAT) );
  NOR2_X1 U602 ( .A1(n556), .A2(n540), .ZN(n541) );
  NAND2_X1 U603 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U604 ( .A(KEYINPUT115), .B(n543), .ZN(n552) );
  NAND2_X1 U605 ( .A1(n576), .A2(n552), .ZN(n544) );
  XNOR2_X1 U606 ( .A(KEYINPUT116), .B(n544), .ZN(n545) );
  XNOR2_X1 U607 ( .A(G113GAT), .B(n545), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n547) );
  NAND2_X1 U609 ( .A1(n552), .A2(n562), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U611 ( .A(G120GAT), .B(n548), .Z(G1341GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n550) );
  NAND2_X1 U613 ( .A1(n552), .A2(n584), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U615 ( .A(G127GAT), .B(n551), .Z(G1342GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n554) );
  NAND2_X1 U617 ( .A1(n552), .A2(n414), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U619 ( .A(G134GAT), .B(n555), .Z(G1343GAT) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(KEYINPUT120), .ZN(n561) );
  NAND2_X1 U621 ( .A1(n557), .A2(n574), .ZN(n558) );
  NOR2_X1 U622 ( .A1(n559), .A2(n558), .ZN(n569) );
  NAND2_X1 U623 ( .A1(n576), .A2(n569), .ZN(n560) );
  XNOR2_X1 U624 ( .A(n561), .B(n560), .ZN(G1344GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n564) );
  NAND2_X1 U626 ( .A1(n569), .A2(n562), .ZN(n563) );
  XNOR2_X1 U627 ( .A(n564), .B(n563), .ZN(n566) );
  XOR2_X1 U628 ( .A(G148GAT), .B(KEYINPUT52), .Z(n565) );
  XNOR2_X1 U629 ( .A(n566), .B(n565), .ZN(G1345GAT) );
  NAND2_X1 U630 ( .A1(n584), .A2(n569), .ZN(n567) );
  XNOR2_X1 U631 ( .A(n567), .B(KEYINPUT122), .ZN(n568) );
  XNOR2_X1 U632 ( .A(G155GAT), .B(n568), .ZN(G1346GAT) );
  NAND2_X1 U633 ( .A1(n569), .A2(n414), .ZN(n570) );
  XNOR2_X1 U634 ( .A(n570), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U635 ( .A1(n572), .A2(n576), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U637 ( .A1(n584), .A2(n572), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n578) );
  AND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n587) );
  NAND2_X1 U641 ( .A1(n587), .A2(n576), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n582) );
  NAND2_X1 U645 ( .A1(n587), .A2(n580), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G204GAT), .B(n583), .ZN(G1353GAT) );
  XOR2_X1 U648 ( .A(G211GAT), .B(KEYINPUT127), .Z(n586) );
  NAND2_X1 U649 ( .A1(n587), .A2(n584), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(G1354GAT) );
  NAND2_X1 U651 ( .A1(n492), .A2(n587), .ZN(n588) );
  XNOR2_X1 U652 ( .A(n588), .B(KEYINPUT62), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

